magic
tech sky130A
magscale 1 2
timestamp 1667937033
<< nwell >>
rect 882 87301 95074 87622
rect 882 86213 95074 86779
rect 882 85135 95074 85691
rect 882 85125 38011 85135
rect 882 84593 11515 84603
rect 882 84047 95074 84593
rect 882 84037 4352 84047
rect 882 83505 6928 83515
rect 882 82959 95074 83505
rect 882 82949 34975 82959
rect 882 82417 7651 82427
rect 882 81871 95074 82417
rect 882 81861 11147 81871
rect 882 81329 4904 81339
rect 882 80783 95074 81329
rect 882 80773 11252 80783
rect 882 80241 17035 80251
rect 882 79695 95074 80241
rect 882 79685 10871 79695
rect 882 79153 4891 79163
rect 882 78607 95074 79153
rect 882 78597 40311 78607
rect 882 78065 7940 78075
rect 882 77519 95074 78065
rect 882 77509 8939 77519
rect 882 76977 5180 76987
rect 882 76431 95074 76977
rect 882 76421 7559 76431
rect 882 75889 25223 75899
rect 882 75343 95074 75889
rect 882 75333 14919 75343
rect 882 74801 37275 74811
rect 882 74255 95074 74801
rect 882 74245 52192 74255
rect 882 73713 4536 73723
rect 882 73167 95074 73713
rect 882 73157 7940 73167
rect 882 72625 12067 72635
rect 882 72079 95074 72625
rect 882 72069 29547 72079
rect 882 71537 33871 71547
rect 882 70991 95074 71537
rect 882 70981 73431 70991
rect 882 70449 7743 70459
rect 882 69903 95074 70449
rect 882 69893 59644 69903
rect 882 69361 10135 69371
rect 882 68815 95074 69361
rect 882 68805 2972 68815
rect 882 68273 4628 68283
rect 882 67727 95074 68273
rect 882 67717 10227 67727
rect 882 67185 24027 67195
rect 882 66639 95074 67185
rect 882 66629 52547 66639
rect 882 66097 4996 66107
rect 882 65551 95074 66097
rect 882 65541 45003 65551
rect 882 65009 5548 65019
rect 882 64463 95074 65009
rect 882 64453 4996 64463
rect 882 63921 8479 63931
rect 882 63375 95074 63921
rect 882 63365 7467 63375
rect 882 62833 43991 62843
rect 882 62287 95074 62833
rect 882 62277 55491 62287
rect 882 61745 14459 61755
rect 882 61199 95074 61745
rect 882 61189 28548 61199
rect 882 60657 35895 60667
rect 882 60111 95074 60657
rect 882 60101 5364 60111
rect 882 59569 21819 59579
rect 882 59023 95074 59569
rect 882 59013 72419 59023
rect 882 58481 14104 58491
rect 882 57935 95074 58481
rect 882 57925 35251 57935
rect 882 57393 4996 57403
rect 882 56847 95074 57393
rect 882 56837 9215 56847
rect 882 56305 35816 56315
rect 882 55759 95074 56305
rect 882 55749 17035 55759
rect 882 54671 95074 55227
rect 882 54661 3971 54671
rect 882 54129 20439 54139
rect 882 53583 95074 54129
rect 882 53573 10779 53583
rect 882 53041 66544 53051
rect 882 52495 95074 53041
rect 882 52485 4904 52495
rect 882 51953 7835 51963
rect 882 51407 95074 51953
rect 882 51397 20176 51407
rect 882 50865 4444 50875
rect 882 50319 95074 50865
rect 882 50309 9583 50319
rect 882 49777 18704 49787
rect 882 49231 95074 49777
rect 882 49221 63403 49231
rect 882 48689 88795 48699
rect 882 48143 95074 48689
rect 882 48133 67635 48143
rect 882 47601 78491 47611
rect 882 47055 95074 47601
rect 882 47045 62220 47055
rect 882 46513 54952 46523
rect 882 45957 95074 46513
rect 882 45425 76283 45435
rect 882 44879 95074 45425
rect 882 44869 62759 44879
rect 882 44337 4720 44347
rect 882 43791 95074 44337
rect 882 43781 2604 43791
rect 882 43249 8755 43259
rect 882 42703 95074 43249
rect 882 42693 4352 42703
rect 882 42161 17771 42171
rect 882 41605 95074 42161
rect 882 41073 21819 41083
rect 882 40517 95074 41073
rect 882 39429 95074 39995
rect 882 38897 73339 38907
rect 882 38351 95074 38897
rect 882 38341 55307 38351
rect 882 37809 15103 37819
rect 882 37263 95074 37809
rect 882 37253 4812 37263
rect 882 36721 80055 36731
rect 882 36175 95074 36721
rect 882 36165 4904 36175
rect 882 35633 11515 35643
rect 882 35087 95074 35633
rect 882 35077 9872 35087
rect 882 34545 11515 34555
rect 882 33999 95074 34545
rect 882 33989 50720 33999
rect 882 33457 27615 33467
rect 882 32911 95074 33457
rect 882 32901 5088 32911
rect 882 32369 39023 32379
rect 882 31823 95074 32369
rect 882 31813 5535 31823
rect 882 31281 14735 31291
rect 882 30735 95074 31281
rect 882 30725 56424 30735
rect 882 30193 10332 30203
rect 882 29647 95074 30193
rect 882 29637 41415 29647
rect 882 29105 15484 29115
rect 882 28559 95074 29105
rect 882 28549 65703 28559
rect 882 28017 49616 28027
rect 882 27471 95074 28017
rect 882 27461 19243 27471
rect 882 26929 19703 26939
rect 882 26383 95074 26929
rect 882 26373 5995 26383
rect 882 25841 10516 25851
rect 882 25295 95074 25841
rect 882 25285 4444 25295
rect 882 24753 37275 24763
rect 882 24207 95074 24753
rect 882 24197 16391 24207
rect 882 23665 10240 23675
rect 882 23119 95074 23665
rect 882 23109 12540 23119
rect 882 22031 95074 22587
rect 882 22021 17219 22031
rect 882 21489 38931 21499
rect 882 20943 95074 21489
rect 882 20933 6087 20943
rect 882 20401 4720 20411
rect 882 19855 95074 20401
rect 882 19845 27983 19855
rect 882 19313 22555 19323
rect 882 18767 95074 19313
rect 882 18757 31847 18767
rect 882 18225 48144 18235
rect 882 17679 95074 18225
rect 882 17669 81067 17679
rect 882 17137 10424 17147
rect 882 16591 95074 17137
rect 882 16581 17863 16591
rect 882 16049 10135 16059
rect 882 15503 95074 16049
rect 882 15493 2420 15503
rect 882 14961 12080 14971
rect 882 14415 95074 14961
rect 882 14405 6100 14415
rect 882 13873 30743 13883
rect 882 13327 95074 13873
rect 882 13317 73431 13327
rect 882 12785 37827 12795
rect 882 12239 95074 12785
rect 882 12229 4339 12239
rect 882 11697 7007 11707
rect 882 11151 95074 11697
rect 882 11141 4628 11151
rect 882 10609 73339 10619
rect 882 10063 95074 10609
rect 882 10053 63035 10063
rect 882 9521 28351 9531
rect 882 8975 95074 9521
rect 882 8965 18428 8975
rect 882 8433 10135 8443
rect 882 7887 95074 8433
rect 882 7877 20176 7887
rect 882 7345 9136 7355
rect 882 6799 95074 7345
rect 882 6789 39036 6799
rect 882 6257 3984 6267
rect 882 5711 95074 6257
rect 882 5701 5535 5711
rect 882 5169 16667 5179
rect 882 4623 95074 5169
rect 882 4613 55767 4623
rect 882 4081 89531 4091
rect 882 3525 95074 4081
rect 882 2437 95074 3003
<< obsli1 >>
rect 920 2159 95036 87601
<< obsm1 >>
rect 920 1980 95114 87848
<< metal2 >>
rect 2318 89200 2374 90000
rect 5262 89200 5318 90000
rect 8206 89200 8262 90000
rect 11150 89200 11206 90000
rect 14094 89200 14150 90000
rect 17038 89200 17094 90000
rect 19982 89200 20038 90000
rect 22926 89200 22982 90000
rect 25870 89200 25926 90000
rect 28814 89200 28870 90000
rect 31758 89200 31814 90000
rect 34702 89200 34758 90000
rect 37646 89200 37702 90000
rect 40590 89200 40646 90000
rect 43534 89200 43590 90000
rect 46478 89200 46534 90000
rect 49422 89200 49478 90000
rect 52366 89200 52422 90000
rect 55310 89200 55366 90000
rect 58254 89200 58310 90000
rect 61198 89200 61254 90000
rect 64142 89200 64198 90000
rect 67086 89200 67142 90000
rect 70030 89200 70086 90000
rect 72974 89200 73030 90000
rect 75918 89200 75974 90000
rect 78862 89200 78918 90000
rect 81806 89200 81862 90000
rect 84750 89200 84806 90000
rect 87694 89200 87750 90000
rect 90638 89200 90694 90000
rect 93582 89200 93638 90000
<< obsm2 >>
rect 1400 89144 2262 89298
rect 2430 89144 5206 89298
rect 5374 89144 8150 89298
rect 8318 89144 11094 89298
rect 11262 89144 14038 89298
rect 14206 89144 16982 89298
rect 17150 89144 19926 89298
rect 20094 89144 22870 89298
rect 23038 89144 25814 89298
rect 25982 89144 28758 89298
rect 28926 89144 31702 89298
rect 31870 89144 34646 89298
rect 34814 89144 37590 89298
rect 37758 89144 40534 89298
rect 40702 89144 43478 89298
rect 43646 89144 46422 89298
rect 46590 89144 49366 89298
rect 49534 89144 52310 89298
rect 52478 89144 55254 89298
rect 55422 89144 58198 89298
rect 58366 89144 61142 89298
rect 61310 89144 64086 89298
rect 64254 89144 67030 89298
rect 67198 89144 69974 89298
rect 70142 89144 72918 89298
rect 73086 89144 75862 89298
rect 76030 89144 78806 89298
rect 78974 89144 81750 89298
rect 81918 89144 84694 89298
rect 84862 89144 87638 89298
rect 87806 89144 90582 89298
rect 90750 89144 93526 89298
rect 93694 89144 95108 89298
rect 1400 1974 95108 89144
<< metal3 >>
rect 95200 86776 96000 86896
rect 95200 84872 96000 84992
rect 95200 82968 96000 83088
rect 95200 81064 96000 81184
rect 95200 79160 96000 79280
rect 95200 77256 96000 77376
rect 95200 75352 96000 75472
rect 95200 73448 96000 73568
rect 95200 71544 96000 71664
rect 95200 69640 96000 69760
rect 95200 67736 96000 67856
rect 95200 65832 96000 65952
rect 95200 63928 96000 64048
rect 95200 62024 96000 62144
rect 95200 60120 96000 60240
rect 95200 58216 96000 58336
rect 95200 56312 96000 56432
rect 95200 54408 96000 54528
rect 95200 52504 96000 52624
rect 95200 50600 96000 50720
rect 95200 48696 96000 48816
rect 95200 46792 96000 46912
rect 95200 44888 96000 45008
rect 95200 42984 96000 43104
rect 95200 41080 96000 41200
rect 95200 39176 96000 39296
rect 95200 37272 96000 37392
rect 95200 35368 96000 35488
rect 95200 33464 96000 33584
rect 95200 31560 96000 31680
rect 95200 29656 96000 29776
rect 95200 27752 96000 27872
rect 95200 25848 96000 25968
rect 95200 23944 96000 24064
rect 95200 22040 96000 22160
rect 95200 20136 96000 20256
rect 95200 18232 96000 18352
rect 95200 16328 96000 16448
rect 95200 14424 96000 14544
rect 95200 12520 96000 12640
rect 95200 10616 96000 10736
rect 95200 8712 96000 8832
rect 95200 6808 96000 6928
rect 95200 4904 96000 5024
rect 95200 3000 96000 3120
<< obsm3 >>
rect 1853 86976 95200 87617
rect 1853 86696 95120 86976
rect 1853 85072 95200 86696
rect 1853 84792 95120 85072
rect 1853 83168 95200 84792
rect 1853 82888 95120 83168
rect 1853 81264 95200 82888
rect 1853 80984 95120 81264
rect 1853 79360 95200 80984
rect 1853 79080 95120 79360
rect 1853 77456 95200 79080
rect 1853 77176 95120 77456
rect 1853 75552 95200 77176
rect 1853 75272 95120 75552
rect 1853 73648 95200 75272
rect 1853 73368 95120 73648
rect 1853 71744 95200 73368
rect 1853 71464 95120 71744
rect 1853 69840 95200 71464
rect 1853 69560 95120 69840
rect 1853 67936 95200 69560
rect 1853 67656 95120 67936
rect 1853 66032 95200 67656
rect 1853 65752 95120 66032
rect 1853 64128 95200 65752
rect 1853 63848 95120 64128
rect 1853 62224 95200 63848
rect 1853 61944 95120 62224
rect 1853 60320 95200 61944
rect 1853 60040 95120 60320
rect 1853 58416 95200 60040
rect 1853 58136 95120 58416
rect 1853 56512 95200 58136
rect 1853 56232 95120 56512
rect 1853 54608 95200 56232
rect 1853 54328 95120 54608
rect 1853 52704 95200 54328
rect 1853 52424 95120 52704
rect 1853 50800 95200 52424
rect 1853 50520 95120 50800
rect 1853 48896 95200 50520
rect 1853 48616 95120 48896
rect 1853 46992 95200 48616
rect 1853 46712 95120 46992
rect 1853 45088 95200 46712
rect 1853 44808 95120 45088
rect 1853 43184 95200 44808
rect 1853 42904 95120 43184
rect 1853 41280 95200 42904
rect 1853 41000 95120 41280
rect 1853 39376 95200 41000
rect 1853 39096 95120 39376
rect 1853 37472 95200 39096
rect 1853 37192 95120 37472
rect 1853 35568 95200 37192
rect 1853 35288 95120 35568
rect 1853 33664 95200 35288
rect 1853 33384 95120 33664
rect 1853 31760 95200 33384
rect 1853 31480 95120 31760
rect 1853 29856 95200 31480
rect 1853 29576 95120 29856
rect 1853 27952 95200 29576
rect 1853 27672 95120 27952
rect 1853 26048 95200 27672
rect 1853 25768 95120 26048
rect 1853 24144 95200 25768
rect 1853 23864 95120 24144
rect 1853 22240 95200 23864
rect 1853 21960 95120 22240
rect 1853 20336 95200 21960
rect 1853 20056 95120 20336
rect 1853 18432 95200 20056
rect 1853 18152 95120 18432
rect 1853 16528 95200 18152
rect 1853 16248 95120 16528
rect 1853 14624 95200 16248
rect 1853 14344 95120 14624
rect 1853 12720 95200 14344
rect 1853 12440 95120 12720
rect 1853 10816 95200 12440
rect 1853 10536 95120 10816
rect 1853 8912 95200 10536
rect 1853 8632 95120 8912
rect 1853 7008 95200 8632
rect 1853 6728 95120 7008
rect 1853 5104 95200 6728
rect 1853 4824 95120 5104
rect 1853 3200 95200 4824
rect 1853 2920 95120 3200
rect 1853 2143 95200 2920
<< metal4 >>
rect 4024 2128 4344 87632
rect 19384 2128 19704 87632
rect 34744 2128 35064 87632
rect 50104 2128 50424 87632
rect 65464 2128 65784 87632
rect 80824 2128 81144 87632
<< obsm4 >>
rect 3371 6835 3944 86733
rect 4424 6835 19304 86733
rect 19784 6835 34664 86733
rect 35144 6835 50024 86733
rect 50504 6835 65384 86733
rect 65864 6835 80744 86733
rect 81224 6835 91757 86733
<< labels >>
rlabel metal3 s 95200 3000 96000 3120 6 A0[0]
port 1 nsew signal input
rlabel metal3 s 95200 4904 96000 5024 6 A0[1]
port 2 nsew signal input
rlabel metal3 s 95200 6808 96000 6928 6 A0[2]
port 3 nsew signal input
rlabel metal3 s 95200 8712 96000 8832 6 A0[3]
port 4 nsew signal input
rlabel metal3 s 95200 10616 96000 10736 6 A0[4]
port 5 nsew signal input
rlabel metal3 s 95200 12520 96000 12640 6 A0[5]
port 6 nsew signal input
rlabel metal3 s 95200 14424 96000 14544 6 A0[6]
port 7 nsew signal input
rlabel metal3 s 95200 56312 96000 56432 6 CLK
port 8 nsew signal input
rlabel metal3 s 95200 25848 96000 25968 6 Di0[0]
port 9 nsew signal input
rlabel metal3 s 95200 44888 96000 45008 6 Di0[10]
port 10 nsew signal input
rlabel metal3 s 95200 46792 96000 46912 6 Di0[11]
port 11 nsew signal input
rlabel metal3 s 95200 48696 96000 48816 6 Di0[12]
port 12 nsew signal input
rlabel metal3 s 95200 50600 96000 50720 6 Di0[13]
port 13 nsew signal input
rlabel metal3 s 95200 52504 96000 52624 6 Di0[14]
port 14 nsew signal input
rlabel metal3 s 95200 54408 96000 54528 6 Di0[15]
port 15 nsew signal input
rlabel metal3 s 95200 58216 96000 58336 6 Di0[16]
port 16 nsew signal input
rlabel metal3 s 95200 60120 96000 60240 6 Di0[17]
port 17 nsew signal input
rlabel metal3 s 95200 62024 96000 62144 6 Di0[18]
port 18 nsew signal input
rlabel metal3 s 95200 63928 96000 64048 6 Di0[19]
port 19 nsew signal input
rlabel metal3 s 95200 27752 96000 27872 6 Di0[1]
port 20 nsew signal input
rlabel metal3 s 95200 65832 96000 65952 6 Di0[20]
port 21 nsew signal input
rlabel metal3 s 95200 67736 96000 67856 6 Di0[21]
port 22 nsew signal input
rlabel metal3 s 95200 69640 96000 69760 6 Di0[22]
port 23 nsew signal input
rlabel metal3 s 95200 71544 96000 71664 6 Di0[23]
port 24 nsew signal input
rlabel metal3 s 95200 73448 96000 73568 6 Di0[24]
port 25 nsew signal input
rlabel metal3 s 95200 75352 96000 75472 6 Di0[25]
port 26 nsew signal input
rlabel metal3 s 95200 77256 96000 77376 6 Di0[26]
port 27 nsew signal input
rlabel metal3 s 95200 79160 96000 79280 6 Di0[27]
port 28 nsew signal input
rlabel metal3 s 95200 81064 96000 81184 6 Di0[28]
port 29 nsew signal input
rlabel metal3 s 95200 82968 96000 83088 6 Di0[29]
port 30 nsew signal input
rlabel metal3 s 95200 29656 96000 29776 6 Di0[2]
port 31 nsew signal input
rlabel metal3 s 95200 84872 96000 84992 6 Di0[30]
port 32 nsew signal input
rlabel metal3 s 95200 86776 96000 86896 6 Di0[31]
port 33 nsew signal input
rlabel metal3 s 95200 31560 96000 31680 6 Di0[3]
port 34 nsew signal input
rlabel metal3 s 95200 33464 96000 33584 6 Di0[4]
port 35 nsew signal input
rlabel metal3 s 95200 35368 96000 35488 6 Di0[5]
port 36 nsew signal input
rlabel metal3 s 95200 37272 96000 37392 6 Di0[6]
port 37 nsew signal input
rlabel metal3 s 95200 39176 96000 39296 6 Di0[7]
port 38 nsew signal input
rlabel metal3 s 95200 41080 96000 41200 6 Di0[8]
port 39 nsew signal input
rlabel metal3 s 95200 42984 96000 43104 6 Di0[9]
port 40 nsew signal input
rlabel metal2 s 2318 89200 2374 90000 6 Do0[0]
port 41 nsew signal output
rlabel metal2 s 31758 89200 31814 90000 6 Do0[10]
port 42 nsew signal output
rlabel metal2 s 34702 89200 34758 90000 6 Do0[11]
port 43 nsew signal output
rlabel metal2 s 37646 89200 37702 90000 6 Do0[12]
port 44 nsew signal output
rlabel metal2 s 40590 89200 40646 90000 6 Do0[13]
port 45 nsew signal output
rlabel metal2 s 43534 89200 43590 90000 6 Do0[14]
port 46 nsew signal output
rlabel metal2 s 46478 89200 46534 90000 6 Do0[15]
port 47 nsew signal output
rlabel metal2 s 49422 89200 49478 90000 6 Do0[16]
port 48 nsew signal output
rlabel metal2 s 52366 89200 52422 90000 6 Do0[17]
port 49 nsew signal output
rlabel metal2 s 55310 89200 55366 90000 6 Do0[18]
port 50 nsew signal output
rlabel metal2 s 58254 89200 58310 90000 6 Do0[19]
port 51 nsew signal output
rlabel metal2 s 5262 89200 5318 90000 6 Do0[1]
port 52 nsew signal output
rlabel metal2 s 61198 89200 61254 90000 6 Do0[20]
port 53 nsew signal output
rlabel metal2 s 64142 89200 64198 90000 6 Do0[21]
port 54 nsew signal output
rlabel metal2 s 67086 89200 67142 90000 6 Do0[22]
port 55 nsew signal output
rlabel metal2 s 70030 89200 70086 90000 6 Do0[23]
port 56 nsew signal output
rlabel metal2 s 72974 89200 73030 90000 6 Do0[24]
port 57 nsew signal output
rlabel metal2 s 75918 89200 75974 90000 6 Do0[25]
port 58 nsew signal output
rlabel metal2 s 78862 89200 78918 90000 6 Do0[26]
port 59 nsew signal output
rlabel metal2 s 81806 89200 81862 90000 6 Do0[27]
port 60 nsew signal output
rlabel metal2 s 84750 89200 84806 90000 6 Do0[28]
port 61 nsew signal output
rlabel metal2 s 87694 89200 87750 90000 6 Do0[29]
port 62 nsew signal output
rlabel metal2 s 8206 89200 8262 90000 6 Do0[2]
port 63 nsew signal output
rlabel metal2 s 90638 89200 90694 90000 6 Do0[30]
port 64 nsew signal output
rlabel metal2 s 93582 89200 93638 90000 6 Do0[31]
port 65 nsew signal output
rlabel metal2 s 11150 89200 11206 90000 6 Do0[3]
port 66 nsew signal output
rlabel metal2 s 14094 89200 14150 90000 6 Do0[4]
port 67 nsew signal output
rlabel metal2 s 17038 89200 17094 90000 6 Do0[5]
port 68 nsew signal output
rlabel metal2 s 19982 89200 20038 90000 6 Do0[6]
port 69 nsew signal output
rlabel metal2 s 22926 89200 22982 90000 6 Do0[7]
port 70 nsew signal output
rlabel metal2 s 25870 89200 25926 90000 6 Do0[8]
port 71 nsew signal output
rlabel metal2 s 28814 89200 28870 90000 6 Do0[9]
port 72 nsew signal output
rlabel metal3 s 95200 23944 96000 24064 6 EN0
port 73 nsew signal input
rlabel metal4 s 19384 2128 19704 87632 6 VGND
port 74 nsew ground bidirectional
rlabel metal4 s 50104 2128 50424 87632 6 VGND
port 74 nsew ground bidirectional
rlabel metal4 s 80824 2128 81144 87632 6 VGND
port 74 nsew ground bidirectional
rlabel metal4 s 4024 2128 4344 87632 6 VPWR
port 75 nsew power bidirectional
rlabel metal4 s 34744 2128 35064 87632 6 VPWR
port 75 nsew power bidirectional
rlabel metal4 s 65464 2128 65784 87632 6 VPWR
port 75 nsew power bidirectional
rlabel metal3 s 95200 16328 96000 16448 6 WE0[0]
port 76 nsew signal input
rlabel metal3 s 95200 18232 96000 18352 6 WE0[1]
port 77 nsew signal input
rlabel metal3 s 95200 20136 96000 20256 6 WE0[2]
port 78 nsew signal input
rlabel metal3 s 95200 22040 96000 22160 6 WE0[3]
port 79 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 96000 90000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 30504172
string GDS_FILE /home/hosni/RAM128/caravel_mgmt_soc_litex/openlane/RAM128/runs/RUN_2022.11.08_19.33.51/results/signoff/RAM128.magic.gds
string GDS_START 166586
<< end >>

