magic
tech sky130A
magscale 1 2
timestamp 1638404839
<< metal1 >>
rect 126330 160080 126336 160132
rect 126388 160120 126394 160132
rect 128354 160120 128360 160132
rect 126388 160092 128360 160120
rect 126388 160080 126394 160092
rect 128354 160080 128360 160092
rect 128412 160080 128418 160132
rect 153010 160080 153016 160132
rect 153068 160120 153074 160132
rect 153068 160092 154620 160120
rect 153068 160080 153074 160092
rect 66714 160012 66720 160064
rect 66772 160052 66778 160064
rect 142798 160052 142804 160064
rect 66772 160024 142804 160052
rect 66772 160012 66778 160024
rect 142798 160012 142804 160024
rect 142856 160012 142862 160064
rect 142890 160012 142896 160064
rect 142948 160052 142954 160064
rect 154482 160052 154488 160064
rect 142948 160024 154488 160052
rect 142948 160012 142954 160024
rect 154482 160012 154488 160024
rect 154540 160012 154546 160064
rect 154592 160052 154620 160092
rect 331186 160092 331444 160120
rect 158806 160052 158812 160064
rect 154592 160024 158812 160052
rect 158806 160012 158812 160024
rect 158864 160012 158870 160064
rect 159910 160012 159916 160064
rect 159968 160052 159974 160064
rect 196158 160052 196164 160064
rect 159968 160024 196164 160052
rect 159968 160012 159974 160024
rect 196158 160012 196164 160024
rect 196216 160012 196222 160064
rect 207750 160012 207756 160064
rect 207808 160052 207814 160064
rect 276106 160052 276112 160064
rect 207808 160024 276112 160052
rect 207808 160012 207814 160024
rect 276106 160012 276112 160024
rect 276164 160012 276170 160064
rect 277486 160012 277492 160064
rect 277544 160052 277550 160064
rect 280154 160052 280160 160064
rect 277544 160024 280160 160052
rect 277544 160012 277550 160024
rect 280154 160012 280160 160024
rect 280212 160012 280218 160064
rect 280798 160012 280804 160064
rect 280856 160052 280862 160064
rect 331186 160052 331214 160092
rect 280856 160024 331214 160052
rect 280856 160012 280862 160024
rect 76742 159944 76748 159996
rect 76800 159984 76806 159996
rect 164510 159984 164516 159996
rect 76800 159956 164516 159984
rect 76800 159944 76806 159956
rect 164510 159944 164516 159956
rect 164568 159944 164574 159996
rect 166626 159944 166632 159996
rect 166684 159984 166690 159996
rect 197630 159984 197636 159996
rect 166684 159956 197636 159984
rect 166684 159944 166690 159956
rect 197630 159944 197636 159956
rect 197688 159944 197694 159996
rect 201034 159944 201040 159996
rect 201092 159984 201098 159996
rect 271874 159984 271880 159996
rect 201092 159956 271880 159984
rect 201092 159944 201098 159956
rect 271874 159944 271880 159956
rect 271932 159944 271938 159996
rect 274910 159944 274916 159996
rect 274968 159984 274974 159996
rect 324406 159984 324412 159996
rect 274968 159956 324412 159984
rect 274968 159944 274974 159956
rect 324406 159944 324412 159956
rect 324464 159944 324470 159996
rect 324498 159944 324504 159996
rect 324556 159984 324562 159996
rect 328362 159984 328368 159996
rect 324556 159956 328368 159984
rect 324556 159944 324562 159956
rect 328362 159944 328368 159956
rect 328420 159944 328426 159996
rect 328454 159944 328460 159996
rect 328512 159984 328518 159996
rect 331306 159984 331312 159996
rect 328512 159956 331312 159984
rect 328512 159944 328518 159956
rect 331306 159944 331312 159956
rect 331364 159944 331370 159996
rect 331416 159984 331444 160092
rect 331490 160012 331496 160064
rect 331548 160052 331554 160064
rect 334066 160052 334072 160064
rect 331548 160024 334072 160052
rect 331548 160012 331554 160024
rect 334066 160012 334072 160024
rect 334124 160012 334130 160064
rect 334618 160012 334624 160064
rect 334676 160052 334682 160064
rect 374730 160052 374736 160064
rect 334676 160024 374736 160052
rect 334676 160012 334682 160024
rect 374730 160012 374736 160024
rect 374788 160012 374794 160064
rect 381630 160012 381636 160064
rect 381688 160052 381694 160064
rect 398834 160052 398840 160064
rect 381688 160024 398840 160052
rect 381688 160012 381694 160024
rect 398834 160012 398840 160024
rect 398892 160012 398898 160064
rect 401778 160012 401784 160064
rect 401836 160052 401842 160064
rect 407574 160052 407580 160064
rect 401836 160024 407580 160052
rect 401836 160012 401842 160024
rect 407574 160012 407580 160024
rect 407632 160012 407638 160064
rect 426986 160012 426992 160064
rect 427044 160052 427050 160064
rect 445294 160052 445300 160064
rect 427044 160024 445300 160052
rect 427044 160012 427050 160024
rect 445294 160012 445300 160024
rect 445352 160012 445358 160064
rect 332594 159984 332600 159996
rect 331416 159956 332600 159984
rect 332594 159944 332600 159956
rect 332652 159944 332658 159996
rect 333698 159944 333704 159996
rect 333756 159984 333762 159996
rect 373994 159984 374000 159996
rect 333756 159956 374000 159984
rect 333756 159944 333762 159956
rect 373994 159944 374000 159956
rect 374052 159944 374058 159996
rect 374914 159944 374920 159996
rect 374972 159984 374978 159996
rect 397914 159984 397920 159996
rect 374972 159956 397920 159984
rect 374972 159944 374978 159956
rect 397914 159944 397920 159956
rect 397972 159944 397978 159996
rect 399202 159944 399208 159996
rect 399260 159984 399266 159996
rect 418246 159984 418252 159996
rect 399260 159956 418252 159984
rect 399260 159944 399266 159956
rect 418246 159944 418252 159956
rect 418304 159944 418310 159996
rect 424410 159944 424416 159996
rect 424468 159984 424474 159996
rect 443454 159984 443460 159996
rect 424468 159956 443460 159984
rect 424468 159944 424474 159956
rect 443454 159944 443460 159956
rect 443512 159944 443518 159996
rect 457990 159944 457996 159996
rect 458048 159984 458054 159996
rect 464890 159984 464896 159996
rect 458048 159956 464896 159984
rect 458048 159944 458054 159956
rect 464890 159944 464896 159956
rect 464948 159944 464954 159996
rect 466454 159944 466460 159996
rect 466512 159984 466518 159996
rect 473354 159984 473360 159996
rect 466512 159956 473360 159984
rect 466512 159944 466518 159956
rect 473354 159944 473360 159956
rect 473412 159944 473418 159996
rect 479058 159944 479064 159996
rect 479116 159984 479122 159996
rect 485222 159984 485228 159996
rect 479116 159956 485228 159984
rect 479116 159944 479122 159956
rect 485222 159944 485228 159956
rect 485280 159944 485286 159996
rect 49878 159876 49884 159928
rect 49936 159916 49942 159928
rect 133598 159916 133604 159928
rect 49936 159888 133604 159916
rect 49936 159876 49942 159888
rect 133598 159876 133604 159888
rect 133656 159876 133662 159928
rect 133690 159876 133696 159928
rect 133748 159916 133754 159928
rect 137094 159916 137100 159928
rect 133748 159888 137100 159916
rect 133748 159876 133754 159888
rect 137094 159876 137100 159888
rect 137152 159876 137158 159928
rect 137278 159876 137284 159928
rect 137336 159916 137342 159928
rect 142706 159916 142712 159928
rect 137336 159888 142712 159916
rect 137336 159876 137342 159888
rect 142706 159876 142712 159888
rect 142764 159876 142770 159928
rect 142798 159876 142804 159928
rect 142856 159916 142862 159928
rect 142856 159888 153148 159916
rect 142856 159876 142862 159888
rect 70026 159808 70032 159860
rect 70084 159848 70090 159860
rect 153010 159848 153016 159860
rect 70084 159820 153016 159848
rect 70084 159808 70090 159820
rect 153010 159808 153016 159820
rect 153068 159808 153074 159860
rect 153120 159848 153148 159888
rect 153194 159876 153200 159928
rect 153252 159916 153258 159928
rect 189718 159916 189724 159928
rect 153252 159888 189724 159916
rect 153252 159876 153258 159888
rect 189718 159876 189724 159888
rect 189776 159876 189782 159928
rect 194318 159876 194324 159928
rect 194376 159916 194382 159928
rect 267550 159916 267556 159928
rect 194376 159888 267556 159916
rect 194376 159876 194382 159888
rect 267550 159876 267556 159888
rect 267608 159876 267614 159928
rect 270770 159876 270776 159928
rect 270828 159916 270834 159928
rect 273346 159916 273352 159928
rect 270828 159888 273352 159916
rect 270828 159876 270834 159888
rect 273346 159876 273352 159888
rect 273404 159876 273410 159928
rect 274082 159876 274088 159928
rect 274140 159916 274146 159928
rect 328546 159916 328552 159928
rect 274140 159888 328552 159916
rect 274140 159876 274146 159888
rect 328546 159876 328552 159888
rect 328604 159876 328610 159928
rect 328730 159876 328736 159928
rect 328788 159916 328794 159928
rect 370038 159916 370044 159928
rect 328788 159888 370044 159916
rect 328788 159876 328794 159888
rect 370038 159876 370044 159888
rect 370096 159876 370102 159928
rect 374086 159876 374092 159928
rect 374144 159916 374150 159928
rect 380710 159916 380716 159928
rect 374144 159888 380716 159916
rect 374144 159876 374150 159888
rect 380710 159876 380716 159888
rect 380768 159876 380774 159928
rect 380802 159876 380808 159928
rect 380860 159916 380866 159928
rect 388622 159916 388628 159928
rect 380860 159888 388628 159916
rect 380860 159876 380866 159888
rect 388622 159876 388628 159888
rect 388680 159876 388686 159928
rect 389174 159876 389180 159928
rect 389232 159916 389238 159928
rect 415946 159916 415952 159928
rect 389232 159888 415952 159916
rect 389232 159876 389238 159888
rect 415946 159876 415952 159888
rect 416004 159876 416010 159928
rect 416038 159876 416044 159928
rect 416096 159916 416102 159928
rect 423398 159916 423404 159928
rect 416096 159888 423404 159916
rect 416096 159876 416102 159888
rect 423398 159876 423404 159888
rect 423456 159876 423462 159928
rect 423582 159876 423588 159928
rect 423640 159916 423646 159928
rect 442810 159916 442816 159928
rect 423640 159888 442816 159916
rect 423640 159876 423646 159888
rect 442810 159876 442816 159888
rect 442868 159876 442874 159928
rect 154390 159848 154396 159860
rect 153120 159820 154396 159848
rect 154390 159808 154396 159820
rect 154448 159808 154454 159860
rect 156506 159808 156512 159860
rect 156564 159848 156570 159860
rect 172422 159848 172428 159860
rect 156564 159820 172428 159848
rect 156564 159808 156570 159820
rect 172422 159808 172428 159820
rect 172480 159808 172486 159860
rect 176654 159808 176660 159860
rect 176712 159848 176718 159860
rect 181990 159848 181996 159860
rect 176712 159820 181996 159848
rect 176712 159808 176718 159820
rect 181990 159808 181996 159820
rect 182048 159808 182054 159860
rect 184290 159808 184296 159860
rect 184348 159848 184354 159860
rect 185026 159848 185032 159860
rect 184348 159820 185032 159848
rect 184348 159808 184354 159820
rect 185026 159808 185032 159820
rect 185084 159808 185090 159860
rect 255498 159848 255504 159860
rect 186286 159820 255504 159848
rect 59998 159740 60004 159792
rect 60056 159780 60062 159792
rect 149054 159780 149060 159792
rect 60056 159752 149060 159780
rect 60056 159740 60062 159752
rect 149054 159740 149060 159752
rect 149112 159740 149118 159792
rect 149790 159740 149796 159792
rect 149848 159780 149854 159792
rect 180794 159780 180800 159792
rect 149848 159752 180800 159780
rect 149848 159740 149854 159752
rect 180794 159740 180800 159752
rect 180852 159740 180858 159792
rect 180886 159740 180892 159792
rect 180944 159780 180950 159792
rect 186286 159780 186314 159820
rect 255498 159808 255504 159820
rect 255556 159808 255562 159860
rect 260650 159808 260656 159860
rect 260708 159848 260714 159860
rect 317138 159848 317144 159860
rect 260708 159820 317144 159848
rect 260708 159808 260714 159820
rect 317138 159808 317144 159820
rect 317196 159808 317202 159860
rect 317708 159820 319024 159848
rect 180944 159752 186314 159780
rect 180944 159740 180950 159752
rect 187602 159740 187608 159792
rect 187660 159780 187666 159792
rect 262214 159780 262220 159792
rect 187660 159752 262220 159780
rect 187660 159740 187666 159752
rect 262214 159740 262220 159752
rect 262272 159740 262278 159792
rect 267366 159740 267372 159792
rect 267424 159780 267430 159792
rect 317708 159780 317736 159820
rect 267424 159752 317736 159780
rect 267424 159740 267430 159752
rect 317782 159740 317788 159792
rect 317840 159780 317846 159792
rect 318886 159780 318892 159792
rect 317840 159752 318892 159780
rect 317840 159740 317846 159752
rect 318886 159740 318892 159752
rect 318944 159740 318950 159792
rect 318996 159780 319024 159820
rect 321094 159808 321100 159860
rect 321152 159848 321158 159860
rect 363230 159848 363236 159860
rect 321152 159820 363236 159848
rect 321152 159808 321158 159820
rect 363230 159808 363236 159820
rect 363288 159808 363294 159860
rect 364794 159808 364800 159860
rect 364852 159848 364858 159860
rect 395522 159848 395528 159860
rect 364852 159820 395528 159848
rect 364852 159808 364858 159820
rect 395522 159808 395528 159820
rect 395580 159808 395586 159860
rect 410150 159808 410156 159860
rect 410208 159848 410214 159860
rect 432506 159848 432512 159860
rect 410208 159820 432512 159848
rect 410208 159808 410214 159820
rect 432506 159808 432512 159820
rect 432564 159808 432570 159860
rect 450446 159808 450452 159860
rect 450504 159848 450510 159860
rect 456794 159848 456800 159860
rect 450504 159820 456800 159848
rect 450504 159808 450510 159820
rect 456794 159808 456800 159820
rect 456852 159808 456858 159860
rect 458910 159808 458916 159860
rect 458968 159848 458974 159860
rect 465350 159848 465356 159860
rect 458968 159820 465356 159848
rect 458968 159808 458974 159820
rect 465350 159808 465356 159820
rect 465408 159808 465414 159860
rect 467282 159808 467288 159860
rect 467340 159848 467346 159860
rect 473446 159848 473452 159860
rect 467340 159820 473452 159848
rect 467340 159808 467346 159820
rect 473446 159808 473452 159820
rect 473504 159808 473510 159860
rect 482370 159808 482376 159860
rect 482428 159848 482434 159860
rect 487338 159848 487344 159860
rect 482428 159820 487344 159848
rect 482428 159808 482434 159820
rect 487338 159808 487344 159820
rect 487396 159808 487402 159860
rect 321554 159780 321560 159792
rect 318996 159752 321560 159780
rect 321554 159740 321560 159752
rect 321612 159740 321618 159792
rect 326982 159740 326988 159792
rect 327040 159780 327046 159792
rect 368934 159780 368940 159792
rect 327040 159752 368940 159780
rect 327040 159740 327046 159752
rect 368934 159740 368940 159752
rect 368992 159740 368998 159792
rect 375742 159740 375748 159792
rect 375800 159780 375806 159792
rect 405826 159780 405832 159792
rect 375800 159752 405832 159780
rect 375800 159740 375806 159752
rect 405826 159740 405832 159752
rect 405884 159740 405890 159792
rect 406838 159740 406844 159792
rect 406896 159780 406902 159792
rect 429930 159780 429936 159792
rect 406896 159752 429936 159780
rect 406896 159740 406902 159752
rect 429930 159740 429936 159752
rect 429988 159740 429994 159792
rect 448790 159740 448796 159792
rect 448848 159780 448854 159792
rect 460198 159780 460204 159792
rect 448848 159752 460204 159780
rect 448848 159740 448854 159752
rect 460198 159740 460204 159752
rect 460256 159740 460262 159792
rect 53282 159672 53288 159724
rect 53340 159712 53346 159724
rect 137278 159712 137284 159724
rect 53340 159684 137284 159712
rect 53340 159672 53346 159684
rect 137278 159672 137284 159684
rect 137336 159672 137342 159724
rect 137370 159672 137376 159724
rect 137428 159712 137434 159724
rect 139302 159712 139308 159724
rect 137428 159684 139308 159712
rect 137428 159672 137434 159684
rect 139302 159672 139308 159684
rect 139360 159672 139366 159724
rect 139762 159672 139768 159724
rect 139820 159712 139826 159724
rect 158714 159712 158720 159724
rect 139820 159684 158720 159712
rect 139820 159672 139826 159684
rect 158714 159672 158720 159684
rect 158772 159672 158778 159724
rect 164142 159712 164148 159724
rect 160756 159684 164148 159712
rect 39850 159604 39856 159656
rect 39908 159644 39914 159656
rect 124030 159644 124036 159656
rect 39908 159616 124036 159644
rect 39908 159604 39914 159616
rect 124030 159604 124036 159616
rect 124088 159604 124094 159656
rect 127158 159604 127164 159656
rect 127216 159644 127222 159656
rect 136266 159644 136272 159656
rect 127216 159616 136272 159644
rect 127216 159604 127222 159616
rect 136266 159604 136272 159616
rect 136324 159604 136330 159656
rect 136358 159604 136364 159656
rect 136416 159644 136422 159656
rect 160756 159644 160784 159684
rect 164142 159672 164148 159684
rect 164200 159672 164206 159724
rect 167454 159672 167460 159724
rect 167512 159712 167518 159724
rect 242986 159712 242992 159724
rect 167512 159684 242992 159712
rect 167512 159672 167518 159684
rect 242986 159672 242992 159684
rect 243044 159672 243050 159724
rect 248046 159672 248052 159724
rect 248104 159712 248110 159724
rect 308490 159712 308496 159724
rect 248104 159684 308496 159712
rect 248104 159672 248110 159684
rect 308490 159672 308496 159684
rect 308548 159672 308554 159724
rect 315298 159672 315304 159724
rect 315356 159712 315362 159724
rect 351270 159712 351276 159724
rect 315356 159684 351276 159712
rect 315356 159672 315362 159684
rect 351270 159672 351276 159684
rect 351328 159672 351334 159724
rect 351362 159672 351368 159724
rect 351420 159712 351426 159724
rect 357802 159712 357808 159724
rect 351420 159684 357808 159712
rect 351420 159672 351426 159684
rect 357802 159672 357808 159684
rect 357860 159672 357866 159724
rect 369026 159672 369032 159724
rect 369084 159712 369090 159724
rect 401042 159712 401048 159724
rect 369084 159684 401048 159712
rect 369084 159672 369090 159684
rect 401042 159672 401048 159684
rect 401100 159672 401106 159724
rect 403434 159672 403440 159724
rect 403492 159712 403498 159724
rect 427354 159712 427360 159724
rect 403492 159684 427360 159712
rect 403492 159672 403498 159684
rect 427354 159672 427360 159684
rect 427412 159672 427418 159724
rect 447134 159672 447140 159724
rect 447192 159712 447198 159724
rect 458174 159712 458180 159724
rect 447192 159684 458180 159712
rect 447192 159672 447198 159684
rect 458174 159672 458180 159684
rect 458232 159672 458238 159724
rect 459738 159672 459744 159724
rect 459796 159712 459802 159724
rect 466546 159712 466552 159724
rect 459796 159684 466552 159712
rect 459796 159672 459802 159684
rect 466546 159672 466552 159684
rect 466604 159672 466610 159724
rect 472342 159672 472348 159724
rect 472400 159712 472406 159724
rect 479426 159712 479432 159724
rect 472400 159684 479432 159712
rect 472400 159672 472406 159684
rect 479426 159672 479432 159684
rect 479484 159672 479490 159724
rect 479886 159672 479892 159724
rect 479944 159712 479950 159724
rect 485958 159712 485964 159724
rect 479944 159684 485964 159712
rect 479944 159672 479950 159684
rect 485958 159672 485964 159684
rect 486016 159672 486022 159724
rect 136416 159616 160784 159644
rect 136416 159604 136422 159616
rect 163222 159604 163228 159656
rect 163280 159644 163286 159656
rect 174078 159644 174084 159656
rect 163280 159616 174084 159644
rect 163280 159604 163286 159616
rect 174078 159604 174084 159616
rect 174136 159604 174142 159656
rect 174170 159604 174176 159656
rect 174228 159644 174234 159656
rect 251174 159644 251180 159656
rect 174228 159616 251180 159644
rect 174228 159604 174234 159616
rect 251174 159604 251180 159616
rect 251232 159604 251238 159656
rect 254762 159604 254768 159656
rect 254820 159644 254826 159656
rect 313734 159644 313740 159656
rect 254820 159616 313740 159644
rect 254820 159604 254826 159616
rect 313734 159604 313740 159616
rect 313792 159604 313798 159656
rect 314378 159604 314384 159656
rect 314436 159644 314442 159656
rect 357526 159644 357532 159656
rect 314436 159616 357532 159644
rect 314436 159604 314442 159616
rect 357526 159604 357532 159616
rect 357584 159604 357590 159656
rect 357618 159604 357624 159656
rect 357676 159644 357682 159656
rect 358814 159644 358820 159656
rect 357676 159616 358820 159644
rect 357676 159604 357682 159616
rect 358814 159604 358820 159616
rect 358872 159604 358878 159656
rect 362310 159604 362316 159656
rect 362368 159644 362374 159656
rect 395246 159644 395252 159656
rect 362368 159616 395252 159644
rect 362368 159604 362374 159616
rect 395246 159604 395252 159616
rect 395304 159604 395310 159656
rect 407666 159604 407672 159656
rect 407724 159644 407730 159656
rect 430666 159644 430672 159656
rect 407724 159616 430672 159644
rect 407724 159604 407730 159616
rect 430666 159604 430672 159616
rect 430724 159604 430730 159656
rect 453850 159604 453856 159656
rect 453908 159644 453914 159656
rect 465074 159644 465080 159656
rect 453908 159616 465080 159644
rect 453908 159604 453914 159616
rect 465074 159604 465080 159616
rect 465132 159604 465138 159656
rect 470594 159604 470600 159656
rect 470652 159644 470658 159656
rect 477678 159644 477684 159656
rect 470652 159616 477684 159644
rect 470652 159604 470658 159616
rect 477678 159604 477684 159616
rect 477736 159604 477742 159656
rect 480714 159604 480720 159656
rect 480772 159644 480778 159656
rect 486510 159644 486516 159656
rect 480772 159616 486516 159644
rect 480772 159604 480778 159616
rect 486510 159604 486516 159616
rect 486568 159604 486574 159656
rect 22186 159536 22192 159588
rect 22244 159576 22250 159588
rect 127250 159576 127256 159588
rect 22244 159548 127256 159576
rect 22244 159536 22250 159548
rect 127250 159536 127256 159548
rect 127308 159536 127314 159588
rect 127618 159536 127624 159588
rect 127676 159576 127682 159588
rect 133690 159576 133696 159588
rect 127676 159548 133696 159576
rect 127676 159536 127682 159548
rect 133690 159536 133696 159548
rect 133748 159536 133754 159588
rect 133782 159536 133788 159588
rect 133840 159576 133846 159588
rect 139486 159576 139492 159588
rect 133840 159548 139492 159576
rect 133840 159536 133846 159548
rect 139486 159536 139492 159548
rect 139544 159536 139550 159588
rect 140590 159536 140596 159588
rect 140648 159576 140654 159588
rect 218146 159576 218152 159588
rect 140648 159548 218152 159576
rect 140648 159536 140654 159548
rect 218146 159536 218152 159548
rect 218204 159536 218210 159588
rect 221182 159536 221188 159588
rect 221240 159576 221246 159588
rect 221240 159548 287468 159576
rect 221240 159536 221246 159548
rect 28902 159468 28908 159520
rect 28960 159508 28966 159520
rect 132862 159508 132868 159520
rect 28960 159480 132868 159508
rect 28960 159468 28966 159480
rect 132862 159468 132868 159480
rect 132920 159468 132926 159520
rect 136542 159508 136548 159520
rect 132972 159480 136548 159508
rect 23014 159400 23020 159452
rect 23072 159440 23078 159452
rect 132972 159440 133000 159480
rect 136542 159468 136548 159480
rect 136600 159468 136606 159520
rect 137186 159468 137192 159520
rect 137244 159508 137250 159520
rect 142798 159508 142804 159520
rect 137244 159480 142804 159508
rect 137244 159468 137250 159480
rect 142798 159468 142804 159480
rect 142856 159468 142862 159520
rect 142982 159468 142988 159520
rect 143040 159508 143046 159520
rect 144454 159508 144460 159520
rect 143040 159480 144460 159508
rect 143040 159468 143046 159480
rect 144454 159468 144460 159480
rect 144512 159468 144518 159520
rect 147306 159468 147312 159520
rect 147364 159508 147370 159520
rect 226334 159508 226340 159520
rect 147364 159480 226340 159508
rect 147364 159468 147370 159480
rect 226334 159468 226340 159480
rect 226392 159468 226398 159520
rect 227898 159468 227904 159520
rect 227956 159508 227962 159520
rect 287330 159508 287336 159520
rect 227956 159480 287336 159508
rect 227956 159468 227962 159480
rect 287330 159468 287336 159480
rect 287388 159468 287394 159520
rect 287440 159508 287468 159548
rect 287514 159536 287520 159588
rect 287572 159576 287578 159588
rect 337010 159576 337016 159588
rect 287572 159548 337016 159576
rect 287572 159536 287578 159548
rect 337010 159536 337016 159548
rect 337068 159536 337074 159588
rect 337856 159548 339724 159576
rect 288066 159508 288072 159520
rect 287440 159480 288072 159508
rect 288066 159468 288072 159480
rect 288124 159468 288130 159520
rect 291654 159468 291660 159520
rect 291712 159508 291718 159520
rect 295058 159508 295064 159520
rect 291712 159480 295064 159508
rect 291712 159468 291718 159480
rect 295058 159468 295064 159480
rect 295116 159468 295122 159520
rect 295150 159468 295156 159520
rect 295208 159508 295214 159520
rect 337856 159508 337884 159548
rect 295208 159480 337884 159508
rect 295208 159468 295214 159480
rect 337930 159468 337936 159520
rect 337988 159508 337994 159520
rect 339494 159508 339500 159520
rect 337988 159480 339500 159508
rect 337988 159468 337994 159480
rect 339494 159468 339500 159480
rect 339552 159468 339558 159520
rect 339696 159508 339724 159548
rect 342162 159536 342168 159588
rect 342220 159576 342226 159588
rect 380526 159576 380532 159588
rect 342220 159548 380532 159576
rect 342220 159536 342226 159548
rect 380526 159536 380532 159548
rect 380584 159536 380590 159588
rect 380710 159536 380716 159588
rect 380768 159576 380774 159588
rect 380768 159548 382964 159576
rect 380768 159536 380774 159548
rect 344554 159508 344560 159520
rect 339696 159480 344560 159508
rect 344554 159468 344560 159480
rect 344612 159468 344618 159520
rect 344646 159468 344652 159520
rect 344704 159508 344710 159520
rect 382550 159508 382556 159520
rect 344704 159480 382556 159508
rect 344704 159468 344710 159480
rect 382550 159468 382556 159480
rect 382608 159468 382614 159520
rect 382936 159508 382964 159548
rect 385770 159536 385776 159588
rect 385828 159576 385834 159588
rect 413186 159576 413192 159588
rect 385828 159548 413192 159576
rect 385828 159536 385834 159548
rect 413186 159536 413192 159548
rect 413244 159536 413250 159588
rect 416866 159536 416872 159588
rect 416924 159576 416930 159588
rect 437658 159576 437664 159588
rect 416924 159548 437664 159576
rect 416924 159536 416930 159548
rect 437658 159536 437664 159548
rect 437716 159536 437722 159588
rect 451274 159536 451280 159588
rect 451332 159576 451338 159588
rect 463694 159576 463700 159588
rect 451332 159548 463700 159576
rect 451332 159536 451338 159548
rect 463694 159536 463700 159548
rect 463752 159536 463758 159588
rect 469766 159536 469772 159588
rect 469824 159576 469830 159588
rect 476114 159576 476120 159588
rect 469824 159548 476120 159576
rect 469824 159536 469830 159548
rect 476114 159536 476120 159548
rect 476172 159536 476178 159588
rect 478138 159536 478144 159588
rect 478196 159576 478202 159588
rect 484578 159576 484584 159588
rect 478196 159548 484584 159576
rect 478196 159536 478202 159548
rect 484578 159536 484584 159548
rect 484636 159536 484642 159588
rect 388714 159508 388720 159520
rect 382936 159480 388720 159508
rect 388714 159468 388720 159480
rect 388772 159468 388778 159520
rect 413554 159468 413560 159520
rect 413612 159508 413618 159520
rect 435082 159508 435088 159520
rect 413612 159480 435088 159508
rect 413612 159468 413618 159480
rect 435082 159468 435088 159480
rect 435140 159468 435146 159520
rect 454678 159468 454684 159520
rect 454736 159508 454742 159520
rect 466638 159508 466644 159520
rect 454736 159480 466644 159508
rect 454736 159468 454742 159480
rect 466638 159468 466644 159480
rect 466696 159468 466702 159520
rect 484026 159468 484032 159520
rect 484084 159508 484090 159520
rect 488994 159508 489000 159520
rect 484084 159480 489000 159508
rect 484084 159468 484090 159480
rect 488994 159468 489000 159480
rect 489052 159468 489058 159520
rect 23072 159412 133000 159440
rect 23072 159400 23078 159412
rect 133046 159400 133052 159452
rect 133104 159440 133110 159452
rect 156598 159440 156604 159452
rect 133104 159412 156604 159440
rect 133104 159400 133110 159412
rect 156598 159400 156604 159412
rect 156656 159400 156662 159452
rect 160738 159400 160744 159452
rect 160796 159440 160802 159452
rect 240318 159440 240324 159452
rect 160796 159412 240324 159440
rect 160796 159400 160802 159412
rect 240318 159400 240324 159412
rect 240376 159400 240382 159452
rect 247218 159400 247224 159452
rect 247276 159440 247282 159452
rect 307754 159440 307760 159452
rect 247276 159412 307760 159440
rect 247276 159400 247282 159412
rect 307754 159400 307760 159412
rect 307812 159400 307818 159452
rect 308582 159400 308588 159452
rect 308640 159440 308646 159452
rect 349798 159440 349804 159452
rect 308640 159412 349804 159440
rect 308640 159400 308646 159412
rect 349798 159400 349804 159412
rect 349856 159400 349862 159452
rect 349890 159400 349896 159452
rect 349948 159440 349954 159452
rect 354214 159440 354220 159452
rect 349948 159412 354220 159440
rect 349948 159400 349954 159412
rect 354214 159400 354220 159412
rect 354272 159400 354278 159452
rect 357618 159440 357624 159452
rect 354324 159412 357624 159440
rect 2866 159332 2872 159384
rect 2924 159372 2930 159384
rect 116118 159372 116124 159384
rect 2924 159344 116124 159372
rect 2924 159332 2930 159344
rect 116118 159332 116124 159344
rect 116176 159332 116182 159384
rect 116210 159332 116216 159384
rect 116268 159372 116274 159384
rect 127618 159372 127624 159384
rect 116268 159344 127624 159372
rect 116268 159332 116274 159344
rect 127618 159332 127624 159344
rect 127676 159332 127682 159384
rect 129642 159332 129648 159384
rect 129700 159372 129706 159384
rect 142890 159372 142896 159384
rect 129700 159344 142896 159372
rect 129700 159332 129706 159344
rect 142890 159332 142896 159344
rect 142948 159332 142954 159384
rect 142982 159332 142988 159384
rect 143040 159372 143046 159384
rect 147122 159372 147128 159384
rect 143040 159344 147128 159372
rect 143040 159332 143046 159344
rect 147122 159332 147128 159344
rect 147180 159332 147186 159384
rect 150618 159332 150624 159384
rect 150676 159372 150682 159384
rect 152734 159372 152740 159384
rect 150676 159344 152740 159372
rect 150676 159332 150682 159344
rect 152734 159332 152740 159344
rect 152792 159332 152798 159384
rect 154022 159332 154028 159384
rect 154080 159372 154086 159384
rect 236730 159372 236736 159384
rect 154080 159344 236736 159372
rect 154080 159332 154086 159344
rect 236730 159332 236736 159344
rect 236788 159332 236794 159384
rect 241330 159332 241336 159384
rect 241388 159372 241394 159384
rect 303430 159372 303436 159384
rect 241388 159344 303436 159372
rect 241388 159332 241394 159344
rect 303430 159332 303436 159344
rect 303488 159332 303494 159384
rect 307662 159332 307668 159384
rect 307720 159372 307726 159384
rect 348786 159372 348792 159384
rect 307720 159344 348792 159372
rect 307720 159332 307726 159344
rect 348786 159332 348792 159344
rect 348844 159332 348850 159384
rect 348878 159332 348884 159384
rect 348936 159372 348942 159384
rect 348936 159344 350534 159372
rect 348936 159332 348942 159344
rect 83458 159264 83464 159316
rect 83516 159304 83522 159316
rect 166994 159304 167000 159316
rect 83516 159276 167000 159304
rect 83516 159264 83522 159276
rect 166994 159264 167000 159276
rect 167052 159264 167058 159316
rect 169938 159264 169944 159316
rect 169996 159304 170002 159316
rect 195330 159304 195336 159316
rect 169996 159276 195336 159304
rect 169996 159264 170002 159276
rect 195330 159264 195336 159276
rect 195388 159264 195394 159316
rect 197722 159264 197728 159316
rect 197780 159304 197786 159316
rect 214374 159304 214380 159316
rect 197780 159276 214380 159304
rect 197780 159264 197786 159276
rect 214374 159264 214380 159276
rect 214432 159264 214438 159316
rect 214466 159264 214472 159316
rect 214524 159304 214530 159316
rect 282822 159304 282828 159316
rect 214524 159276 282828 159304
rect 214524 159264 214530 159276
rect 282822 159264 282828 159276
rect 282880 159264 282886 159316
rect 287330 159264 287336 159316
rect 287388 159304 287394 159316
rect 293218 159304 293224 159316
rect 287388 159276 293224 159304
rect 287388 159264 287394 159276
rect 293218 159264 293224 159276
rect 293276 159264 293282 159316
rect 294230 159264 294236 159316
rect 294288 159304 294294 159316
rect 343634 159304 343640 159316
rect 294288 159276 343640 159304
rect 294288 159264 294294 159276
rect 343634 159264 343640 159276
rect 343692 159264 343698 159316
rect 343818 159264 343824 159316
rect 343876 159304 343882 159316
rect 349982 159304 349988 159316
rect 343876 159276 349988 159304
rect 343876 159264 343882 159276
rect 349982 159264 349988 159276
rect 350040 159264 350046 159316
rect 350506 159304 350534 159344
rect 351270 159332 351276 159384
rect 351328 159372 351334 159384
rect 354324 159372 354352 159412
rect 357618 159400 357624 159412
rect 357676 159400 357682 159452
rect 358078 159400 358084 159452
rect 358136 159440 358142 159452
rect 392394 159440 392400 159452
rect 358136 159412 392400 159440
rect 358136 159400 358142 159412
rect 392394 159400 392400 159412
rect 392452 159400 392458 159452
rect 395062 159400 395068 159452
rect 395120 159440 395126 159452
rect 405642 159440 405648 159452
rect 395120 159412 405648 159440
rect 395120 159400 395126 159412
rect 405642 159400 405648 159412
rect 405700 159400 405706 159452
rect 420270 159400 420276 159452
rect 420328 159440 420334 159452
rect 440326 159440 440332 159452
rect 420328 159412 440332 159440
rect 420328 159400 420334 159412
rect 440326 159400 440332 159412
rect 440384 159400 440390 159452
rect 452102 159400 452108 159452
rect 452160 159440 452166 159452
rect 464246 159440 464252 159452
rect 452160 159412 464252 159440
rect 452160 159400 452166 159412
rect 464246 159400 464252 159412
rect 464304 159400 464310 159452
rect 468938 159400 468944 159452
rect 468996 159440 469002 159452
rect 475010 159440 475016 159452
rect 468996 159412 475016 159440
rect 468996 159400 469002 159412
rect 475010 159400 475016 159412
rect 475068 159400 475074 159452
rect 476482 159400 476488 159452
rect 476540 159440 476546 159452
rect 483290 159440 483296 159452
rect 476540 159412 483296 159440
rect 476540 159400 476546 159412
rect 483290 159400 483296 159412
rect 483348 159400 483354 159452
rect 518802 159400 518808 159452
rect 518860 159440 518866 159452
rect 521838 159440 521844 159452
rect 518860 159412 521844 159440
rect 518860 159400 518866 159412
rect 521838 159400 521844 159412
rect 521896 159400 521902 159452
rect 351328 159344 354352 159372
rect 351328 159332 351334 159344
rect 355594 159332 355600 159384
rect 355652 159372 355658 159384
rect 390738 159372 390744 159384
rect 355652 159344 390744 159372
rect 355652 159332 355658 159344
rect 390738 159332 390744 159344
rect 390796 159332 390802 159384
rect 404262 159332 404268 159384
rect 404320 159372 404326 159384
rect 427998 159372 428004 159384
rect 404320 159344 428004 159372
rect 404320 159332 404326 159344
rect 427998 159332 428004 159344
rect 428056 159332 428062 159384
rect 446030 159372 446036 159384
rect 431926 159344 446036 159372
rect 385586 159304 385592 159316
rect 350506 159276 385592 159304
rect 385586 159264 385592 159276
rect 385644 159264 385650 159316
rect 388346 159264 388352 159316
rect 388404 159304 388410 159316
rect 401594 159304 401600 159316
rect 388404 159276 401600 159304
rect 388404 159264 388410 159276
rect 401594 159264 401600 159276
rect 401652 159264 401658 159316
rect 427814 159264 427820 159316
rect 427872 159304 427878 159316
rect 431926 159304 431954 159344
rect 446030 159332 446036 159344
rect 446088 159332 446094 159384
rect 453022 159332 453028 159384
rect 453080 159372 453086 159384
rect 465258 159372 465264 159384
rect 453080 159344 465264 159372
rect 453080 159332 453086 159344
rect 465258 159332 465264 159344
rect 465316 159332 465322 159384
rect 468110 159332 468116 159384
rect 468168 159372 468174 159384
rect 474734 159372 474740 159384
rect 468168 159344 474740 159372
rect 468168 159332 468174 159344
rect 474734 159332 474740 159344
rect 474792 159332 474798 159384
rect 477310 159332 477316 159384
rect 477368 159372 477374 159384
rect 483106 159372 483112 159384
rect 477368 159344 483112 159372
rect 477368 159332 477374 159344
rect 483106 159332 483112 159344
rect 483164 159332 483170 159384
rect 518710 159332 518716 159384
rect 518768 159372 518774 159384
rect 522666 159372 522672 159384
rect 518768 159344 522672 159372
rect 518768 159332 518774 159344
rect 522666 159332 522672 159344
rect 522724 159332 522730 159384
rect 427872 159276 431954 159304
rect 427872 159264 427878 159276
rect 90174 159196 90180 159248
rect 90232 159236 90238 159248
rect 173250 159236 173256 159248
rect 90232 159208 173256 159236
rect 90232 159196 90238 159208
rect 173250 159196 173256 159208
rect 173308 159196 173314 159248
rect 173342 159196 173348 159248
rect 173400 159236 173406 159248
rect 195238 159236 195244 159248
rect 173400 159208 195244 159236
rect 173400 159196 173406 159208
rect 195238 159196 195244 159208
rect 195296 159196 195302 159248
rect 196894 159196 196900 159248
rect 196952 159236 196958 159248
rect 211798 159236 211804 159248
rect 196952 159208 211804 159236
rect 196952 159196 196958 159208
rect 211798 159196 211804 159208
rect 211856 159196 211862 159248
rect 213638 159196 213644 159248
rect 213696 159236 213702 159248
rect 279786 159236 279792 159248
rect 213696 159208 279792 159236
rect 213696 159196 213702 159208
rect 279786 159196 279792 159208
rect 279844 159196 279850 159248
rect 281626 159196 281632 159248
rect 281684 159236 281690 159248
rect 328454 159236 328460 159248
rect 281684 159208 328460 159236
rect 281684 159196 281690 159208
rect 328454 159196 328460 159208
rect 328512 159196 328518 159248
rect 332042 159196 332048 159248
rect 332100 159236 332106 159248
rect 334526 159236 334532 159248
rect 332100 159208 334532 159236
rect 332100 159196 332106 159208
rect 334526 159196 334532 159208
rect 334584 159196 334590 159248
rect 335446 159196 335452 159248
rect 335504 159236 335510 159248
rect 375374 159236 375380 159248
rect 335504 159208 375380 159236
rect 335504 159196 335510 159208
rect 375374 159196 375380 159208
rect 375432 159196 375438 159248
rect 391658 159196 391664 159248
rect 391716 159236 391722 159248
rect 403894 159236 403900 159248
rect 391716 159208 403900 159236
rect 391716 159196 391722 159208
rect 403894 159196 403900 159208
rect 403952 159196 403958 159248
rect 457162 159196 457168 159248
rect 457220 159236 457226 159248
rect 464614 159236 464620 159248
rect 457220 159208 464620 159236
rect 457220 159196 457226 159208
rect 464614 159196 464620 159208
rect 464672 159196 464678 159248
rect 63310 159128 63316 159180
rect 63368 159168 63374 159180
rect 102134 159168 102140 159180
rect 63368 159140 102140 159168
rect 63368 159128 63374 159140
rect 102134 159128 102140 159140
rect 102192 159128 102198 159180
rect 103606 159128 103612 159180
rect 103664 159168 103670 159180
rect 183094 159168 183100 159180
rect 103664 159140 183100 159168
rect 103664 159128 103670 159140
rect 183094 159128 183100 159140
rect 183152 159128 183158 159180
rect 193490 159128 193496 159180
rect 193548 159168 193554 159180
rect 223574 159168 223580 159180
rect 193548 159140 223580 159168
rect 193548 159128 193554 159140
rect 223574 159128 223580 159140
rect 223632 159128 223638 159180
rect 234614 159128 234620 159180
rect 234672 159168 234678 159180
rect 298370 159168 298376 159180
rect 234672 159140 298376 159168
rect 234672 159128 234678 159140
rect 298370 159128 298376 159140
rect 298428 159128 298434 159180
rect 301866 159128 301872 159180
rect 301924 159168 301930 159180
rect 349706 159168 349712 159180
rect 301924 159140 349712 159168
rect 301924 159128 301930 159140
rect 349706 159128 349712 159140
rect 349764 159128 349770 159180
rect 353294 159168 353300 159180
rect 349908 159140 353300 159168
rect 80146 159060 80152 159112
rect 80204 159100 80210 159112
rect 89714 159100 89720 159112
rect 80204 159072 89720 159100
rect 80204 159060 80210 159072
rect 89714 159060 89720 159072
rect 89772 159060 89778 159112
rect 96890 159060 96896 159112
rect 96948 159100 96954 159112
rect 173986 159100 173992 159112
rect 96948 159072 173992 159100
rect 96948 159060 96954 159072
rect 173986 159060 173992 159072
rect 174044 159060 174050 159112
rect 174078 159060 174084 159112
rect 174136 159100 174142 159112
rect 179046 159100 179052 159112
rect 174136 159072 179052 159100
rect 174136 159060 174142 159072
rect 179046 159060 179052 159072
rect 179104 159060 179110 159112
rect 180794 159060 180800 159112
rect 180852 159100 180858 159112
rect 181622 159100 181628 159112
rect 180852 159072 181628 159100
rect 180852 159060 180858 159072
rect 181622 159060 181628 159072
rect 181680 159060 181686 159112
rect 186774 159060 186780 159112
rect 186832 159100 186838 159112
rect 214558 159100 214564 159112
rect 186832 159072 214564 159100
rect 186832 159060 186838 159072
rect 214558 159060 214564 159072
rect 214616 159060 214622 159112
rect 220354 159060 220360 159112
rect 220412 159100 220418 159112
rect 229370 159100 229376 159112
rect 220412 159072 229376 159100
rect 220412 159060 220418 159072
rect 229370 159060 229376 159072
rect 229428 159060 229434 159112
rect 230474 159060 230480 159112
rect 230532 159100 230538 159112
rect 294506 159100 294512 159112
rect 230532 159072 294512 159100
rect 230532 159060 230538 159072
rect 294506 159060 294512 159072
rect 294564 159060 294570 159112
rect 300946 159060 300952 159112
rect 301004 159100 301010 159112
rect 349062 159100 349068 159112
rect 301004 159072 349068 159100
rect 301004 159060 301010 159072
rect 349062 159060 349068 159072
rect 349120 159060 349126 159112
rect 92750 158992 92756 159044
rect 92808 159032 92814 159044
rect 116026 159032 116032 159044
rect 92808 159004 116032 159032
rect 92808 158992 92814 159004
rect 116026 158992 116032 159004
rect 116084 158992 116090 159044
rect 116118 158992 116124 159044
rect 116176 159032 116182 159044
rect 118694 159032 118700 159044
rect 116176 159004 118700 159032
rect 116176 158992 116182 159004
rect 118694 158992 118700 159004
rect 118752 158992 118758 159044
rect 119614 158992 119620 159044
rect 119672 159032 119678 159044
rect 133782 159032 133788 159044
rect 119672 159004 133788 159032
rect 119672 158992 119678 159004
rect 133782 158992 133788 159004
rect 133840 158992 133846 159044
rect 133874 158992 133880 159044
rect 133932 159032 133938 159044
rect 210234 159032 210240 159044
rect 133932 159004 210240 159032
rect 133932 158992 133938 159004
rect 210234 158992 210240 159004
rect 210292 158992 210298 159044
rect 210326 158992 210332 159044
rect 210384 159032 210390 159044
rect 214006 159032 214012 159044
rect 210384 159004 214012 159032
rect 210384 158992 210390 159004
rect 214006 158992 214012 159004
rect 214064 158992 214070 159044
rect 214374 158992 214380 159044
rect 214432 159032 214438 159044
rect 215386 159032 215392 159044
rect 214432 159004 215392 159032
rect 214432 158992 214438 159004
rect 215386 158992 215392 159004
rect 215444 158992 215450 159044
rect 224218 158992 224224 159044
rect 224276 159032 224282 159044
rect 227714 159032 227720 159044
rect 224276 159004 227720 159032
rect 224276 158992 224282 159004
rect 227714 158992 227720 159004
rect 227772 158992 227778 159044
rect 233786 158992 233792 159044
rect 233844 159032 233850 159044
rect 291654 159032 291660 159044
rect 233844 159004 291660 159032
rect 233844 158992 233850 159004
rect 291654 158992 291660 159004
rect 291712 158992 291718 159044
rect 291746 158992 291752 159044
rect 291804 159032 291810 159044
rect 293954 159032 293960 159044
rect 291804 159004 293960 159032
rect 291804 158992 291810 159004
rect 293954 158992 293960 159004
rect 294012 158992 294018 159044
rect 298462 158992 298468 159044
rect 298520 159032 298526 159044
rect 299474 159032 299480 159044
rect 298520 159004 299480 159032
rect 298520 158992 298526 159004
rect 299474 158992 299480 159004
rect 299532 158992 299538 159044
rect 306834 158992 306840 159044
rect 306892 159032 306898 159044
rect 349908 159032 349936 159140
rect 353294 159128 353300 159140
rect 353352 159128 353358 159180
rect 353846 159128 353852 159180
rect 353904 159168 353910 159180
rect 357710 159168 357716 159180
rect 353904 159140 357716 159168
rect 353904 159128 353910 159140
rect 357710 159128 357716 159140
rect 357768 159128 357774 159180
rect 357802 159128 357808 159180
rect 357860 159168 357866 159180
rect 387610 159168 387616 159180
rect 357860 159140 387616 159168
rect 357860 159128 357866 159140
rect 387610 159128 387616 159140
rect 387668 159128 387674 159180
rect 392486 159128 392492 159180
rect 392544 159168 392550 159180
rect 415670 159168 415676 159180
rect 392544 159140 415676 159168
rect 392544 159128 392550 159140
rect 415670 159128 415676 159140
rect 415728 159128 415734 159180
rect 461394 159128 461400 159180
rect 461452 159168 461458 159180
rect 468018 159168 468024 159180
rect 461452 159140 468024 159168
rect 461452 159128 461458 159140
rect 468018 159128 468024 159140
rect 468076 159128 468082 159180
rect 349982 159060 349988 159112
rect 350040 159100 350046 159112
rect 377766 159100 377772 159112
rect 350040 159072 377772 159100
rect 350040 159060 350046 159072
rect 377766 159060 377772 159072
rect 377824 159060 377830 159112
rect 380894 159100 380900 159112
rect 378704 159072 380900 159100
rect 306892 159004 349936 159032
rect 306892 158992 306898 159004
rect 350074 158992 350080 159044
rect 350132 159032 350138 159044
rect 354858 159032 354864 159044
rect 350132 159004 354864 159032
rect 350132 158992 350138 159004
rect 354858 158992 354864 159004
rect 354916 158992 354922 159044
rect 357618 159032 357624 159044
rect 354968 159004 357624 159032
rect 113634 158924 113640 158976
rect 113692 158964 113698 158976
rect 120074 158964 120080 158976
rect 113692 158936 120080 158964
rect 113692 158924 113698 158936
rect 120074 158924 120080 158936
rect 120132 158924 120138 158976
rect 120442 158924 120448 158976
rect 120500 158964 120506 158976
rect 120500 158936 122696 158964
rect 120500 158924 120506 158936
rect 106182 158856 106188 158908
rect 106240 158896 106246 158908
rect 122558 158896 122564 158908
rect 106240 158868 122564 158896
rect 106240 158856 106246 158868
rect 122558 158856 122564 158868
rect 122616 158856 122622 158908
rect 122668 158896 122696 158936
rect 122742 158924 122748 158976
rect 122800 158964 122806 158976
rect 186406 158964 186412 158976
rect 122800 158936 186412 158964
rect 122800 158924 122806 158936
rect 186406 158924 186412 158936
rect 186464 158924 186470 158976
rect 195238 158924 195244 158976
rect 195296 158964 195302 158976
rect 195296 158936 200804 158964
rect 195296 158924 195302 158936
rect 194502 158896 194508 158908
rect 122668 158868 194508 158896
rect 194502 158856 194508 158868
rect 194560 158856 194566 158908
rect 195330 158856 195336 158908
rect 195388 158896 195394 158908
rect 198734 158896 198740 158908
rect 195388 158868 198740 158896
rect 195388 158856 195394 158868
rect 198734 158856 198740 158868
rect 198792 158856 198798 158908
rect 200776 158896 200804 158936
rect 203610 158924 203616 158976
rect 203668 158964 203674 158976
rect 233142 158964 233148 158976
rect 203668 158936 233148 158964
rect 203668 158924 203674 158936
rect 233142 158924 233148 158936
rect 233200 158924 233206 158976
rect 240502 158924 240508 158976
rect 240560 158964 240566 158976
rect 300854 158964 300860 158976
rect 240560 158936 300860 158964
rect 240560 158924 240566 158936
rect 300854 158924 300860 158936
rect 300912 158924 300918 158976
rect 310238 158924 310244 158976
rect 310296 158964 310302 158976
rect 310698 158964 310704 158976
rect 310296 158936 310704 158964
rect 310296 158924 310302 158936
rect 310698 158924 310704 158936
rect 310756 158924 310762 158976
rect 313550 158924 313556 158976
rect 313608 158964 313614 158976
rect 354968 158964 354996 159004
rect 357618 158992 357624 159004
rect 357676 158992 357682 159044
rect 357710 158992 357716 159044
rect 357768 159032 357774 159044
rect 378704 159032 378732 159072
rect 380894 159060 380900 159072
rect 380952 159060 380958 159112
rect 390830 159060 390836 159112
rect 390888 159100 390894 159112
rect 391934 159100 391940 159112
rect 390888 159072 391940 159100
rect 390888 159060 390894 159072
rect 391934 159060 391940 159072
rect 391992 159060 391998 159112
rect 422754 159060 422760 159112
rect 422812 159100 422818 159112
rect 424962 159100 424968 159112
rect 422812 159072 424968 159100
rect 422812 159060 422818 159072
rect 424962 159060 424968 159072
rect 425020 159060 425026 159112
rect 460566 159060 460572 159112
rect 460624 159100 460630 159112
rect 466454 159100 466460 159112
rect 460624 159072 466460 159100
rect 460624 159060 460630 159072
rect 466454 159060 466460 159072
rect 466512 159060 466518 159112
rect 473170 159060 473176 159112
rect 473228 159100 473234 159112
rect 478874 159100 478880 159112
rect 473228 159072 478880 159100
rect 473228 159060 473234 159072
rect 478874 159060 478880 159072
rect 478932 159060 478938 159112
rect 481542 159060 481548 159112
rect 481600 159100 481606 159112
rect 487246 159100 487252 159112
rect 481600 159072 487252 159100
rect 481600 159060 481606 159072
rect 487246 159060 487252 159072
rect 487304 159060 487310 159112
rect 357768 159004 378732 159032
rect 378888 159004 379514 159032
rect 357768 158992 357774 159004
rect 365162 158964 365168 158976
rect 313608 158936 354996 158964
rect 355244 158936 365168 158964
rect 313608 158924 313614 158936
rect 204070 158896 204076 158908
rect 200776 158868 204076 158896
rect 204070 158856 204076 158868
rect 204128 158856 204134 158908
rect 206922 158856 206928 158908
rect 206980 158896 206986 158908
rect 233878 158896 233884 158908
rect 206980 158868 233884 158896
rect 206980 158856 206986 158868
rect 233878 158856 233884 158868
rect 233936 158856 233942 158908
rect 253934 158856 253940 158908
rect 253992 158896 253998 158908
rect 311986 158896 311992 158908
rect 253992 158868 311992 158896
rect 253992 158856 253998 158868
rect 311986 158856 311992 158868
rect 312044 158856 312050 158908
rect 318610 158856 318616 158908
rect 318668 158896 318674 158908
rect 319162 158896 319168 158908
rect 318668 158868 319168 158896
rect 318668 158856 318674 158868
rect 319162 158856 319168 158868
rect 319220 158856 319226 158908
rect 324038 158896 324044 158908
rect 320008 158868 324044 158896
rect 102778 158788 102784 158840
rect 102836 158828 102842 158840
rect 123938 158828 123944 158840
rect 102836 158800 123944 158828
rect 102836 158788 102842 158800
rect 123938 158788 123944 158800
rect 123996 158788 124002 158840
rect 124030 158788 124036 158840
rect 124088 158828 124094 158840
rect 135162 158828 135168 158840
rect 124088 158800 135168 158828
rect 124088 158788 124094 158800
rect 135162 158788 135168 158800
rect 135220 158788 135226 158840
rect 136266 158788 136272 158840
rect 136324 158828 136330 158840
rect 196066 158828 196072 158840
rect 136324 158800 196072 158828
rect 136324 158788 136330 158800
rect 196066 158788 196072 158800
rect 196124 158788 196130 158840
rect 200206 158788 200212 158840
rect 200264 158828 200270 158840
rect 224218 158828 224224 158840
rect 200264 158800 224224 158828
rect 200264 158788 200270 158800
rect 224218 158788 224224 158800
rect 224276 158788 224282 158840
rect 224586 158788 224592 158840
rect 224644 158828 224650 158840
rect 230750 158828 230756 158840
rect 224644 158800 230756 158828
rect 224644 158788 224650 158800
rect 230750 158788 230756 158800
rect 230808 158788 230814 158840
rect 243906 158788 243912 158840
rect 243964 158828 243970 158840
rect 246114 158828 246120 158840
rect 243964 158800 246120 158828
rect 243964 158788 243970 158800
rect 246114 158788 246120 158800
rect 246172 158788 246178 158840
rect 261478 158788 261484 158840
rect 261536 158828 261542 158840
rect 318702 158828 318708 158840
rect 261536 158800 318708 158828
rect 261536 158788 261542 158800
rect 318702 158788 318708 158800
rect 318760 158788 318766 158840
rect 99466 158720 99472 158772
rect 99524 158760 99530 158772
rect 113634 158760 113640 158772
rect 99524 158732 113640 158760
rect 99524 158720 99530 158732
rect 113634 158720 113640 158732
rect 113692 158720 113698 158772
rect 113726 158720 113732 158772
rect 113784 158760 113790 158772
rect 122742 158760 122748 158772
rect 113784 158732 122748 158760
rect 113784 158720 113790 158732
rect 122742 158720 122748 158732
rect 122800 158720 122806 158772
rect 122926 158720 122932 158772
rect 122984 158760 122990 158772
rect 142982 158760 142988 158772
rect 122984 158732 142988 158760
rect 122984 158720 122990 158732
rect 142982 158720 142988 158732
rect 143040 158720 143046 158772
rect 143074 158720 143080 158772
rect 143132 158760 143138 158772
rect 176470 158760 176476 158772
rect 143132 158732 176476 158760
rect 143132 158720 143138 158732
rect 176470 158720 176476 158732
rect 176528 158720 176534 158772
rect 180058 158720 180064 158772
rect 180116 158760 180122 158772
rect 202874 158760 202880 158772
rect 180116 158732 202880 158760
rect 180116 158720 180122 158732
rect 202874 158720 202880 158732
rect 202932 158720 202938 158772
rect 204438 158720 204444 158772
rect 204496 158760 204502 158772
rect 219894 158760 219900 158772
rect 204496 158732 219900 158760
rect 204496 158720 204502 158732
rect 219894 158720 219900 158732
rect 219952 158720 219958 158772
rect 227070 158720 227076 158772
rect 227128 158760 227134 158772
rect 241422 158760 241428 158772
rect 227128 158732 241428 158760
rect 227128 158720 227134 158732
rect 241422 158720 241428 158732
rect 241480 158720 241486 158772
rect 244734 158720 244740 158772
rect 244792 158760 244798 158772
rect 245746 158760 245752 158772
rect 244792 158732 245752 158760
rect 244792 158720 244798 158732
rect 245746 158720 245752 158732
rect 245804 158720 245810 158772
rect 251450 158720 251456 158772
rect 251508 158760 251514 158772
rect 252922 158760 252928 158772
rect 251508 158732 252928 158760
rect 251508 158720 251514 158732
rect 252922 158720 252928 158732
rect 252980 158720 252986 158772
rect 268194 158720 268200 158772
rect 268252 158760 268258 158772
rect 320008 158760 320036 158868
rect 324038 158856 324044 158868
rect 324096 158856 324102 158908
rect 324406 158856 324412 158908
rect 324464 158896 324470 158908
rect 328454 158896 328460 158908
rect 324464 158868 328460 158896
rect 324464 158856 324470 158868
rect 328454 158856 328460 158868
rect 328512 158856 328518 158908
rect 328638 158856 328644 158908
rect 328696 158896 328702 158908
rect 355244 158896 355272 158936
rect 365162 158924 365168 158936
rect 365220 158924 365226 158976
rect 371510 158924 371516 158976
rect 371568 158964 371574 158976
rect 378888 158964 378916 159004
rect 371568 158936 378916 158964
rect 379486 158964 379514 159004
rect 382458 158992 382464 159044
rect 382516 159032 382522 159044
rect 411346 159032 411352 159044
rect 382516 159004 411352 159032
rect 382516 158992 382522 159004
rect 411346 158992 411352 159004
rect 411404 158992 411410 159044
rect 463050 158992 463056 159044
rect 463108 159032 463114 159044
rect 469214 159032 469220 159044
rect 463108 159004 469220 159032
rect 463108 158992 463114 159004
rect 469214 158992 469220 159004
rect 469272 158992 469278 159044
rect 471422 158992 471428 159044
rect 471480 159032 471486 159044
rect 477586 159032 477592 159044
rect 471480 159004 477592 159032
rect 471480 158992 471486 159004
rect 477586 158992 477592 159004
rect 477644 158992 477650 159044
rect 397362 158964 397368 158976
rect 379486 158936 397368 158964
rect 371568 158924 371574 158936
rect 397362 158924 397368 158936
rect 397420 158924 397426 158976
rect 419350 158924 419356 158976
rect 419408 158964 419414 158976
rect 423490 158964 423496 158976
rect 419408 158936 423496 158964
rect 419408 158924 419414 158936
rect 423490 158924 423496 158936
rect 423548 158924 423554 158976
rect 465626 158924 465632 158976
rect 465684 158964 465690 158976
rect 472526 158964 472532 158976
rect 465684 158936 472532 158964
rect 465684 158924 465690 158936
rect 472526 158924 472532 158936
rect 472584 158924 472590 158976
rect 474826 158924 474832 158976
rect 474884 158964 474890 158976
rect 481634 158964 481640 158976
rect 474884 158936 481640 158964
rect 474884 158924 474890 158936
rect 481634 158924 481640 158936
rect 481692 158924 481698 158976
rect 506566 158924 506572 158976
rect 506624 158964 506630 158976
rect 508406 158964 508412 158976
rect 506624 158936 508412 158964
rect 506624 158924 506630 158936
rect 508406 158924 508412 158936
rect 508464 158924 508470 158976
rect 516686 158924 516692 158976
rect 516744 158964 516750 158976
rect 520182 158964 520188 158976
rect 516744 158936 520188 158964
rect 516744 158924 516750 158936
rect 520182 158924 520188 158936
rect 520240 158924 520246 158976
rect 363046 158896 363052 158908
rect 328696 158868 355272 158896
rect 355336 158868 363052 158896
rect 328696 158856 328702 158868
rect 355336 158828 355364 158868
rect 363046 158856 363052 158868
rect 363104 158856 363110 158908
rect 363966 158856 363972 158908
rect 364024 158896 364030 158908
rect 385862 158896 385868 158908
rect 364024 158868 385868 158896
rect 364024 158856 364030 158868
rect 385862 158856 385868 158868
rect 385920 158856 385926 158908
rect 411806 158856 411812 158908
rect 411864 158896 411870 158908
rect 413738 158896 413744 158908
rect 411864 158868 413744 158896
rect 411864 158856 411870 158868
rect 413738 158856 413744 158868
rect 413796 158856 413802 158908
rect 455506 158856 455512 158908
rect 455564 158896 455570 158908
rect 463602 158896 463608 158908
rect 455564 158868 463608 158896
rect 455564 158856 455570 158868
rect 463602 158856 463608 158868
rect 463660 158856 463666 158908
rect 464706 158856 464712 158908
rect 464764 158896 464770 158908
rect 471422 158896 471428 158908
rect 464764 158868 471428 158896
rect 464764 158856 464770 158868
rect 471422 158856 471428 158868
rect 471480 158856 471486 158908
rect 473998 158856 474004 158908
rect 474056 158896 474062 158908
rect 481358 158896 481364 158908
rect 474056 158868 481364 158896
rect 474056 158856 474062 158868
rect 481358 158856 481364 158868
rect 481416 158856 481422 158908
rect 508314 158856 508320 158908
rect 508372 158896 508378 158908
rect 509234 158896 509240 158908
rect 508372 158868 509240 158896
rect 508372 158856 508378 158868
rect 509234 158856 509240 158868
rect 509292 158856 509298 158908
rect 509326 158856 509332 158908
rect 509384 158896 509390 158908
rect 511810 158896 511816 158908
rect 509384 158868 511816 158896
rect 509384 158856 509390 158868
rect 511810 158856 511816 158868
rect 511868 158856 511874 158908
rect 515030 158856 515036 158908
rect 515088 158896 515094 158908
rect 518526 158896 518532 158908
rect 515088 158868 518532 158896
rect 515088 158856 515094 158868
rect 518526 158856 518532 158868
rect 518584 158856 518590 158908
rect 321526 158800 355364 158828
rect 268252 158732 320036 158760
rect 268252 158720 268258 158732
rect 320266 158720 320272 158772
rect 320324 158760 320330 158772
rect 321526 158760 321554 158800
rect 357250 158788 357256 158840
rect 357308 158828 357314 158840
rect 380986 158828 380992 158840
rect 357308 158800 380992 158828
rect 357308 158788 357314 158800
rect 380986 158788 380992 158800
rect 381044 158788 381050 158840
rect 398374 158788 398380 158840
rect 398432 158828 398438 158840
rect 404630 158828 404636 158840
rect 398432 158800 404636 158828
rect 398432 158788 398438 158800
rect 404630 158788 404636 158800
rect 404688 158788 404694 158840
rect 408494 158788 408500 158840
rect 408552 158828 408558 158840
rect 411254 158828 411260 158840
rect 408552 158800 411260 158828
rect 408552 158788 408558 158800
rect 411254 158788 411260 158800
rect 411312 158788 411318 158840
rect 456334 158788 456340 158840
rect 456392 158828 456398 158840
rect 463510 158828 463516 158840
rect 456392 158800 463516 158828
rect 456392 158788 456398 158800
rect 463510 158788 463516 158800
rect 463568 158788 463574 158840
rect 463878 158788 463884 158840
rect 463936 158828 463942 158840
rect 471514 158828 471520 158840
rect 463936 158800 471520 158828
rect 463936 158788 463942 158800
rect 471514 158788 471520 158800
rect 471572 158788 471578 158840
rect 507946 158788 507952 158840
rect 508004 158828 508010 158840
rect 510062 158828 510068 158840
rect 508004 158800 510068 158828
rect 508004 158788 508010 158800
rect 510062 158788 510068 158800
rect 510120 158788 510126 158840
rect 512178 158788 512184 158840
rect 512236 158828 512242 158840
rect 514294 158828 514300 158840
rect 512236 158800 514300 158828
rect 512236 158788 512242 158800
rect 514294 158788 514300 158800
rect 514352 158788 514358 158840
rect 514846 158788 514852 158840
rect 514904 158828 514910 158840
rect 517606 158828 517612 158840
rect 514904 158800 517612 158828
rect 514904 158788 514910 158800
rect 517606 158788 517612 158800
rect 517664 158788 517670 158840
rect 320324 158732 321554 158760
rect 320324 158720 320330 158732
rect 322014 158720 322020 158772
rect 322072 158760 322078 158772
rect 322072 158732 327856 158760
rect 322072 158720 322078 158732
rect 80974 158652 80980 158704
rect 81032 158692 81038 158704
rect 180794 158692 180800 158704
rect 81032 158664 180800 158692
rect 81032 158652 81038 158664
rect 180794 158652 180800 158664
rect 180852 158652 180858 158704
rect 181714 158652 181720 158704
rect 181772 158692 181778 158704
rect 256786 158692 256792 158704
rect 181772 158664 256792 158692
rect 181772 158652 181778 158664
rect 256786 158652 256792 158664
rect 256844 158652 256850 158704
rect 327828 158692 327856 158732
rect 327902 158720 327908 158772
rect 327960 158760 327966 158772
rect 327960 158732 367324 158760
rect 327960 158720 327966 158732
rect 328638 158692 328644 158704
rect 327828 158664 328644 158692
rect 328638 158652 328644 158664
rect 328696 158652 328702 158704
rect 367296 158692 367324 158732
rect 367370 158720 367376 158772
rect 367428 158760 367434 158772
rect 386046 158760 386052 158772
rect 367428 158732 386052 158760
rect 367428 158720 367434 158732
rect 386046 158720 386052 158732
rect 386104 158720 386110 158772
rect 387518 158720 387524 158772
rect 387576 158760 387582 158772
rect 390554 158760 390560 158772
rect 387576 158732 390560 158760
rect 387576 158720 387582 158732
rect 390554 158720 390560 158732
rect 390612 158720 390618 158772
rect 405090 158720 405096 158772
rect 405148 158760 405154 158772
rect 408862 158760 408868 158772
rect 405148 158732 408868 158760
rect 405148 158720 405154 158732
rect 408862 158720 408868 158732
rect 408920 158720 408926 158772
rect 412634 158720 412640 158772
rect 412692 158760 412698 158772
rect 419534 158760 419540 158772
rect 412692 158732 419540 158760
rect 412692 158720 412698 158732
rect 419534 158720 419540 158732
rect 419592 158720 419598 158772
rect 462222 158720 462228 158772
rect 462280 158760 462286 158772
rect 467926 158760 467932 158772
rect 462280 158732 467932 158760
rect 462280 158720 462286 158732
rect 467926 158720 467932 158732
rect 467984 158720 467990 158772
rect 475654 158720 475660 158772
rect 475712 158760 475718 158772
rect 482646 158760 482652 158772
rect 475712 158732 482652 158760
rect 475712 158720 475718 158732
rect 482646 158720 482652 158732
rect 482704 158720 482710 158772
rect 505278 158720 505284 158772
rect 505336 158760 505342 158772
rect 506750 158760 506756 158772
rect 505336 158732 506756 158760
rect 505336 158720 505342 158732
rect 506750 158720 506756 158732
rect 506808 158720 506814 158772
rect 509602 158720 509608 158772
rect 509660 158760 509666 158772
rect 510890 158760 510896 158772
rect 509660 158732 510896 158760
rect 509660 158720 509666 158732
rect 510890 158720 510896 158732
rect 510948 158720 510954 158772
rect 510982 158720 510988 158772
rect 511040 158760 511046 158772
rect 512638 158760 512644 158772
rect 511040 158732 512644 158760
rect 511040 158720 511046 158732
rect 512638 158720 512644 158732
rect 512696 158720 512702 158772
rect 513558 158720 513564 158772
rect 513616 158760 513622 158772
rect 515950 158760 515956 158772
rect 513616 158732 515956 158760
rect 513616 158720 513622 158732
rect 515950 158720 515956 158732
rect 516008 158720 516014 158772
rect 368474 158692 368480 158704
rect 367296 158664 368480 158692
rect 368474 158652 368480 158664
rect 368532 158652 368538 158704
rect 70854 158584 70860 158636
rect 70912 158624 70918 158636
rect 172698 158624 172704 158636
rect 70912 158596 172704 158624
rect 70912 158584 70918 158596
rect 172698 158584 172704 158596
rect 172756 158584 172762 158636
rect 174998 158584 175004 158636
rect 175056 158624 175062 158636
rect 252738 158624 252744 158636
rect 175056 158596 252744 158624
rect 175056 158584 175062 158596
rect 252738 158584 252744 158596
rect 252796 158584 252802 158636
rect 74258 158516 74264 158568
rect 74316 158556 74322 158568
rect 175366 158556 175372 158568
rect 74316 158528 175372 158556
rect 74316 158516 74322 158528
rect 175366 158516 175372 158528
rect 175424 158516 175430 158568
rect 178402 158516 178408 158568
rect 178460 158556 178466 158568
rect 255406 158556 255412 158568
rect 178460 158528 255412 158556
rect 178460 158516 178466 158528
rect 255406 158516 255412 158528
rect 255464 158516 255470 158568
rect 60826 158448 60832 158500
rect 60884 158488 60890 158500
rect 164326 158488 164332 158500
rect 60884 158460 164332 158488
rect 60884 158448 60890 158460
rect 164326 158448 164332 158460
rect 164384 158448 164390 158500
rect 164418 158448 164424 158500
rect 164476 158488 164482 158500
rect 242434 158488 242440 158500
rect 164476 158460 242440 158488
rect 164476 158448 164482 158460
rect 242434 158448 242440 158460
rect 242492 158448 242498 158500
rect 64138 158380 64144 158432
rect 64196 158420 64202 158432
rect 162118 158420 162124 158432
rect 64196 158392 162124 158420
rect 64196 158380 64202 158392
rect 162118 158380 162124 158392
rect 162176 158380 162182 158432
rect 162228 158392 167684 158420
rect 67542 158312 67548 158364
rect 67600 158352 67606 158364
rect 162228 158352 162256 158392
rect 67600 158324 162256 158352
rect 67600 158312 67606 158324
rect 162302 158312 162308 158364
rect 162360 158352 162366 158364
rect 167546 158352 167552 158364
rect 162360 158324 167552 158352
rect 162360 158312 162366 158324
rect 167546 158312 167552 158324
rect 167604 158312 167610 158364
rect 167656 158352 167684 158392
rect 168282 158380 168288 158432
rect 168340 158420 168346 158432
rect 247586 158420 247592 158432
rect 168340 158392 247592 158420
rect 168340 158380 168346 158392
rect 247586 158380 247592 158392
rect 247644 158380 247650 158432
rect 170582 158352 170588 158364
rect 167656 158324 170588 158352
rect 170582 158312 170588 158324
rect 170640 158312 170646 158364
rect 171686 158312 171692 158364
rect 171744 158352 171750 158364
rect 249886 158352 249892 158364
rect 171744 158324 249892 158352
rect 171744 158312 171750 158324
rect 249886 158312 249892 158324
rect 249944 158312 249950 158364
rect 54110 158244 54116 158296
rect 54168 158284 54174 158296
rect 153010 158284 153016 158296
rect 54168 158256 153016 158284
rect 54168 158244 54174 158256
rect 153010 158244 153016 158256
rect 153068 158244 153074 158296
rect 157426 158284 157432 158296
rect 153396 158256 157432 158284
rect 47394 158176 47400 158228
rect 47452 158216 47458 158228
rect 153102 158216 153108 158228
rect 47452 158188 153108 158216
rect 47452 158176 47458 158188
rect 153102 158176 153108 158188
rect 153160 158176 153166 158228
rect 153396 158216 153424 158256
rect 157426 158244 157432 158256
rect 157484 158244 157490 158296
rect 158254 158244 158260 158296
rect 158312 158284 158318 158296
rect 161934 158284 161940 158296
rect 158312 158256 161940 158284
rect 158312 158244 158318 158256
rect 161934 158244 161940 158256
rect 161992 158244 161998 158296
rect 162210 158244 162216 158296
rect 162268 158284 162274 158296
rect 164878 158284 164884 158296
rect 162268 158256 164884 158284
rect 162268 158244 162274 158256
rect 164878 158244 164884 158256
rect 164936 158244 164942 158296
rect 164970 158244 164976 158296
rect 165028 158284 165034 158296
rect 245010 158284 245016 158296
rect 165028 158256 245016 158284
rect 165028 158244 165034 158256
rect 245010 158244 245016 158256
rect 245068 158244 245074 158296
rect 153304 158188 153424 158216
rect 50706 158108 50712 158160
rect 50764 158148 50770 158160
rect 153304 158148 153332 158188
rect 154850 158176 154856 158228
rect 154908 158216 154914 158228
rect 164602 158216 164608 158228
rect 154908 158188 164608 158216
rect 154908 158176 154914 158188
rect 164602 158176 164608 158188
rect 164660 158176 164666 158228
rect 164786 158176 164792 158228
rect 164844 158216 164850 158228
rect 237466 158216 237472 158228
rect 164844 158188 237472 158216
rect 164844 158176 164850 158188
rect 237466 158176 237472 158188
rect 237524 158176 237530 158228
rect 249794 158176 249800 158228
rect 249852 158216 249858 158228
rect 309870 158216 309876 158228
rect 249852 158188 309876 158216
rect 249852 158176 249858 158188
rect 309870 158176 309876 158188
rect 309928 158176 309934 158228
rect 50764 158120 153332 158148
rect 50764 158108 50770 158120
rect 153470 158108 153476 158160
rect 153528 158148 153534 158160
rect 155126 158148 155132 158160
rect 153528 158120 155132 158148
rect 153528 158108 153534 158120
rect 155126 158108 155132 158120
rect 155184 158108 155190 158160
rect 155218 158108 155224 158160
rect 155276 158148 155282 158160
rect 160094 158148 160100 158160
rect 155276 158120 160100 158148
rect 155276 158108 155282 158120
rect 160094 158108 160100 158120
rect 160152 158108 160158 158160
rect 161566 158108 161572 158160
rect 161624 158148 161630 158160
rect 164418 158148 164424 158160
rect 161624 158120 164424 158148
rect 161624 158108 161630 158120
rect 164418 158108 164424 158120
rect 164476 158108 164482 158160
rect 164878 158108 164884 158160
rect 164936 158148 164942 158160
rect 238846 158148 238852 158160
rect 164936 158120 238852 158148
rect 164936 158108 164942 158120
rect 238846 158108 238852 158120
rect 238904 158108 238910 158160
rect 246390 158108 246396 158160
rect 246448 158148 246454 158160
rect 307294 158148 307300 158160
rect 246448 158120 307300 158148
rect 246448 158108 246454 158120
rect 307294 158108 307300 158120
rect 307352 158108 307358 158160
rect 37274 158040 37280 158092
rect 37332 158080 37338 158092
rect 146294 158080 146300 158092
rect 37332 158052 146300 158080
rect 37332 158040 37338 158052
rect 146294 158040 146300 158052
rect 146352 158040 146358 158092
rect 148134 158040 148140 158092
rect 148192 158080 148198 158092
rect 231946 158080 231952 158092
rect 148192 158052 231952 158080
rect 148192 158040 148198 158052
rect 231946 158040 231952 158052
rect 232004 158040 232010 158092
rect 239674 158040 239680 158092
rect 239732 158080 239738 158092
rect 302326 158080 302332 158092
rect 239732 158052 302332 158080
rect 239732 158040 239738 158052
rect 302326 158040 302332 158052
rect 302384 158040 302390 158092
rect 382 157972 388 158024
rect 440 158012 446 158024
rect 118878 158012 118884 158024
rect 440 157984 118884 158012
rect 440 157972 446 157984
rect 118878 157972 118884 157984
rect 118936 157972 118942 158024
rect 134702 157972 134708 158024
rect 134760 158012 134766 158024
rect 221918 158012 221924 158024
rect 134760 157984 221924 158012
rect 134760 157972 134766 157984
rect 221918 157972 221924 157984
rect 221976 157972 221982 158024
rect 236362 157972 236368 158024
rect 236420 158012 236426 158024
rect 299658 158012 299664 158024
rect 236420 157984 299664 158012
rect 236420 157972 236426 157984
rect 299658 157972 299664 157984
rect 299716 157972 299722 158024
rect 77570 157904 77576 157956
rect 77628 157944 77634 157956
rect 178034 157944 178040 157956
rect 77628 157916 178040 157944
rect 77628 157904 77634 157916
rect 178034 157904 178040 157916
rect 178092 157904 178098 157956
rect 185302 157944 185308 157956
rect 180996 157916 185308 157944
rect 87690 157836 87696 157888
rect 87748 157876 87754 157888
rect 180996 157876 181024 157916
rect 185302 157904 185308 157916
rect 185360 157904 185366 157956
rect 188430 157904 188436 157956
rect 188488 157944 188494 157956
rect 263042 157944 263048 157956
rect 188488 157916 263048 157944
rect 188488 157904 188494 157916
rect 263042 157904 263048 157916
rect 263100 157904 263106 157956
rect 188522 157876 188528 157888
rect 87748 157848 181024 157876
rect 181456 157848 188528 157876
rect 87748 157836 87754 157848
rect 91002 157768 91008 157820
rect 91060 157808 91066 157820
rect 181456 157808 181484 157848
rect 188522 157836 188528 157848
rect 188580 157836 188586 157888
rect 190086 157836 190092 157888
rect 190144 157876 190150 157888
rect 264330 157876 264336 157888
rect 190144 157848 264336 157876
rect 190144 157836 190150 157848
rect 264330 157836 264336 157848
rect 264388 157836 264394 157888
rect 91060 157780 181484 157808
rect 91060 157768 91066 157780
rect 181530 157768 181536 157820
rect 181588 157808 181594 157820
rect 191098 157808 191104 157820
rect 181588 157780 191104 157808
rect 181588 157768 181594 157780
rect 191098 157768 191104 157780
rect 191156 157768 191162 157820
rect 195146 157768 195152 157820
rect 195204 157808 195210 157820
rect 267734 157808 267740 157820
rect 195204 157780 267740 157808
rect 195204 157768 195210 157780
rect 267734 157768 267740 157780
rect 267792 157768 267798 157820
rect 84286 157700 84292 157752
rect 84344 157740 84350 157752
rect 182358 157740 182364 157752
rect 84344 157712 182364 157740
rect 84344 157700 84350 157712
rect 182358 157700 182364 157712
rect 182416 157700 182422 157752
rect 185118 157700 185124 157752
rect 185176 157740 185182 157752
rect 260466 157740 260472 157752
rect 185176 157712 260472 157740
rect 185176 157700 185182 157712
rect 260466 157700 260472 157712
rect 260524 157700 260530 157752
rect 94406 157632 94412 157684
rect 94464 157672 94470 157684
rect 181530 157672 181536 157684
rect 94464 157644 181536 157672
rect 94464 157632 94470 157644
rect 181530 157632 181536 157644
rect 181588 157632 181594 157684
rect 181622 157632 181628 157684
rect 181680 157672 181686 157684
rect 200298 157672 200304 157684
rect 181680 157644 200304 157672
rect 181680 157632 181686 157644
rect 200298 157632 200304 157644
rect 200356 157632 200362 157684
rect 202874 157632 202880 157684
rect 202932 157672 202938 157684
rect 255866 157672 255872 157684
rect 202932 157644 255872 157672
rect 202932 157632 202938 157644
rect 255866 157632 255872 157644
rect 255924 157632 255930 157684
rect 111150 157564 111156 157616
rect 111208 157604 111214 157616
rect 200574 157604 200580 157616
rect 111208 157576 200580 157604
rect 111208 157564 111214 157576
rect 200574 157564 200580 157576
rect 200632 157564 200638 157616
rect 200758 157564 200764 157616
rect 200816 157604 200822 157616
rect 203978 157604 203984 157616
rect 200816 157576 203984 157604
rect 200816 157564 200822 157576
rect 203978 157564 203984 157576
rect 204036 157564 204042 157616
rect 204070 157564 204076 157616
rect 204128 157604 204134 157616
rect 251450 157604 251456 157616
rect 204128 157576 251456 157604
rect 204128 157564 204134 157576
rect 251450 157564 251456 157576
rect 251508 157564 251514 157616
rect 107838 157496 107844 157548
rect 107896 157536 107902 157548
rect 200206 157536 200212 157548
rect 107896 157508 200212 157536
rect 107896 157496 107902 157508
rect 200206 157496 200212 157508
rect 200264 157496 200270 157548
rect 200298 157496 200304 157548
rect 200356 157536 200362 157548
rect 233510 157536 233516 157548
rect 200356 157508 233516 157536
rect 200356 157496 200362 157508
rect 233510 157496 233516 157508
rect 233568 157496 233574 157548
rect 117866 157428 117872 157480
rect 117924 157468 117930 157480
rect 209130 157468 209136 157480
rect 117924 157440 209136 157468
rect 117924 157428 117930 157440
rect 209130 157428 209136 157440
rect 209188 157428 209194 157480
rect 233142 157428 233148 157480
rect 233200 157468 233206 157480
rect 273806 157468 273812 157480
rect 233200 157440 273812 157468
rect 233200 157428 233206 157440
rect 273806 157428 273812 157440
rect 273864 157428 273870 157480
rect 107010 157360 107016 157412
rect 107068 157400 107074 157412
rect 107746 157400 107752 157412
rect 107068 157372 107752 157400
rect 107068 157360 107074 157372
rect 107746 157360 107752 157372
rect 107804 157360 107810 157412
rect 141418 157360 141424 157412
rect 141476 157400 141482 157412
rect 226886 157400 226892 157412
rect 141476 157372 226892 157400
rect 141476 157360 141482 157372
rect 226886 157360 226892 157372
rect 226944 157360 226950 157412
rect 45646 157292 45652 157344
rect 45704 157332 45710 157344
rect 153838 157332 153844 157344
rect 45704 157304 153844 157332
rect 45704 157292 45710 157304
rect 153838 157292 153844 157304
rect 153896 157292 153902 157344
rect 191834 157292 191840 157344
rect 191892 157332 191898 157344
rect 265158 157332 265164 157344
rect 191892 157304 265164 157332
rect 191892 157292 191898 157304
rect 265158 157292 265164 157304
rect 265216 157292 265222 157344
rect 49050 157224 49056 157276
rect 49108 157264 49114 157276
rect 156414 157264 156420 157276
rect 49108 157236 156420 157264
rect 49108 157224 49114 157236
rect 156414 157224 156420 157236
rect 156472 157224 156478 157276
rect 156598 157224 156604 157276
rect 156656 157264 156662 157276
rect 219986 157264 219992 157276
rect 156656 157236 219992 157264
rect 156656 157224 156662 157236
rect 219986 157224 219992 157236
rect 220044 157224 220050 157276
rect 283374 157224 283380 157276
rect 283432 157264 283438 157276
rect 335538 157264 335544 157276
rect 283432 157236 335544 157264
rect 283432 157224 283438 157236
rect 335538 157224 335544 157236
rect 335596 157224 335602 157276
rect 38930 157156 38936 157208
rect 38988 157196 38994 157208
rect 148778 157196 148784 157208
rect 38988 157168 148784 157196
rect 38988 157156 38994 157168
rect 148778 157156 148784 157168
rect 148836 157156 148842 157208
rect 151814 157156 151820 157208
rect 151872 157196 151878 157208
rect 152918 157196 152924 157208
rect 151872 157168 152924 157196
rect 151872 157156 151878 157168
rect 152918 157156 152924 157168
rect 152976 157156 152982 157208
rect 158714 157156 158720 157208
rect 158772 157196 158778 157208
rect 166166 157196 166172 157208
rect 158772 157168 166172 157196
rect 158772 157156 158778 157168
rect 166166 157156 166172 157168
rect 166224 157156 166230 157208
rect 166258 157156 166264 157208
rect 166316 157196 166322 157208
rect 171134 157196 171140 157208
rect 166316 157168 171140 157196
rect 166316 157156 166322 157168
rect 171134 157156 171140 157168
rect 171192 157156 171198 157208
rect 172422 157156 172428 157208
rect 172480 157196 172486 157208
rect 179690 157196 179696 157208
rect 172480 157168 179696 157196
rect 172480 157156 172486 157168
rect 179690 157156 179696 157168
rect 179748 157156 179754 157208
rect 183370 157156 183376 157208
rect 183428 157196 183434 157208
rect 258166 157196 258172 157208
rect 183428 157168 258172 157196
rect 183428 157156 183434 157168
rect 258166 157156 258172 157168
rect 258224 157156 258230 157208
rect 273254 157156 273260 157208
rect 273312 157196 273318 157208
rect 327626 157196 327632 157208
rect 273312 157168 327632 157196
rect 273312 157156 273318 157168
rect 327626 157156 327632 157168
rect 327684 157156 327690 157208
rect 31386 157088 31392 157140
rect 31444 157128 31450 157140
rect 142982 157128 142988 157140
rect 31444 157100 142988 157128
rect 31444 157088 31450 157100
rect 142982 157088 142988 157100
rect 143040 157088 143046 157140
rect 151538 157088 151544 157140
rect 151596 157128 151602 157140
rect 234798 157128 234804 157140
rect 151596 157100 234804 157128
rect 151596 157088 151602 157100
rect 234798 157088 234804 157100
rect 234856 157088 234862 157140
rect 279970 157088 279976 157140
rect 280028 157128 280034 157140
rect 333054 157128 333060 157140
rect 280028 157100 333060 157128
rect 280028 157088 280034 157100
rect 333054 157088 333060 157100
rect 333112 157088 333118 157140
rect 28074 157020 28080 157072
rect 28132 157060 28138 157072
rect 139946 157060 139952 157072
rect 28132 157032 139952 157060
rect 28132 157020 28138 157032
rect 139946 157020 139952 157032
rect 140004 157020 140010 157072
rect 142246 157020 142252 157072
rect 142304 157060 142310 157072
rect 227806 157060 227812 157072
rect 142304 157032 227812 157060
rect 142304 157020 142310 157032
rect 227806 157020 227812 157032
rect 227864 157020 227870 157072
rect 276658 157020 276664 157072
rect 276716 157060 276722 157072
rect 330478 157060 330484 157072
rect 276716 157032 330484 157060
rect 276716 157020 276722 157032
rect 330478 157020 330484 157032
rect 330536 157020 330542 157072
rect 24670 156952 24676 157004
rect 24728 156992 24734 157004
rect 137186 156992 137192 157004
rect 24728 156964 137192 156992
rect 24728 156952 24734 156964
rect 137186 156952 137192 156964
rect 137244 156952 137250 157004
rect 144822 156952 144828 157004
rect 144880 156992 144886 157004
rect 229554 156992 229560 157004
rect 144880 156964 229560 156992
rect 144880 156952 144886 156964
rect 229554 156952 229560 156964
rect 229612 156952 229618 157004
rect 232958 156952 232964 157004
rect 233016 156992 233022 157004
rect 297082 156992 297088 157004
rect 233016 156964 297088 156992
rect 233016 156952 233022 156964
rect 297082 156952 297088 156964
rect 297140 156952 297146 157004
rect 17954 156884 17960 156936
rect 18012 156924 18018 156936
rect 132678 156924 132684 156936
rect 18012 156896 132684 156924
rect 18012 156884 18018 156896
rect 132678 156884 132684 156896
rect 132736 156884 132742 156936
rect 138106 156884 138112 156936
rect 138164 156924 138170 156936
rect 224494 156924 224500 156936
rect 138164 156896 224500 156924
rect 138164 156884 138170 156896
rect 224494 156884 224500 156896
rect 224552 156884 224558 156936
rect 229646 156884 229652 156936
rect 229704 156924 229710 156936
rect 294046 156924 294052 156936
rect 229704 156896 294052 156924
rect 229704 156884 229710 156896
rect 294046 156884 294052 156896
rect 294104 156884 294110 156936
rect 296806 156884 296812 156936
rect 296864 156924 296870 156936
rect 345842 156924 345848 156936
rect 296864 156896 345848 156924
rect 296864 156884 296870 156896
rect 345842 156884 345848 156896
rect 345900 156884 345906 156936
rect 21358 156816 21364 156868
rect 21416 156856 21422 156868
rect 135254 156856 135260 156868
rect 21416 156828 135260 156856
rect 21416 156816 21422 156828
rect 135254 156816 135260 156828
rect 135312 156816 135318 156868
rect 135530 156816 135536 156868
rect 135588 156856 135594 156868
rect 222562 156856 222568 156868
rect 135588 156828 222568 156856
rect 135588 156816 135594 156828
rect 222562 156816 222568 156828
rect 222620 156816 222626 156868
rect 222838 156816 222844 156868
rect 222896 156856 222902 156868
rect 289354 156856 289360 156868
rect 222896 156828 289360 156856
rect 222896 156816 222902 156828
rect 289354 156816 289360 156828
rect 289412 156816 289418 156868
rect 300118 156816 300124 156868
rect 300176 156856 300182 156868
rect 348050 156856 348056 156868
rect 300176 156828 348056 156856
rect 300176 156816 300182 156828
rect 348050 156816 348056 156828
rect 348108 156816 348114 156868
rect 127986 156748 127992 156800
rect 128044 156788 128050 156800
rect 216858 156788 216864 156800
rect 128044 156760 216864 156788
rect 128044 156748 128050 156760
rect 216858 156748 216864 156760
rect 216916 156748 216922 156800
rect 219526 156748 219532 156800
rect 219584 156788 219590 156800
rect 286778 156788 286784 156800
rect 219584 156760 286784 156788
rect 219584 156748 219590 156760
rect 286778 156748 286784 156760
rect 286836 156748 286842 156800
rect 290090 156748 290096 156800
rect 290148 156788 290154 156800
rect 339678 156788 339684 156800
rect 290148 156760 339684 156788
rect 290148 156748 290154 156760
rect 339678 156748 339684 156760
rect 339736 156748 339742 156800
rect 14642 156680 14648 156732
rect 14700 156720 14706 156732
rect 130102 156720 130108 156732
rect 14700 156692 130108 156720
rect 14700 156680 14706 156692
rect 130102 156680 130108 156692
rect 130160 156680 130166 156732
rect 138934 156680 138940 156732
rect 138992 156720 138998 156732
rect 225138 156720 225144 156732
rect 138992 156692 225144 156720
rect 138992 156680 138998 156692
rect 225138 156680 225144 156692
rect 225196 156680 225202 156732
rect 293402 156680 293408 156732
rect 293460 156720 293466 156732
rect 343266 156720 343272 156732
rect 293460 156692 343272 156720
rect 293460 156680 293466 156692
rect 343266 156680 343272 156692
rect 343324 156680 343330 156732
rect 2038 156612 2044 156664
rect 2096 156652 2102 156664
rect 120442 156652 120448 156664
rect 2096 156624 120448 156652
rect 2096 156612 2102 156624
rect 120442 156612 120448 156624
rect 120500 156612 120506 156664
rect 121270 156612 121276 156664
rect 121328 156652 121334 156664
rect 211338 156652 211344 156664
rect 121328 156624 211344 156652
rect 121328 156612 121334 156624
rect 211338 156612 211344 156624
rect 211396 156612 211402 156664
rect 216122 156612 216128 156664
rect 216180 156652 216186 156664
rect 284202 156652 284208 156664
rect 216180 156624 284208 156652
rect 216180 156612 216186 156624
rect 284202 156612 284208 156624
rect 284260 156612 284266 156664
rect 286686 156612 286692 156664
rect 286744 156652 286750 156664
rect 338206 156652 338212 156664
rect 286744 156624 338212 156652
rect 286744 156612 286750 156624
rect 338206 156612 338212 156624
rect 338264 156612 338270 156664
rect 521838 156612 521844 156664
rect 521896 156652 521902 156664
rect 523494 156652 523500 156664
rect 521896 156624 523500 156652
rect 521896 156612 521902 156624
rect 523494 156612 523500 156624
rect 523552 156612 523558 156664
rect 69198 156544 69204 156596
rect 69256 156584 69262 156596
rect 166258 156584 166264 156596
rect 69256 156556 166264 156584
rect 69256 156544 69262 156556
rect 166258 156544 166264 156556
rect 166316 156544 166322 156596
rect 166350 156544 166356 156596
rect 166408 156584 166414 156596
rect 175918 156584 175924 156596
rect 166408 156556 175924 156584
rect 166408 156544 166414 156556
rect 175918 156544 175924 156556
rect 175976 156544 175982 156596
rect 179598 156584 179604 156596
rect 176028 156556 179604 156584
rect 79318 156476 79324 156528
rect 79376 156516 79382 156528
rect 176028 156516 176056 156556
rect 179598 156544 179604 156556
rect 179656 156544 179662 156596
rect 179690 156544 179696 156596
rect 179748 156584 179754 156596
rect 191006 156584 191012 156596
rect 179748 156556 191012 156584
rect 179748 156544 179754 156556
rect 191006 156544 191012 156556
rect 191064 156544 191070 156596
rect 191190 156544 191196 156596
rect 191248 156584 191254 156596
rect 191248 156556 195974 156584
rect 191248 156544 191254 156556
rect 79376 156488 176056 156516
rect 79376 156476 79382 156488
rect 176194 156476 176200 156528
rect 176252 156516 176258 156528
rect 176252 156488 193904 156516
rect 176252 156476 176258 156488
rect 12066 156408 12072 156460
rect 12124 156448 12130 156460
rect 109034 156448 109040 156460
rect 12124 156420 109040 156448
rect 12124 156408 12130 156420
rect 109034 156408 109040 156420
rect 109092 156408 109098 156460
rect 115382 156408 115388 156460
rect 115440 156448 115446 156460
rect 187878 156448 187884 156460
rect 115440 156420 187884 156448
rect 115440 156408 115446 156420
rect 187878 156408 187884 156420
rect 187936 156408 187942 156460
rect 89346 156340 89352 156392
rect 89404 156380 89410 156392
rect 187234 156380 187240 156392
rect 89404 156352 187240 156380
rect 89404 156340 89410 156352
rect 187234 156340 187240 156352
rect 187292 156340 187298 156392
rect 193674 156380 193680 156392
rect 190288 156352 193680 156380
rect 97718 156272 97724 156324
rect 97776 156312 97782 156324
rect 190288 156312 190316 156352
rect 193674 156340 193680 156352
rect 193732 156340 193738 156392
rect 193876 156380 193904 156488
rect 195946 156448 195974 156556
rect 200666 156544 200672 156596
rect 200724 156584 200730 156596
rect 200724 156556 201816 156584
rect 200724 156544 200730 156556
rect 198550 156476 198556 156528
rect 198608 156516 198614 156528
rect 200850 156516 200856 156528
rect 198608 156488 200856 156516
rect 198608 156476 198614 156488
rect 200850 156476 200856 156488
rect 200908 156476 200914 156528
rect 201788 156516 201816 156556
rect 201862 156544 201868 156596
rect 201920 156584 201926 156596
rect 273254 156584 273260 156596
rect 201920 156556 273260 156584
rect 201920 156544 201926 156556
rect 273254 156544 273260 156556
rect 273312 156544 273318 156596
rect 202690 156516 202696 156528
rect 201788 156488 202696 156516
rect 202690 156476 202696 156488
rect 202748 156476 202754 156528
rect 206094 156476 206100 156528
rect 206152 156516 206158 156528
rect 276014 156516 276020 156528
rect 206152 156488 276020 156516
rect 206152 156476 206158 156488
rect 276014 156476 276020 156488
rect 276072 156476 276078 156528
rect 207198 156448 207204 156460
rect 195946 156420 207204 156448
rect 207198 156408 207204 156420
rect 207256 156408 207262 156460
rect 209406 156408 209412 156460
rect 209464 156448 209470 156460
rect 279050 156448 279056 156460
rect 209464 156420 279056 156448
rect 209464 156408 209470 156420
rect 279050 156408 279056 156420
rect 279108 156408 279114 156460
rect 225782 156380 225788 156392
rect 193876 156352 225788 156380
rect 225782 156340 225788 156352
rect 225840 156340 225846 156392
rect 226242 156340 226248 156392
rect 226300 156380 226306 156392
rect 291930 156380 291936 156392
rect 226300 156352 291936 156380
rect 226300 156340 226306 156352
rect 291930 156340 291936 156352
rect 291988 156340 291994 156392
rect 97776 156284 190316 156312
rect 97776 156272 97782 156284
rect 191006 156272 191012 156324
rect 191064 156312 191070 156324
rect 238662 156312 238668 156324
rect 191064 156284 238668 156312
rect 191064 156272 191070 156284
rect 238662 156272 238668 156284
rect 238720 156272 238726 156324
rect 15470 156204 15476 156256
rect 15528 156244 15534 156256
rect 109678 156244 109684 156256
rect 15528 156216 109684 156244
rect 15528 156204 15534 156216
rect 109678 156204 109684 156216
rect 109736 156204 109742 156256
rect 114554 156204 114560 156256
rect 114612 156244 114618 156256
rect 206554 156244 206560 156256
rect 114612 156216 206560 156244
rect 114612 156204 114618 156216
rect 206554 156204 206560 156216
rect 206612 156204 206618 156256
rect 211798 156204 211804 156256
rect 211856 156244 211862 156256
rect 269482 156244 269488 156256
rect 211856 156216 269488 156244
rect 211856 156204 211862 156216
rect 269482 156204 269488 156216
rect 269540 156204 269546 156256
rect 109494 156136 109500 156188
rect 109552 156176 109558 156188
rect 200666 156176 200672 156188
rect 109552 156148 200672 156176
rect 109552 156136 109558 156148
rect 200666 156136 200672 156148
rect 200724 156136 200730 156188
rect 200758 156136 200764 156188
rect 200816 156176 200822 156188
rect 213914 156176 213920 156188
rect 200816 156148 213920 156176
rect 200816 156136 200822 156148
rect 213914 156136 213920 156148
rect 213972 156136 213978 156188
rect 260834 156176 260840 156188
rect 219406 156148 260840 156176
rect 124582 156068 124588 156120
rect 124640 156108 124646 156120
rect 214190 156108 214196 156120
rect 124640 156080 214196 156108
rect 124640 156068 124646 156080
rect 214190 156068 214196 156080
rect 214248 156068 214254 156120
rect 214558 156068 214564 156120
rect 214616 156108 214622 156120
rect 219406 156108 219434 156148
rect 260834 156136 260840 156148
rect 260892 156136 260898 156188
rect 214616 156080 219434 156108
rect 214616 156068 214622 156080
rect 223574 156068 223580 156120
rect 223632 156108 223638 156120
rect 266446 156108 266452 156120
rect 223632 156080 266452 156108
rect 223632 156068 223638 156080
rect 266446 156068 266452 156080
rect 266504 156068 266510 156120
rect 125502 156000 125508 156052
rect 125560 156040 125566 156052
rect 200758 156040 200764 156052
rect 125560 156012 200764 156040
rect 125560 156000 125566 156012
rect 200758 156000 200764 156012
rect 200816 156000 200822 156052
rect 200850 156000 200856 156052
rect 200908 156040 200914 156052
rect 270586 156040 270592 156052
rect 200908 156012 270592 156040
rect 200908 156000 200914 156012
rect 270586 156000 270592 156012
rect 270644 156000 270650 156052
rect 11238 155932 11244 155984
rect 11296 155972 11302 155984
rect 127434 155972 127440 155984
rect 11296 155944 127440 155972
rect 11296 155932 11302 155944
rect 127434 155932 127440 155944
rect 127492 155932 127498 155984
rect 131390 155932 131396 155984
rect 131448 155972 131454 155984
rect 218238 155972 218244 155984
rect 131448 155944 218244 155972
rect 131448 155932 131454 155944
rect 218238 155932 218244 155944
rect 218296 155932 218302 155984
rect 75914 155864 75920 155916
rect 75972 155904 75978 155916
rect 177022 155904 177028 155916
rect 75972 155876 177028 155904
rect 75972 155864 75978 155876
rect 177022 155864 177028 155876
rect 177080 155864 177086 155916
rect 179230 155864 179236 155916
rect 179288 155904 179294 155916
rect 255682 155904 255688 155916
rect 179288 155876 255688 155904
rect 179288 155864 179294 155876
rect 255682 155864 255688 155876
rect 255740 155864 255746 155916
rect 292574 155864 292580 155916
rect 292632 155904 292638 155916
rect 342346 155904 342352 155916
rect 292632 155876 342352 155904
rect 292632 155864 292638 155876
rect 342346 155864 342352 155876
rect 342404 155864 342410 155916
rect 75086 155796 75092 155848
rect 75144 155836 75150 155848
rect 176378 155836 176384 155848
rect 75144 155808 176384 155836
rect 75144 155796 75150 155808
rect 176378 155796 176384 155808
rect 176436 155796 176442 155848
rect 176470 155796 176476 155848
rect 176528 155836 176534 155848
rect 185670 155836 185676 155848
rect 176528 155808 185676 155836
rect 176528 155796 176534 155808
rect 185670 155796 185676 155808
rect 185728 155796 185734 155848
rect 185946 155796 185952 155848
rect 186004 155836 186010 155848
rect 261110 155836 261116 155848
rect 186004 155808 261116 155836
rect 186004 155796 186010 155808
rect 261110 155796 261116 155808
rect 261168 155796 261174 155848
rect 299290 155796 299296 155848
rect 299348 155836 299354 155848
rect 347866 155836 347872 155848
rect 299348 155808 347872 155836
rect 299348 155796 299354 155808
rect 347866 155796 347872 155808
rect 347924 155796 347930 155848
rect 43162 155728 43168 155780
rect 43220 155768 43226 155780
rect 75822 155768 75828 155780
rect 43220 155740 75828 155768
rect 43220 155728 43226 155740
rect 75822 155728 75828 155740
rect 75880 155728 75886 155780
rect 78398 155728 78404 155780
rect 78456 155768 78462 155780
rect 178954 155768 178960 155780
rect 78456 155740 178960 155768
rect 78456 155728 78462 155740
rect 178954 155728 178960 155740
rect 179012 155728 179018 155780
rect 179046 155728 179052 155780
rect 179104 155768 179110 155780
rect 185762 155768 185768 155780
rect 179104 155740 185768 155768
rect 179104 155728 179110 155740
rect 185762 155728 185768 155740
rect 185820 155728 185826 155780
rect 185854 155728 185860 155780
rect 185912 155768 185918 155780
rect 258534 155768 258540 155780
rect 185912 155740 258540 155768
rect 185912 155728 185918 155740
rect 258534 155728 258540 155740
rect 258592 155728 258598 155780
rect 295978 155728 295984 155780
rect 296036 155768 296042 155780
rect 345198 155768 345204 155780
rect 296036 155740 345204 155768
rect 296036 155728 296042 155740
rect 345198 155728 345204 155740
rect 345256 155728 345262 155780
rect 46566 155660 46572 155712
rect 46624 155700 46630 155712
rect 69658 155700 69664 155712
rect 46624 155672 69664 155700
rect 46624 155660 46630 155672
rect 69658 155660 69664 155672
rect 69716 155660 69722 155712
rect 71682 155660 71688 155712
rect 71740 155700 71746 155712
rect 173066 155700 173072 155712
rect 71740 155672 173072 155700
rect 71740 155660 71746 155672
rect 173066 155660 173072 155672
rect 173124 155660 173130 155712
rect 173158 155660 173164 155712
rect 173216 155700 173222 155712
rect 250806 155700 250812 155712
rect 173216 155672 250812 155700
rect 173216 155660 173222 155672
rect 250806 155660 250812 155672
rect 250864 155660 250870 155712
rect 289262 155660 289268 155712
rect 289320 155700 289326 155712
rect 340046 155700 340052 155712
rect 289320 155672 340052 155700
rect 289320 155660 289326 155672
rect 340046 155660 340052 155672
rect 340104 155660 340110 155712
rect 36446 155592 36452 155644
rect 36504 155632 36510 155644
rect 63494 155632 63500 155644
rect 36504 155604 63500 155632
rect 36504 155592 36510 155604
rect 63494 155592 63500 155604
rect 63552 155592 63558 155644
rect 64966 155592 64972 155644
rect 65024 155632 65030 155644
rect 168650 155632 168656 155644
rect 65024 155604 168656 155632
rect 65024 155592 65030 155604
rect 168650 155592 168656 155604
rect 168708 155592 168714 155644
rect 169110 155592 169116 155644
rect 169168 155632 169174 155644
rect 247126 155632 247132 155644
rect 169168 155604 247132 155632
rect 169168 155592 169174 155604
rect 247126 155592 247132 155604
rect 247184 155592 247190 155644
rect 269942 155592 269948 155644
rect 270000 155632 270006 155644
rect 325326 155632 325332 155644
rect 270000 155604 325332 155632
rect 270000 155592 270006 155604
rect 325326 155592 325332 155604
rect 325384 155592 325390 155644
rect 51534 155524 51540 155576
rect 51592 155564 51598 155576
rect 158346 155564 158352 155576
rect 51592 155536 158352 155564
rect 51592 155524 51598 155536
rect 158346 155524 158352 155536
rect 158404 155524 158410 155576
rect 159082 155524 159088 155576
rect 159140 155564 159146 155576
rect 240594 155564 240600 155576
rect 159140 155536 240600 155564
rect 159140 155524 159146 155536
rect 240594 155524 240600 155536
rect 240652 155524 240658 155576
rect 266538 155524 266544 155576
rect 266596 155564 266602 155576
rect 321830 155564 321836 155576
rect 266596 155536 321836 155564
rect 266596 155524 266602 155536
rect 321830 155524 321836 155536
rect 321888 155524 321894 155576
rect 340414 155524 340420 155576
rect 340472 155564 340478 155576
rect 379238 155564 379244 155576
rect 340472 155536 379244 155564
rect 340472 155524 340478 155536
rect 379238 155524 379244 155536
rect 379296 155524 379302 155576
rect 54938 155456 54944 155508
rect 54996 155496 55002 155508
rect 160922 155496 160928 155508
rect 54996 155468 160928 155496
rect 54996 155456 55002 155468
rect 160922 155456 160928 155468
rect 160980 155456 160986 155508
rect 162394 155456 162400 155508
rect 162452 155496 162458 155508
rect 243078 155496 243084 155508
rect 162452 155468 243084 155496
rect 162452 155456 162458 155468
rect 243078 155456 243084 155468
rect 243136 155456 243142 155508
rect 263226 155456 263232 155508
rect 263284 155496 263290 155508
rect 320174 155496 320180 155508
rect 263284 155468 320180 155496
rect 263284 155456 263290 155468
rect 320174 155456 320180 155468
rect 320232 155456 320238 155508
rect 337102 155456 337108 155508
rect 337160 155496 337166 155508
rect 376662 155496 376668 155508
rect 337160 155468 376668 155496
rect 337160 155456 337166 155468
rect 376662 155456 376668 155468
rect 376720 155456 376726 155508
rect 48222 155388 48228 155440
rect 48280 155428 48286 155440
rect 151722 155428 151728 155440
rect 48280 155400 151728 155428
rect 48280 155388 48286 155400
rect 151722 155388 151728 155400
rect 151780 155388 151786 155440
rect 152734 155388 152740 155440
rect 152792 155428 152798 155440
rect 155586 155428 155592 155440
rect 152792 155400 155592 155428
rect 152792 155388 152798 155400
rect 155586 155388 155592 155400
rect 155644 155388 155650 155440
rect 155678 155388 155684 155440
rect 155736 155428 155742 155440
rect 237558 155428 237564 155440
rect 155736 155400 237564 155428
rect 155736 155388 155742 155400
rect 237558 155388 237564 155400
rect 237616 155388 237622 155440
rect 259822 155388 259828 155440
rect 259880 155428 259886 155440
rect 317598 155428 317604 155440
rect 259880 155400 317604 155428
rect 259880 155388 259886 155400
rect 317598 155388 317604 155400
rect 317656 155388 317662 155440
rect 332870 155388 332876 155440
rect 332928 155428 332934 155440
rect 373442 155428 373448 155440
rect 332928 155400 373448 155428
rect 332928 155388 332934 155400
rect 373442 155388 373448 155400
rect 373500 155388 373506 155440
rect 4522 155320 4528 155372
rect 4580 155360 4586 155372
rect 122006 155360 122012 155372
rect 4580 155332 122012 155360
rect 4580 155320 4586 155332
rect 122006 155320 122012 155332
rect 122064 155320 122070 155372
rect 123754 155320 123760 155372
rect 123812 155360 123818 155372
rect 128446 155360 128452 155372
rect 123812 155332 128452 155360
rect 123812 155320 123818 155332
rect 128446 155320 128452 155332
rect 128504 155320 128510 155372
rect 148962 155320 148968 155372
rect 149020 155360 149026 155372
rect 232866 155360 232872 155372
rect 149020 155332 232872 155360
rect 149020 155320 149026 155332
rect 232866 155320 232872 155332
rect 232924 155320 232930 155372
rect 256510 155320 256516 155372
rect 256568 155360 256574 155372
rect 315022 155360 315028 155372
rect 256568 155332 315028 155360
rect 256568 155320 256574 155332
rect 315022 155320 315028 155332
rect 315080 155320 315086 155372
rect 329558 155320 329564 155372
rect 329616 155360 329622 155372
rect 370866 155360 370872 155372
rect 329616 155332 370872 155360
rect 329616 155320 329622 155332
rect 370866 155320 370872 155332
rect 370924 155320 370930 155372
rect 376570 155320 376576 155372
rect 376628 155360 376634 155372
rect 406838 155360 406844 155372
rect 376628 155332 406844 155360
rect 376628 155320 376634 155332
rect 406838 155320 406844 155332
rect 406896 155320 406902 155372
rect 8754 155252 8760 155304
rect 8812 155292 8818 155304
rect 125594 155292 125600 155304
rect 8812 155264 125600 155292
rect 8812 155252 8818 155264
rect 125594 155252 125600 155264
rect 125652 155252 125658 155304
rect 132218 155252 132224 155304
rect 132276 155292 132282 155304
rect 219526 155292 219532 155304
rect 132276 155264 219532 155292
rect 132276 155252 132282 155264
rect 219526 155252 219532 155264
rect 219584 155252 219590 155304
rect 243170 155252 243176 155304
rect 243228 155292 243234 155304
rect 243228 155264 248414 155292
rect 243228 155252 243234 155264
rect 5350 155184 5356 155236
rect 5408 155224 5414 155236
rect 123018 155224 123024 155236
rect 5408 155196 123024 155224
rect 5408 155184 5414 155196
rect 123018 155184 123024 155196
rect 123076 155184 123082 155236
rect 128814 155184 128820 155236
rect 128872 155224 128878 155236
rect 217410 155224 217416 155236
rect 128872 155196 217416 155224
rect 128872 155184 128878 155196
rect 217410 155184 217416 155196
rect 217468 155184 217474 155236
rect 233878 155184 233884 155236
rect 233936 155224 233942 155236
rect 243538 155224 243544 155236
rect 233936 155196 243544 155224
rect 233936 155184 233942 155196
rect 243538 155184 243544 155196
rect 243596 155184 243602 155236
rect 248386 155224 248414 155264
rect 253106 155252 253112 155304
rect 253164 155292 253170 155304
rect 312446 155292 312452 155304
rect 253164 155264 312452 155292
rect 253164 155252 253170 155264
rect 312446 155252 312452 155264
rect 312504 155252 312510 155304
rect 373166 155252 373172 155304
rect 373224 155292 373230 155304
rect 403158 155292 403164 155304
rect 373224 155264 403164 155292
rect 373224 155252 373230 155264
rect 403158 155252 403164 155264
rect 403216 155252 403222 155304
rect 304718 155224 304724 155236
rect 248386 155196 304724 155224
rect 304718 155184 304724 155196
rect 304776 155184 304782 155236
rect 306006 155184 306012 155236
rect 306064 155224 306070 155236
rect 352926 155224 352932 155236
rect 306064 155196 352932 155224
rect 306064 155184 306070 155196
rect 352926 155184 352932 155196
rect 352984 155184 352990 155236
rect 369854 155184 369860 155236
rect 369912 155224 369918 155236
rect 401686 155224 401692 155236
rect 369912 155196 401692 155224
rect 369912 155184 369918 155196
rect 401686 155184 401692 155196
rect 401744 155184 401750 155236
rect 56594 155116 56600 155168
rect 56652 155156 56658 155168
rect 76466 155156 76472 155168
rect 56652 155128 76472 155156
rect 56652 155116 56658 155128
rect 76466 155116 76472 155128
rect 76524 155116 76530 155168
rect 81802 155116 81808 155168
rect 81860 155156 81866 155168
rect 181346 155156 181352 155168
rect 81860 155128 181352 155156
rect 81860 155116 81866 155128
rect 181346 155116 181352 155128
rect 181404 155116 181410 155168
rect 182542 155116 182548 155168
rect 182600 155156 182606 155168
rect 185394 155156 185400 155168
rect 182600 155128 185400 155156
rect 182600 155116 182606 155128
rect 185394 155116 185400 155128
rect 185452 155116 185458 155168
rect 185486 155116 185492 155168
rect 185544 155156 185550 155168
rect 185544 155128 189212 155156
rect 185544 155116 185550 155128
rect 73430 155048 73436 155100
rect 73488 155088 73494 155100
rect 81434 155088 81440 155100
rect 73488 155060 81440 155088
rect 73488 155048 73494 155060
rect 81434 155048 81440 155060
rect 81492 155048 81498 155100
rect 88518 155048 88524 155100
rect 88576 155088 88582 155100
rect 186590 155088 186596 155100
rect 88576 155060 186596 155088
rect 88576 155048 88582 155060
rect 186590 155048 186596 155060
rect 186648 155048 186654 155100
rect 189184 155088 189212 155128
rect 189258 155116 189264 155168
rect 189316 155156 189322 155168
rect 263778 155156 263784 155168
rect 189316 155128 263784 155156
rect 189316 155116 189322 155128
rect 263778 155116 263784 155128
rect 263836 155116 263842 155168
rect 302694 155116 302700 155168
rect 302752 155156 302758 155168
rect 349338 155156 349344 155168
rect 302752 155128 349344 155156
rect 302752 155116 302758 155128
rect 349338 155116 349344 155128
rect 349396 155116 349402 155168
rect 192386 155088 192392 155100
rect 189184 155060 192392 155088
rect 192386 155048 192392 155060
rect 192444 155048 192450 155100
rect 192662 155048 192668 155100
rect 192720 155088 192726 155100
rect 266262 155088 266268 155100
rect 192720 155060 266268 155088
rect 192720 155048 192726 155060
rect 266262 155048 266268 155060
rect 266320 155048 266326 155100
rect 312722 155048 312728 155100
rect 312780 155088 312786 155100
rect 357894 155088 357900 155100
rect 312780 155060 357900 155088
rect 312780 155048 312786 155060
rect 357894 155048 357900 155060
rect 357952 155048 357958 155100
rect 91830 154980 91836 155032
rect 91888 155020 91894 155032
rect 189166 155020 189172 155032
rect 91888 154992 189172 155020
rect 91888 154980 91894 154992
rect 189166 154980 189172 154992
rect 189224 154980 189230 155032
rect 195974 154980 195980 155032
rect 196032 155020 196038 155032
rect 268838 155020 268844 155032
rect 196032 154992 268844 155020
rect 196032 154980 196038 154992
rect 268838 154980 268844 154992
rect 268896 154980 268902 155032
rect 86034 154912 86040 154964
rect 86092 154952 86098 154964
rect 183554 154952 183560 154964
rect 86092 154924 183560 154952
rect 86092 154912 86098 154924
rect 183554 154912 183560 154924
rect 183612 154912 183618 154964
rect 185578 154912 185584 154964
rect 185636 154952 185642 154964
rect 191742 154952 191748 154964
rect 185636 154924 191748 154952
rect 185636 154912 185642 154924
rect 191742 154912 191748 154924
rect 191800 154912 191806 154964
rect 199378 154912 199384 154964
rect 199436 154952 199442 154964
rect 271414 154952 271420 154964
rect 199436 154924 271420 154952
rect 199436 154912 199442 154924
rect 271414 154912 271420 154924
rect 271472 154912 271478 154964
rect 96062 154844 96068 154896
rect 96120 154884 96126 154896
rect 185486 154884 185492 154896
rect 96120 154856 185492 154884
rect 96120 154844 96126 154856
rect 185486 154844 185492 154856
rect 185544 154844 185550 154896
rect 185670 154844 185676 154896
rect 185728 154884 185734 154896
rect 185728 154856 195974 154884
rect 185728 154844 185734 154856
rect 98638 154776 98644 154828
rect 98696 154816 98702 154828
rect 194318 154816 194324 154828
rect 98696 154788 194324 154816
rect 98696 154776 98702 154788
rect 194318 154776 194324 154788
rect 194376 154776 194382 154828
rect 195946 154816 195974 154856
rect 202782 154844 202788 154896
rect 202840 154884 202846 154896
rect 273438 154884 273444 154896
rect 202840 154856 273444 154884
rect 202840 154844 202846 154856
rect 273438 154844 273444 154856
rect 273496 154844 273502 154896
rect 228358 154816 228364 154828
rect 195946 154788 228364 154816
rect 228358 154776 228364 154788
rect 228416 154776 228422 154828
rect 281626 154816 281632 154828
rect 229756 154788 281632 154816
rect 95234 154708 95240 154760
rect 95292 154748 95298 154760
rect 185578 154748 185584 154760
rect 95292 154720 185584 154748
rect 95292 154708 95298 154720
rect 185578 154708 185584 154720
rect 185636 154708 185642 154760
rect 185762 154708 185768 154760
rect 185820 154748 185826 154760
rect 229646 154748 229652 154760
rect 185820 154720 229652 154748
rect 185820 154708 185826 154720
rect 229646 154708 229652 154720
rect 229704 154708 229710 154760
rect 118786 154640 118792 154692
rect 118844 154680 118850 154692
rect 209774 154680 209780 154692
rect 118844 154652 209780 154680
rect 118844 154640 118850 154652
rect 209774 154640 209780 154652
rect 209832 154640 209838 154692
rect 212810 154640 212816 154692
rect 212868 154680 212874 154692
rect 229756 154680 229784 154788
rect 281626 154776 281632 154788
rect 281684 154776 281690 154828
rect 229830 154708 229836 154760
rect 229888 154748 229894 154760
rect 242894 154748 242900 154760
rect 229888 154720 242900 154748
rect 229888 154708 229894 154720
rect 242894 154708 242900 154720
rect 242952 154708 242958 154760
rect 243538 154708 243544 154760
rect 243596 154748 243602 154760
rect 276474 154748 276480 154760
rect 243596 154720 276480 154748
rect 243596 154708 243602 154720
rect 276474 154708 276480 154720
rect 276532 154708 276538 154760
rect 212868 154652 229784 154680
rect 212868 154640 212874 154652
rect 241422 154640 241428 154692
rect 241480 154680 241486 154692
rect 292574 154680 292580 154692
rect 241480 154652 292580 154680
rect 241480 154640 241486 154652
rect 292574 154640 292580 154652
rect 292632 154640 292638 154692
rect 122098 154572 122104 154624
rect 122156 154612 122162 154624
rect 212258 154612 212264 154624
rect 122156 154584 212264 154612
rect 122156 154572 122162 154584
rect 212258 154572 212264 154584
rect 212316 154572 212322 154624
rect 227714 154572 227720 154624
rect 227772 154612 227778 154624
rect 272058 154612 272064 154624
rect 227772 154584 272064 154612
rect 227772 154572 227778 154584
rect 272058 154572 272064 154584
rect 272116 154572 272122 154624
rect 58342 154504 58348 154556
rect 58400 154544 58406 154556
rect 58400 154516 152504 154544
rect 58400 154504 58406 154516
rect 44174 154436 44180 154488
rect 44232 154476 44238 154488
rect 146754 154476 146760 154488
rect 44232 154448 146760 154476
rect 44232 154436 44238 154448
rect 146754 154436 146760 154448
rect 146812 154436 146818 154488
rect 147030 154436 147036 154488
rect 147088 154476 147094 154488
rect 148318 154476 148324 154488
rect 147088 154448 148324 154476
rect 147088 154436 147094 154448
rect 148318 154436 148324 154448
rect 148376 154436 148382 154488
rect 41506 154368 41512 154420
rect 41564 154408 41570 154420
rect 146570 154408 146576 154420
rect 41564 154380 146576 154408
rect 41564 154368 41570 154380
rect 146570 154368 146576 154380
rect 146628 154368 146634 154420
rect 146938 154368 146944 154420
rect 146996 154408 147002 154420
rect 152366 154408 152372 154420
rect 146996 154380 152372 154408
rect 146996 154368 147002 154380
rect 152366 154368 152372 154380
rect 152424 154368 152430 154420
rect 152476 154408 152504 154516
rect 152734 154504 152740 154556
rect 152792 154544 152798 154556
rect 210510 154544 210516 154556
rect 152792 154516 210516 154544
rect 152792 154504 152798 154516
rect 210510 154504 210516 154516
rect 210568 154504 210574 154556
rect 215294 154504 215300 154556
rect 215352 154544 215358 154556
rect 283190 154544 283196 154556
rect 215352 154516 283196 154544
rect 215352 154504 215358 154516
rect 283190 154504 283196 154516
rect 283248 154504 283254 154556
rect 285858 154504 285864 154556
rect 285916 154544 285922 154556
rect 337470 154544 337476 154556
rect 285916 154516 337476 154544
rect 285916 154504 285922 154516
rect 337470 154504 337476 154516
rect 337528 154504 337534 154556
rect 352282 154504 352288 154556
rect 352340 154544 352346 154556
rect 388898 154544 388904 154556
rect 352340 154516 388904 154544
rect 352340 154504 352346 154516
rect 388898 154504 388904 154516
rect 388956 154504 388962 154556
rect 153010 154436 153016 154488
rect 153068 154476 153074 154488
rect 207842 154476 207848 154488
rect 153068 154448 207848 154476
rect 153068 154436 153074 154448
rect 207842 154436 207848 154448
rect 207900 154436 207906 154488
rect 211246 154436 211252 154488
rect 211304 154476 211310 154488
rect 280982 154476 280988 154488
rect 211304 154448 280988 154476
rect 211304 154436 211310 154448
rect 280982 154436 280988 154448
rect 281040 154436 281046 154488
rect 281718 154436 281724 154488
rect 281776 154476 281782 154488
rect 334894 154476 334900 154488
rect 281776 154448 334900 154476
rect 281776 154436 281782 154448
rect 334894 154436 334900 154448
rect 334952 154436 334958 154488
rect 349246 154436 349252 154488
rect 349304 154476 349310 154488
rect 386322 154476 386328 154488
rect 349304 154448 386328 154476
rect 349304 154436 349310 154448
rect 386322 154436 386328 154448
rect 386380 154436 386386 154488
rect 163314 154408 163320 154420
rect 152476 154380 163320 154408
rect 163314 154368 163320 154380
rect 163372 154368 163378 154420
rect 164142 154368 164148 154420
rect 164200 154408 164206 154420
rect 165706 154408 165712 154420
rect 164200 154380 165712 154408
rect 164200 154368 164206 154380
rect 165706 154368 165712 154380
rect 165764 154368 165770 154420
rect 165798 154368 165804 154420
rect 165856 154408 165862 154420
rect 175918 154408 175924 154420
rect 165856 154380 175924 154408
rect 165856 154368 165862 154380
rect 175918 154368 175924 154380
rect 175976 154368 175982 154420
rect 176010 154368 176016 154420
rect 176068 154408 176074 154420
rect 181254 154408 181260 154420
rect 176068 154380 181260 154408
rect 176068 154368 176074 154380
rect 181254 154368 181260 154380
rect 181312 154368 181318 154420
rect 181990 154368 181996 154420
rect 182048 154408 182054 154420
rect 254026 154408 254032 154420
rect 182048 154380 254032 154408
rect 182048 154368 182054 154380
rect 254026 154368 254032 154380
rect 254084 154368 254090 154420
rect 258258 154368 258264 154420
rect 258316 154408 258322 154420
rect 316954 154408 316960 154420
rect 258316 154380 316960 154408
rect 258316 154368 258322 154380
rect 316954 154368 316960 154380
rect 317012 154368 317018 154420
rect 345566 154368 345572 154420
rect 345624 154408 345630 154420
rect 383838 154408 383844 154420
rect 345624 154380 383844 154408
rect 345624 154368 345630 154380
rect 383838 154368 383844 154380
rect 383896 154368 383902 154420
rect 116026 154300 116032 154352
rect 116084 154340 116090 154352
rect 121914 154340 121920 154352
rect 116084 154312 121920 154340
rect 116084 154300 116090 154312
rect 121914 154300 121920 154312
rect 121972 154300 121978 154352
rect 123938 154300 123944 154352
rect 123996 154340 124002 154352
rect 127342 154340 127348 154352
rect 123996 154312 127348 154340
rect 123996 154300 124002 154312
rect 127342 154300 127348 154312
rect 127400 154300 127406 154352
rect 127526 154300 127532 154352
rect 127584 154340 127590 154352
rect 189810 154340 189816 154352
rect 127584 154312 189816 154340
rect 127584 154300 127590 154312
rect 189810 154300 189816 154312
rect 189868 154300 189874 154352
rect 191190 154300 191196 154352
rect 191248 154340 191254 154352
rect 202046 154340 202052 154352
rect 191248 154312 202052 154340
rect 191248 154300 191254 154312
rect 202046 154300 202052 154312
rect 202104 154300 202110 154352
rect 208578 154300 208584 154352
rect 208636 154340 208642 154352
rect 278406 154340 278412 154352
rect 208636 154312 278412 154340
rect 208636 154300 208642 154312
rect 278406 154300 278412 154312
rect 278464 154300 278470 154352
rect 278774 154300 278780 154352
rect 278832 154340 278838 154352
rect 332410 154340 332416 154352
rect 278832 154312 332416 154340
rect 278832 154300 278838 154312
rect 332410 154300 332416 154312
rect 332468 154300 332474 154352
rect 342254 154300 342260 154352
rect 342312 154340 342318 154352
rect 381170 154340 381176 154352
rect 342312 154312 381176 154340
rect 342312 154300 342318 154312
rect 381170 154300 381176 154312
rect 381228 154300 381234 154352
rect 400306 154300 400312 154352
rect 400364 154340 400370 154352
rect 425514 154340 425520 154352
rect 400364 154312 425520 154340
rect 400364 154300 400370 154312
rect 425514 154300 425520 154312
rect 425572 154300 425578 154352
rect 30558 154232 30564 154284
rect 30616 154272 30622 154284
rect 137278 154272 137284 154284
rect 30616 154244 137284 154272
rect 30616 154232 30622 154244
rect 137278 154232 137284 154244
rect 137336 154232 137342 154284
rect 189534 154272 189540 154284
rect 137388 154244 189540 154272
rect 26878 154164 26884 154216
rect 26936 154204 26942 154216
rect 136082 154204 136088 154216
rect 26936 154176 136088 154204
rect 26936 154164 26942 154176
rect 136082 154164 136088 154176
rect 136140 154164 136146 154216
rect 137388 154204 137416 154244
rect 189534 154232 189540 154244
rect 189592 154232 189598 154284
rect 191006 154232 191012 154284
rect 191064 154272 191070 154284
rect 199470 154272 199476 154284
rect 191064 154244 199476 154272
rect 191064 154232 191070 154244
rect 199470 154232 199476 154244
rect 199528 154232 199534 154284
rect 204530 154232 204536 154284
rect 204588 154272 204594 154284
rect 274634 154272 274640 154284
rect 204588 154244 274640 154272
rect 204588 154232 204594 154244
rect 274634 154232 274640 154244
rect 274692 154232 274698 154284
rect 275094 154232 275100 154284
rect 275152 154272 275158 154284
rect 329926 154272 329932 154284
rect 275152 154244 329932 154272
rect 275152 154232 275158 154244
rect 329926 154232 329932 154244
rect 329984 154232 329990 154284
rect 339586 154232 339592 154284
rect 339644 154272 339650 154284
rect 378594 154272 378600 154284
rect 339644 154244 378600 154272
rect 339644 154232 339650 154244
rect 378594 154232 378600 154244
rect 378652 154232 378658 154284
rect 393406 154232 393412 154284
rect 393464 154272 393470 154284
rect 419718 154272 419724 154284
rect 393464 154244 419724 154272
rect 393464 154232 393470 154244
rect 419718 154232 419724 154244
rect 419776 154232 419782 154284
rect 137204 154176 137416 154204
rect 23474 154096 23480 154148
rect 23532 154136 23538 154148
rect 137094 154136 137100 154148
rect 23532 154108 137100 154136
rect 23532 154096 23538 154108
rect 137094 154096 137100 154108
rect 137152 154096 137158 154148
rect 13814 154028 13820 154080
rect 13872 154068 13878 154080
rect 129458 154068 129464 154080
rect 13872 154040 129464 154068
rect 13872 154028 13878 154040
rect 129458 154028 129464 154040
rect 129516 154028 129522 154080
rect 129550 154028 129556 154080
rect 129608 154068 129614 154080
rect 137204 154068 137232 154176
rect 139486 154164 139492 154216
rect 139544 154204 139550 154216
rect 146938 154204 146944 154216
rect 139544 154176 146944 154204
rect 139544 154164 139550 154176
rect 146938 154164 146944 154176
rect 146996 154164 147002 154216
rect 147122 154164 147128 154216
rect 147180 154204 147186 154216
rect 147180 154176 148088 154204
rect 147180 154164 147186 154176
rect 137554 154096 137560 154148
rect 137612 154136 137618 154148
rect 146846 154136 146852 154148
rect 137612 154108 146852 154136
rect 137612 154096 137618 154108
rect 146846 154096 146852 154108
rect 146904 154096 146910 154148
rect 148060 154136 148088 154176
rect 148226 154164 148232 154216
rect 148284 154204 148290 154216
rect 153194 154204 153200 154216
rect 148284 154176 153200 154204
rect 148284 154164 148290 154176
rect 153194 154164 153200 154176
rect 153252 154164 153258 154216
rect 154482 154164 154488 154216
rect 154540 154204 154546 154216
rect 175826 154204 175832 154216
rect 154540 154176 175832 154204
rect 154540 154164 154546 154176
rect 175826 154164 175832 154176
rect 175884 154164 175890 154216
rect 176102 154164 176108 154216
rect 176160 154204 176166 154216
rect 253382 154204 253388 154216
rect 176160 154176 253388 154204
rect 176160 154164 176166 154176
rect 253382 154164 253388 154176
rect 253440 154164 253446 154216
rect 255314 154164 255320 154216
rect 255372 154204 255378 154216
rect 314378 154204 314384 154216
rect 255372 154176 314384 154204
rect 255372 154164 255378 154176
rect 314378 154164 314384 154176
rect 314436 154164 314442 154216
rect 335630 154164 335636 154216
rect 335688 154204 335694 154216
rect 376018 154204 376024 154216
rect 335688 154176 376024 154204
rect 335688 154164 335694 154176
rect 376018 154164 376024 154176
rect 376076 154164 376082 154216
rect 386598 154164 386604 154216
rect 386656 154204 386662 154216
rect 414566 154204 414572 154216
rect 386656 154176 414572 154204
rect 386656 154164 386662 154176
rect 414566 154164 414572 154176
rect 414624 154164 414630 154216
rect 166258 154136 166264 154148
rect 148060 154108 166264 154136
rect 166258 154096 166264 154108
rect 166316 154096 166322 154148
rect 166350 154096 166356 154148
rect 166408 154136 166414 154148
rect 175734 154136 175740 154148
rect 166408 154108 175740 154136
rect 166408 154096 166414 154108
rect 175734 154096 175740 154108
rect 175792 154096 175798 154148
rect 175918 154096 175924 154148
rect 175976 154136 175982 154148
rect 245654 154136 245660 154148
rect 175976 154108 245660 154136
rect 175976 154096 175982 154108
rect 245654 154096 245660 154108
rect 245712 154096 245718 154148
rect 248414 154096 248420 154148
rect 248472 154136 248478 154148
rect 309226 154136 309232 154148
rect 248472 154108 309232 154136
rect 248472 154096 248478 154108
rect 309226 154096 309232 154108
rect 309284 154096 309290 154148
rect 325694 154096 325700 154148
rect 325752 154136 325758 154148
rect 368290 154136 368296 154148
rect 325752 154108 368296 154136
rect 325752 154096 325758 154108
rect 368290 154096 368296 154108
rect 368348 154096 368354 154148
rect 389726 154096 389732 154148
rect 389784 154136 389790 154148
rect 417142 154136 417148 154148
rect 389784 154108 417148 154136
rect 389784 154096 389790 154108
rect 417142 154096 417148 154108
rect 417200 154096 417206 154148
rect 129608 154040 137232 154068
rect 129608 154028 129614 154040
rect 137278 154028 137284 154080
rect 137336 154068 137342 154080
rect 142338 154068 142344 154080
rect 137336 154040 142344 154068
rect 137336 154028 137342 154040
rect 142338 154028 142344 154040
rect 142396 154028 142402 154080
rect 144914 154028 144920 154080
rect 144972 154068 144978 154080
rect 144972 154040 147996 154068
rect 144972 154028 144978 154040
rect 16574 153960 16580 154012
rect 16632 154000 16638 154012
rect 132034 154000 132040 154012
rect 16632 153972 132040 154000
rect 16632 153960 16638 153972
rect 132034 153960 132040 153972
rect 132092 153960 132098 154012
rect 136082 153960 136088 154012
rect 136140 154000 136146 154012
rect 139762 154000 139768 154012
rect 136140 153972 139768 154000
rect 136140 153960 136146 153972
rect 139762 153960 139768 153972
rect 139820 153960 139826 154012
rect 474 153892 480 153944
rect 532 153932 538 153944
rect 119798 153932 119804 153944
rect 532 153904 119804 153932
rect 532 153892 538 153904
rect 119798 153892 119804 153904
rect 119856 153892 119862 153944
rect 120074 153892 120080 153944
rect 120132 153932 120138 153944
rect 120132 153904 121868 153932
rect 120132 153892 120138 153904
rect 2958 153824 2964 153876
rect 3016 153864 3022 153876
rect 121730 153864 121736 153876
rect 3016 153836 121736 153864
rect 3016 153824 3022 153836
rect 121730 153824 121736 153836
rect 121788 153824 121794 153876
rect 121840 153864 121868 153904
rect 121914 153892 121920 153944
rect 121972 153932 121978 153944
rect 127526 153932 127532 153944
rect 121972 153904 127532 153932
rect 121972 153892 121978 153904
rect 127526 153892 127532 153904
rect 127584 153892 127590 153944
rect 146662 153932 146668 153944
rect 127636 153904 146668 153932
rect 127636 153864 127664 153904
rect 146662 153892 146668 153904
rect 146720 153892 146726 153944
rect 146754 153892 146760 153944
rect 146812 153932 146818 153944
rect 147766 153932 147772 153944
rect 146812 153904 147772 153932
rect 146812 153892 146818 153904
rect 147766 153892 147772 153904
rect 147824 153892 147830 153944
rect 147968 153932 147996 154040
rect 152918 154028 152924 154080
rect 152976 154068 152982 154080
rect 235442 154068 235448 154080
rect 152976 154040 235448 154068
rect 152976 154028 152982 154040
rect 235442 154028 235448 154040
rect 235500 154028 235506 154080
rect 245562 154028 245568 154080
rect 245620 154068 245626 154080
rect 306650 154068 306656 154080
rect 245620 154040 306656 154068
rect 245620 154028 245626 154040
rect 306650 154028 306656 154040
rect 306708 154028 306714 154080
rect 316126 154028 316132 154080
rect 316184 154068 316190 154080
rect 360654 154068 360660 154080
rect 316184 154040 360660 154068
rect 316184 154028 316190 154040
rect 360654 154028 360660 154040
rect 360712 154028 360718 154080
rect 363138 154028 363144 154080
rect 363196 154068 363202 154080
rect 396534 154068 396540 154080
rect 363196 154040 396540 154068
rect 363196 154028 363202 154040
rect 396534 154028 396540 154040
rect 396592 154028 396598 154080
rect 400122 154028 400128 154080
rect 400180 154068 400186 154080
rect 424870 154068 424876 154080
rect 400180 154040 424876 154068
rect 400180 154028 400186 154040
rect 424870 154028 424876 154040
rect 424928 154028 424934 154080
rect 148318 153960 148324 154012
rect 148376 154000 148382 154012
rect 230934 154000 230940 154012
rect 148376 153972 230940 154000
rect 148376 153960 148382 153972
rect 230934 153960 230940 153972
rect 230992 153960 230998 154012
rect 231854 153960 231860 154012
rect 231912 154000 231918 154012
rect 296438 154000 296444 154012
rect 231912 153972 296444 154000
rect 231912 153960 231918 153972
rect 296438 153960 296444 153972
rect 296496 153960 296502 154012
rect 322842 153960 322848 154012
rect 322900 154000 322906 154012
rect 365806 154000 365812 154012
rect 322900 153972 365812 154000
rect 322900 153960 322906 153972
rect 365806 153960 365812 153972
rect 365864 153960 365870 154012
rect 379606 153960 379612 154012
rect 379664 154000 379670 154012
rect 409414 154000 409420 154012
rect 379664 153972 409420 154000
rect 379664 153960 379670 153972
rect 409414 153960 409420 153972
rect 409472 153960 409478 154012
rect 230290 153932 230296 153944
rect 147968 153904 230296 153932
rect 230290 153892 230296 153904
rect 230348 153892 230354 153944
rect 234706 153892 234712 153944
rect 234764 153932 234770 153944
rect 299014 153932 299020 153944
rect 234764 153904 299020 153932
rect 234764 153892 234770 153904
rect 299014 153892 299020 153904
rect 299072 153892 299078 153944
rect 318794 153892 318800 153944
rect 318852 153932 318858 153944
rect 363138 153932 363144 153944
rect 318852 153904 363144 153932
rect 318852 153892 318858 153904
rect 363138 153892 363144 153904
rect 363196 153892 363202 153944
rect 383286 153892 383292 153944
rect 383344 153932 383350 153944
rect 411990 153932 411996 153944
rect 383344 153904 411996 153932
rect 383344 153892 383350 153904
rect 411990 153892 411996 153904
rect 412048 153892 412054 153944
rect 421098 153892 421104 153944
rect 421156 153932 421162 153944
rect 440878 153932 440884 153944
rect 421156 153904 440884 153932
rect 421156 153892 421162 153904
rect 440878 153892 440884 153904
rect 440936 153892 440942 153944
rect 121840 153836 127664 153864
rect 128354 153824 128360 153876
rect 128412 153864 128418 153876
rect 215478 153864 215484 153876
rect 128412 153836 215484 153864
rect 128412 153824 128418 153836
rect 215478 153824 215484 153836
rect 215536 153824 215542 153876
rect 218054 153824 218060 153876
rect 218112 153864 218118 153876
rect 286134 153864 286140 153876
rect 218112 153836 286140 153864
rect 218112 153824 218118 153836
rect 286134 153824 286140 153836
rect 286192 153824 286198 153876
rect 309134 153824 309140 153876
rect 309192 153864 309198 153876
rect 355502 153864 355508 153876
rect 309192 153836 355508 153864
rect 309192 153824 309198 153836
rect 355502 153824 355508 153836
rect 355560 153824 355566 153876
rect 356054 153824 356060 153876
rect 356112 153864 356118 153876
rect 391474 153864 391480 153876
rect 356112 153836 391480 153864
rect 356112 153824 356118 153836
rect 391474 153824 391480 153836
rect 391532 153824 391538 153876
rect 396074 153824 396080 153876
rect 396132 153864 396138 153876
rect 422294 153864 422300 153876
rect 396132 153836 422300 153864
rect 396132 153824 396138 153836
rect 422294 153824 422300 153836
rect 422352 153824 422358 153876
rect 62114 153756 62120 153808
rect 62172 153796 62178 153808
rect 166166 153796 166172 153808
rect 62172 153768 166172 153796
rect 62172 153756 62178 153768
rect 166166 153756 166172 153768
rect 166224 153756 166230 153808
rect 166258 153756 166264 153808
rect 166316 153796 166322 153808
rect 212902 153796 212908 153808
rect 166316 153768 212908 153796
rect 166316 153756 166322 153768
rect 212902 153756 212908 153768
rect 212960 153756 212966 153808
rect 224954 153756 224960 153808
rect 225012 153796 225018 153808
rect 291286 153796 291292 153808
rect 225012 153768 291292 153796
rect 225012 153756 225018 153768
rect 291286 153756 291292 153768
rect 291344 153756 291350 153808
rect 358998 153756 359004 153808
rect 359056 153796 359062 153808
rect 394050 153796 394056 153808
rect 359056 153768 394056 153796
rect 359056 153756 359062 153768
rect 394050 153756 394056 153768
rect 394108 153756 394114 153808
rect 425238 153756 425244 153808
rect 425296 153796 425302 153808
rect 432690 153796 432696 153808
rect 425296 153768 432696 153796
rect 425296 153756 425302 153768
rect 432690 153756 432696 153768
rect 432748 153756 432754 153808
rect 71774 153688 71780 153740
rect 71832 153728 71838 153740
rect 173894 153728 173900 153740
rect 71832 153700 173900 153728
rect 71832 153688 71838 153700
rect 173894 153688 173900 153700
rect 173952 153688 173958 153740
rect 175826 153688 175832 153740
rect 175884 153728 175890 153740
rect 218054 153728 218060 153740
rect 175884 153700 218060 153728
rect 175884 153688 175890 153700
rect 218054 153688 218060 153700
rect 218112 153688 218118 153740
rect 227990 153688 227996 153740
rect 228048 153728 228054 153740
rect 293862 153728 293868 153740
rect 228048 153700 293868 153728
rect 228048 153688 228054 153700
rect 293862 153688 293868 153700
rect 293920 153688 293926 153740
rect 365714 153688 365720 153740
rect 365772 153728 365778 153740
rect 399110 153728 399116 153740
rect 365772 153700 399116 153728
rect 365772 153688 365778 153700
rect 399110 153688 399116 153700
rect 399168 153688 399174 153740
rect 81894 153620 81900 153672
rect 81952 153660 81958 153672
rect 175642 153660 175648 153672
rect 81952 153632 175648 153660
rect 81952 153620 81958 153632
rect 175642 153620 175648 153632
rect 175700 153620 175706 153672
rect 175734 153620 175740 153672
rect 175792 153660 175798 153672
rect 223206 153660 223212 153672
rect 175792 153632 223212 153660
rect 175792 153620 175798 153632
rect 223206 153620 223212 153632
rect 223264 153620 223270 153672
rect 241514 153620 241520 153672
rect 241572 153660 241578 153672
rect 304074 153660 304080 153672
rect 241572 153632 304080 153660
rect 241572 153620 241578 153632
rect 304074 153620 304080 153632
rect 304132 153620 304138 153672
rect 101306 153552 101312 153604
rect 101364 153592 101370 153604
rect 101364 153564 191144 153592
rect 101364 153552 101370 153564
rect 104894 153484 104900 153536
rect 104952 153524 104958 153536
rect 191006 153524 191012 153536
rect 104952 153496 191012 153524
rect 104952 153484 104958 153496
rect 191006 153484 191012 153496
rect 191064 153484 191070 153536
rect 191116 153524 191144 153564
rect 191282 153552 191288 153604
rect 191340 153592 191346 153604
rect 236086 153592 236092 153604
rect 191340 153564 236092 153592
rect 191340 153552 191346 153564
rect 236086 153552 236092 153564
rect 236144 153552 236150 153604
rect 238938 153552 238944 153604
rect 238996 153592 239002 153604
rect 301590 153592 301596 153604
rect 238996 153564 301596 153592
rect 238996 153552 239002 153564
rect 301590 153552 301596 153564
rect 301648 153552 301654 153604
rect 196894 153524 196900 153536
rect 191116 153496 196900 153524
rect 196894 153484 196900 153496
rect 196952 153484 196958 153536
rect 198734 153484 198740 153536
rect 198792 153524 198798 153536
rect 248874 153524 248880 153536
rect 198792 153496 248880 153524
rect 198792 153484 198798 153496
rect 248874 153484 248880 153496
rect 248932 153484 248938 153536
rect 251542 153484 251548 153536
rect 251600 153524 251606 153536
rect 311802 153524 311808 153536
rect 251600 153496 311808 153524
rect 251600 153484 251606 153496
rect 311802 153484 311808 153496
rect 311860 153484 311866 153536
rect 107930 153416 107936 153468
rect 107988 153456 107994 153468
rect 191190 153456 191196 153468
rect 107988 153428 191196 153456
rect 107988 153416 107994 153428
rect 191190 153416 191196 153428
rect 191248 153416 191254 153468
rect 191282 153416 191288 153468
rect 191340 153456 191346 153468
rect 194962 153456 194968 153468
rect 191340 153428 194968 153456
rect 191340 153416 191346 153428
rect 194962 153416 194968 153428
rect 195020 153416 195026 153468
rect 196158 153416 196164 153468
rect 196216 153456 196222 153468
rect 241238 153456 241244 153468
rect 196216 153428 241244 153456
rect 196216 153416 196222 153428
rect 241238 153416 241244 153428
rect 241296 153416 241302 153468
rect 264974 153416 264980 153468
rect 265032 153456 265038 153468
rect 321738 153456 321744 153468
rect 265032 153428 321744 153456
rect 265032 153416 265038 153428
rect 321738 153416 321744 153428
rect 321796 153416 321802 153468
rect 426158 153416 426164 153468
rect 426216 153456 426222 153468
rect 429470 153456 429476 153468
rect 426216 153428 429476 153456
rect 426216 153416 426222 153428
rect 429470 153416 429476 153428
rect 429528 153416 429534 153468
rect 111794 153348 111800 153400
rect 111852 153388 111858 153400
rect 204622 153388 204628 153400
rect 111852 153360 204628 153388
rect 111852 153348 111858 153360
rect 204622 153348 204628 153360
rect 204680 153348 204686 153400
rect 262398 153348 262404 153400
rect 262456 153388 262462 153400
rect 319530 153388 319536 153400
rect 262456 153360 319536 153388
rect 262456 153348 262462 153360
rect 319530 153348 319536 153360
rect 319588 153348 319594 153400
rect 112254 153280 112260 153332
rect 112312 153320 112318 153332
rect 205266 153320 205272 153332
rect 112312 153292 205272 153320
rect 112312 153280 112318 153292
rect 205266 153280 205272 153292
rect 205324 153280 205330 153332
rect 269114 153280 269120 153332
rect 269172 153320 269178 153332
rect 274542 153320 274548 153332
rect 269172 153292 274548 153320
rect 269172 153280 269178 153292
rect 274542 153280 274548 153292
rect 274600 153280 274606 153332
rect 274634 153280 274640 153332
rect 274692 153320 274698 153332
rect 275830 153320 275836 153332
rect 274692 153292 275836 153320
rect 274692 153280 274698 153292
rect 275830 153280 275836 153292
rect 275888 153280 275894 153332
rect 275922 153280 275928 153332
rect 275980 153320 275986 153332
rect 324682 153320 324688 153332
rect 275980 153292 324688 153320
rect 275980 153280 275986 153292
rect 324682 153280 324688 153292
rect 324740 153280 324746 153332
rect 34514 153212 34520 153264
rect 34572 153252 34578 153264
rect 145558 153252 145564 153264
rect 34572 153224 145564 153252
rect 34572 153212 34578 153224
rect 145558 153212 145564 153224
rect 145616 153212 145622 153264
rect 146662 153212 146668 153264
rect 146720 153252 146726 153264
rect 189442 153252 189448 153264
rect 146720 153224 189448 153252
rect 146720 153212 146726 153224
rect 189442 153212 189448 153224
rect 189500 153212 189506 153264
rect 189534 153212 189540 153264
rect 189592 153252 189598 153264
rect 197538 153252 197544 153264
rect 189592 153224 197544 153252
rect 189592 153212 189598 153224
rect 197538 153212 197544 153224
rect 197596 153212 197602 153264
rect 197630 153212 197636 153264
rect 197688 153252 197694 153264
rect 246298 153252 246304 153264
rect 197688 153224 246304 153252
rect 197688 153212 197694 153224
rect 246298 153212 246304 153224
rect 246356 153212 246362 153264
rect 271966 153212 271972 153264
rect 272024 153252 272030 153264
rect 327258 153252 327264 153264
rect 272024 153224 327264 153252
rect 272024 153212 272030 153224
rect 327258 153212 327264 153224
rect 327316 153212 327322 153264
rect 360838 153212 360844 153264
rect 360896 153252 360902 153264
rect 360896 153224 365116 153252
rect 360896 153212 360902 153224
rect 107746 153144 107752 153196
rect 107804 153184 107810 153196
rect 200758 153184 200764 153196
rect 107804 153156 200764 153184
rect 107804 153144 107810 153156
rect 200758 153144 200764 153156
rect 200816 153144 200822 153196
rect 218146 153144 218152 153196
rect 218204 153184 218210 153196
rect 226242 153184 226248 153196
rect 218204 153156 226248 153184
rect 218204 153144 218210 153156
rect 226242 153144 226248 153156
rect 226300 153144 226306 153196
rect 226334 153144 226340 153196
rect 226392 153184 226398 153196
rect 231578 153184 231584 153196
rect 226392 153156 231584 153184
rect 226392 153144 226398 153156
rect 231578 153144 231584 153156
rect 231636 153144 231642 153196
rect 237190 153144 237196 153196
rect 237248 153184 237254 153196
rect 300302 153184 300308 153196
rect 237248 153156 300308 153184
rect 237248 153144 237254 153156
rect 300302 153144 300308 153156
rect 300360 153144 300366 153196
rect 300854 153144 300860 153196
rect 300912 153184 300918 153196
rect 302878 153184 302884 153196
rect 300912 153156 302884 153184
rect 300912 153144 300918 153156
rect 302878 153144 302884 153156
rect 302936 153144 302942 153196
rect 303614 153144 303620 153196
rect 303672 153184 303678 153196
rect 351638 153184 351644 153196
rect 303672 153156 351644 153184
rect 303672 153144 303678 153156
rect 351638 153144 351644 153156
rect 351696 153144 351702 153196
rect 354766 153144 354772 153196
rect 354824 153184 354830 153196
rect 364978 153184 364984 153196
rect 354824 153156 364984 153184
rect 354824 153144 354830 153156
rect 364978 153144 364984 153156
rect 365036 153144 365042 153196
rect 365088 153184 365116 153224
rect 395154 153184 395160 153196
rect 365088 153156 395160 153184
rect 395154 153144 395160 153156
rect 395212 153144 395218 153196
rect 395522 153144 395528 153196
rect 395580 153184 395586 153196
rect 397822 153184 397828 153196
rect 395580 153156 397828 153184
rect 395580 153144 395586 153156
rect 397822 153144 397828 153156
rect 397880 153144 397886 153196
rect 401594 153144 401600 153196
rect 401652 153184 401658 153196
rect 415854 153184 415860 153196
rect 401652 153156 415860 153184
rect 401652 153144 401658 153156
rect 415854 153144 415860 153156
rect 415912 153144 415918 153196
rect 416958 153144 416964 153196
rect 417016 153184 417022 153196
rect 438302 153184 438308 153196
rect 417016 153156 438308 153184
rect 417016 153144 417022 153156
rect 438302 153144 438308 153156
rect 438360 153144 438366 153196
rect 438854 153144 438860 153196
rect 438912 153184 438918 153196
rect 442442 153184 442448 153196
rect 438912 153156 442448 153184
rect 438912 153144 438918 153156
rect 442442 153144 442448 153156
rect 442500 153144 442506 153196
rect 442902 153144 442908 153196
rect 442960 153184 442966 153196
rect 457622 153184 457628 153196
rect 442960 153156 457628 153184
rect 442960 153144 442966 153156
rect 457622 153144 457628 153156
rect 457680 153144 457686 153196
rect 458174 153144 458180 153196
rect 458232 153184 458238 153196
rect 460750 153184 460756 153196
rect 458232 153156 460756 153184
rect 458232 153144 458238 153156
rect 460750 153144 460756 153156
rect 460808 153144 460814 153196
rect 463602 153144 463608 153196
rect 463660 153184 463666 153196
rect 467190 153184 467196 153196
rect 463660 153156 467196 153184
rect 463660 153144 463666 153156
rect 467190 153144 467196 153156
rect 467248 153144 467254 153196
rect 471514 153144 471520 153196
rect 471572 153184 471578 153196
rect 473630 153184 473636 153196
rect 471572 153156 473636 153184
rect 471572 153144 471578 153156
rect 473630 153144 473636 153156
rect 473688 153144 473694 153196
rect 474734 153144 474740 153196
rect 474792 153184 474798 153196
rect 476850 153184 476856 153196
rect 474792 153156 476856 153184
rect 474792 153144 474798 153156
rect 476850 153144 476856 153156
rect 476908 153144 476914 153196
rect 477586 153144 477592 153196
rect 477644 153184 477650 153196
rect 479334 153184 479340 153196
rect 477644 153156 479340 153184
rect 477644 153144 477650 153156
rect 479334 153144 479340 153156
rect 479392 153144 479398 153196
rect 483198 153144 483204 153196
rect 483256 153184 483262 153196
rect 488442 153184 488448 153196
rect 483256 153156 488448 153184
rect 483256 153144 483262 153156
rect 488442 153144 488448 153156
rect 488500 153144 488506 153196
rect 489914 153144 489920 153196
rect 489972 153184 489978 153196
rect 493502 153184 493508 153196
rect 489972 153156 493508 153184
rect 489972 153144 489978 153156
rect 493502 153144 493508 153156
rect 493560 153144 493566 153196
rect 494146 153144 494152 153196
rect 494204 153184 494210 153196
rect 496722 153184 496728 153196
rect 494204 153156 496728 153184
rect 494204 153144 494210 153156
rect 496722 153144 496728 153156
rect 496780 153144 496786 153196
rect 496814 153144 496820 153196
rect 496872 153184 496878 153196
rect 499298 153184 499304 153196
rect 496872 153156 499304 153184
rect 496872 153144 496878 153156
rect 499298 153144 499304 153156
rect 499356 153144 499362 153196
rect 500862 153144 500868 153196
rect 500920 153184 500926 153196
rect 501874 153184 501880 153196
rect 500920 153156 501880 153184
rect 500920 153144 500926 153156
rect 501874 153144 501880 153156
rect 501932 153144 501938 153196
rect 503346 153144 503352 153196
rect 503404 153184 503410 153196
rect 503806 153184 503812 153196
rect 503404 153156 503812 153184
rect 503404 153144 503410 153156
rect 503806 153144 503812 153156
rect 503864 153144 503870 153196
rect 511626 153144 511632 153196
rect 511684 153184 511690 153196
rect 513466 153184 513472 153196
rect 511684 153156 513472 153184
rect 511684 153144 511690 153156
rect 513466 153144 513472 153156
rect 513524 153144 513530 153196
rect 514202 153144 514208 153196
rect 514260 153184 514266 153196
rect 516134 153184 516140 153196
rect 514260 153156 516140 153184
rect 514260 153144 514266 153156
rect 516134 153144 516140 153156
rect 516192 153144 516198 153196
rect 30190 153076 30196 153128
rect 30248 153116 30254 153128
rect 110966 153116 110972 153128
rect 30248 153088 110972 153116
rect 30248 153076 30254 153088
rect 110966 153076 110972 153088
rect 111024 153076 111030 153128
rect 116394 153076 116400 153128
rect 116452 153116 116458 153128
rect 208486 153116 208492 153128
rect 116452 153088 208492 153116
rect 116452 153076 116458 153088
rect 208486 153076 208492 153088
rect 208544 153076 208550 153128
rect 214006 153076 214012 153128
rect 214064 153116 214070 153128
rect 279326 153116 279332 153128
rect 214064 153088 279332 153116
rect 214064 153076 214070 153088
rect 279326 153076 279332 153088
rect 279384 153076 279390 153128
rect 279786 153076 279792 153128
rect 279844 153116 279850 153128
rect 282270 153116 282276 153128
rect 279844 153088 282276 153116
rect 279844 153076 279850 153088
rect 282270 153076 282276 153088
rect 282328 153076 282334 153128
rect 284294 153076 284300 153128
rect 284352 153116 284358 153128
rect 336826 153116 336832 153128
rect 284352 153088 336832 153116
rect 284352 153076 284358 153088
rect 336826 153076 336832 153088
rect 336884 153076 336890 153128
rect 337010 153076 337016 153128
rect 337068 153116 337074 153128
rect 338758 153116 338764 153128
rect 337068 153088 338764 153116
rect 337068 153076 337074 153088
rect 338758 153076 338764 153088
rect 338816 153076 338822 153128
rect 340874 153076 340880 153128
rect 340932 153116 340938 153128
rect 379882 153116 379888 153128
rect 340932 153088 379888 153116
rect 340932 153076 340938 153088
rect 379882 153076 379888 153088
rect 379940 153076 379946 153128
rect 384942 153076 384948 153128
rect 385000 153116 385006 153128
rect 413094 153116 413100 153128
rect 385000 153088 413100 153116
rect 385000 153076 385006 153088
rect 413094 153076 413100 153088
rect 413152 153076 413158 153128
rect 414106 153076 414112 153128
rect 414164 153116 414170 153128
rect 431862 153116 431868 153128
rect 414164 153088 431868 153116
rect 414164 153076 414170 153088
rect 431862 153076 431868 153088
rect 431920 153076 431926 153128
rect 431954 153076 431960 153128
rect 432012 153116 432018 153128
rect 432782 153116 432788 153128
rect 432012 153088 432788 153116
rect 432012 153076 432018 153088
rect 432782 153076 432788 153088
rect 432840 153076 432846 153128
rect 437934 153076 437940 153128
rect 437992 153116 437998 153128
rect 454402 153116 454408 153128
rect 437992 153088 454408 153116
rect 437992 153076 437998 153088
rect 454402 153076 454408 153088
rect 454460 153076 454466 153128
rect 463510 153076 463516 153128
rect 463568 153116 463574 153128
rect 467834 153116 467840 153128
rect 463568 153088 467840 153116
rect 463568 153076 463574 153088
rect 467834 153076 467840 153088
rect 467892 153076 467898 153128
rect 471422 153076 471428 153128
rect 471480 153116 471486 153128
rect 474274 153116 474280 153128
rect 471480 153088 474280 153116
rect 471480 153076 471486 153088
rect 474274 153076 474280 153088
rect 474332 153076 474338 153128
rect 475010 153076 475016 153128
rect 475068 153116 475074 153128
rect 477494 153116 477500 153128
rect 475068 153088 477500 153116
rect 475068 153076 475074 153088
rect 477494 153076 477500 153088
rect 477552 153076 477558 153128
rect 484394 153076 484400 153128
rect 484452 153116 484458 153128
rect 489638 153116 489644 153128
rect 484452 153088 489644 153116
rect 484452 153076 484458 153088
rect 489638 153076 489644 153088
rect 489696 153076 489702 153128
rect 491294 153076 491300 153128
rect 491352 153116 491358 153128
rect 494790 153116 494796 153128
rect 491352 153088 494796 153116
rect 491352 153076 491358 153088
rect 494790 153076 494796 153088
rect 494848 153076 494854 153128
rect 495434 153076 495440 153128
rect 495492 153116 495498 153128
rect 498010 153116 498016 153128
rect 495492 153088 498016 153116
rect 495492 153076 495498 153088
rect 498010 153076 498016 153088
rect 498068 153076 498074 153128
rect 500954 153076 500960 153128
rect 501012 153116 501018 153128
rect 502518 153116 502524 153128
rect 501012 153088 502524 153116
rect 501012 153076 501018 153088
rect 502518 153076 502524 153088
rect 502576 153076 502582 153128
rect 512914 153076 512920 153128
rect 512972 153116 512978 153128
rect 515122 153116 515128 153128
rect 512972 153088 515128 153116
rect 512972 153076 512978 153088
rect 515122 153076 515128 153088
rect 515180 153076 515186 153128
rect 23290 153008 23296 153060
rect 23348 153048 23354 153060
rect 108022 153048 108028 153060
rect 23348 153020 108028 153048
rect 23348 153008 23354 153020
rect 108022 153008 108028 153020
rect 108080 153008 108086 153060
rect 110322 153008 110328 153060
rect 110380 153048 110386 153060
rect 203334 153048 203340 153060
rect 110380 153020 203340 153048
rect 110380 153008 110386 153020
rect 203334 153008 203340 153020
rect 203392 153008 203398 153060
rect 210234 153008 210240 153060
rect 210292 153048 210298 153060
rect 221274 153048 221280 153060
rect 210292 153020 221280 153048
rect 210292 153008 210298 153020
rect 221274 153008 221280 153020
rect 221332 153008 221338 153060
rect 230566 153008 230572 153060
rect 230624 153048 230630 153060
rect 295794 153048 295800 153060
rect 230624 153020 295800 153048
rect 230624 153008 230630 153020
rect 295794 153008 295800 153020
rect 295852 153008 295858 153060
rect 305178 153008 305184 153060
rect 305236 153048 305242 153060
rect 352282 153048 352288 153060
rect 305236 153020 352288 153048
rect 305236 153008 305242 153020
rect 352282 153008 352288 153020
rect 352340 153008 352346 153060
rect 358906 153008 358912 153060
rect 358964 153048 358970 153060
rect 364886 153048 364892 153060
rect 358964 153020 364892 153048
rect 358964 153008 358970 153020
rect 364886 153008 364892 153020
rect 364944 153008 364950 153060
rect 364978 153008 364984 153060
rect 365036 153048 365042 153060
rect 390186 153048 390192 153060
rect 365036 153020 390192 153048
rect 365036 153008 365042 153020
rect 390186 153008 390192 153020
rect 390244 153008 390250 153060
rect 391934 153008 391940 153060
rect 391992 153048 391998 153060
rect 417786 153048 417792 153060
rect 391992 153020 417792 153048
rect 391992 153008 391998 153020
rect 417786 153008 417792 153020
rect 417844 153008 417850 153060
rect 418154 153008 418160 153060
rect 418212 153048 418218 153060
rect 438946 153048 438952 153060
rect 418212 153020 438952 153048
rect 418212 153008 418218 153020
rect 438946 153008 438952 153020
rect 439004 153008 439010 153060
rect 440418 153008 440424 153060
rect 440476 153048 440482 153060
rect 455690 153048 455696 153060
rect 440476 153020 455696 153048
rect 440476 153008 440482 153020
rect 455690 153008 455696 153020
rect 455748 153008 455754 153060
rect 464614 153008 464620 153060
rect 464672 153048 464678 153060
rect 468386 153048 468392 153060
rect 464672 153020 468392 153048
rect 464672 153008 464678 153020
rect 468386 153008 468392 153020
rect 468444 153008 468450 153060
rect 472526 153008 472532 153060
rect 472584 153048 472590 153060
rect 474918 153048 474924 153060
rect 472584 153020 474924 153048
rect 472584 153008 472590 153020
rect 474918 153008 474924 153020
rect 474976 153008 474982 153060
rect 476114 153008 476120 153060
rect 476172 153048 476178 153060
rect 478230 153048 478236 153060
rect 476172 153020 478236 153048
rect 476172 153008 476178 153020
rect 478230 153008 478236 153020
rect 478288 153008 478294 153060
rect 490006 153008 490012 153060
rect 490064 153048 490070 153060
rect 494146 153048 494152 153060
rect 490064 153020 494152 153048
rect 490064 153008 490070 153020
rect 494146 153008 494152 153020
rect 494204 153008 494210 153060
rect 495986 153008 495992 153060
rect 496044 153048 496050 153060
rect 498654 153048 498660 153060
rect 496044 153020 498660 153048
rect 496044 153008 496050 153020
rect 498654 153008 498660 153020
rect 498712 153008 498718 153060
rect 499666 153008 499672 153060
rect 499724 153048 499730 153060
rect 501230 153048 501236 153060
rect 499724 153020 501236 153048
rect 499724 153008 499730 153020
rect 501230 153008 501236 153020
rect 501288 153008 501294 153060
rect 9490 152940 9496 152992
rect 9548 152980 9554 152992
rect 92566 152980 92572 152992
rect 9548 152952 92572 152980
rect 9548 152940 9554 152952
rect 92566 152940 92572 152952
rect 92624 152940 92630 152992
rect 99558 152940 99564 152992
rect 99616 152980 99622 152992
rect 195606 152980 195612 152992
rect 99616 152952 195612 152980
rect 99616 152940 99622 152952
rect 195606 152940 195612 152952
rect 195664 152940 195670 152992
rect 196066 152940 196072 152992
rect 196124 152980 196130 152992
rect 216122 152980 216128 152992
rect 196124 152952 216128 152980
rect 196124 152940 196130 152952
rect 216122 152940 216128 152952
rect 216180 152940 216186 152992
rect 216674 152940 216680 152992
rect 216732 152980 216738 152992
rect 284846 152980 284852 152992
rect 216732 152952 284852 152980
rect 216732 152940 216738 152952
rect 284846 152940 284852 152952
rect 284904 152940 284910 152992
rect 290182 152940 290188 152992
rect 290240 152980 290246 152992
rect 341334 152980 341340 152992
rect 290240 152952 341340 152980
rect 290240 152940 290246 152952
rect 341334 152940 341340 152952
rect 341392 152940 341398 152992
rect 346394 152940 346400 152992
rect 346452 152980 346458 152992
rect 346452 152952 383654 152980
rect 346452 152940 346458 152952
rect 93302 152872 93308 152924
rect 93360 152912 93366 152924
rect 190454 152912 190460 152924
rect 93360 152884 190460 152912
rect 93360 152872 93366 152884
rect 190454 152872 190460 152884
rect 190512 152872 190518 152924
rect 194502 152872 194508 152924
rect 194560 152912 194566 152924
rect 211062 152912 211068 152924
rect 194560 152884 211068 152912
rect 194560 152872 194566 152884
rect 211062 152872 211068 152884
rect 211120 152872 211126 152924
rect 211154 152872 211160 152924
rect 211212 152912 211218 152924
rect 280338 152912 280344 152924
rect 211212 152884 280344 152912
rect 211212 152872 211218 152884
rect 280338 152872 280344 152884
rect 280396 152872 280402 152924
rect 284110 152872 284116 152924
rect 284168 152912 284174 152924
rect 336182 152912 336188 152924
rect 284168 152884 336188 152912
rect 284168 152872 284174 152884
rect 336182 152872 336188 152884
rect 336240 152872 336246 152924
rect 338114 152872 338120 152924
rect 338172 152912 338178 152924
rect 377950 152912 377956 152924
rect 338172 152884 377956 152912
rect 338172 152872 338178 152884
rect 377950 152872 377956 152884
rect 378008 152872 378014 152924
rect 380894 152872 380900 152924
rect 380952 152912 380958 152924
rect 383194 152912 383200 152924
rect 380952 152884 383200 152912
rect 380952 152872 380958 152884
rect 383194 152872 383200 152884
rect 383252 152872 383258 152924
rect 383626 152912 383654 152952
rect 383746 152940 383752 152992
rect 383804 152980 383810 152992
rect 412634 152980 412640 152992
rect 383804 152952 412640 152980
rect 383804 152940 383810 152952
rect 412634 152940 412640 152952
rect 412692 152940 412698 152992
rect 415210 152940 415216 152992
rect 415268 152980 415274 152992
rect 436370 152980 436376 152992
rect 415268 152952 436376 152980
rect 415268 152940 415274 152952
rect 436370 152940 436376 152952
rect 436428 152940 436434 152992
rect 436462 152940 436468 152992
rect 436520 152980 436526 152992
rect 442350 152980 442356 152992
rect 436520 152952 442356 152980
rect 436520 152940 436526 152952
rect 442350 152940 442356 152952
rect 442408 152940 442414 152992
rect 442442 152940 442448 152992
rect 442500 152980 442506 152992
rect 446766 152980 446772 152992
rect 442500 152952 446772 152980
rect 442500 152940 442506 152952
rect 446766 152940 446772 152952
rect 446824 152940 446830 152992
rect 464890 152940 464896 152992
rect 464948 152980 464954 152992
rect 469122 152980 469128 152992
rect 464948 152952 469128 152980
rect 464948 152940 464954 152952
rect 469122 152940 469128 152952
rect 469180 152940 469186 152992
rect 473354 152940 473360 152992
rect 473412 152980 473418 152992
rect 475562 152980 475568 152992
rect 473412 152952 475568 152980
rect 473412 152940 473418 152952
rect 475562 152940 475568 152952
rect 475620 152940 475626 152992
rect 494238 152940 494244 152992
rect 494296 152980 494302 152992
rect 497366 152980 497372 152992
rect 494296 152952 497372 152980
rect 494296 152940 494302 152952
rect 497366 152940 497372 152952
rect 497424 152940 497430 152992
rect 384390 152912 384396 152924
rect 383626 152884 384396 152912
rect 384390 152872 384396 152884
rect 384448 152872 384454 152924
rect 388438 152872 388444 152924
rect 388496 152912 388502 152924
rect 408770 152912 408776 152924
rect 388496 152884 408776 152912
rect 388496 152872 388502 152884
rect 408770 152872 408776 152884
rect 408828 152872 408834 152924
rect 410702 152872 410708 152924
rect 410760 152912 410766 152924
rect 433150 152912 433156 152924
rect 410760 152884 433156 152912
rect 410760 152872 410766 152884
rect 433150 152872 433156 152884
rect 433208 152872 433214 152924
rect 434714 152872 434720 152924
rect 434772 152912 434778 152924
rect 451826 152912 451832 152924
rect 434772 152884 451832 152912
rect 434772 152872 434778 152884
rect 451826 152872 451832 152884
rect 451884 152872 451890 152924
rect 465350 152872 465356 152924
rect 465408 152912 465414 152924
rect 469766 152912 469772 152924
rect 465408 152884 469772 152912
rect 465408 152872 465414 152884
rect 469766 152872 469772 152884
rect 469824 152872 469830 152924
rect 473446 152872 473452 152924
rect 473504 152912 473510 152924
rect 476206 152912 476212 152924
rect 473504 152884 476212 152912
rect 473504 152872 473510 152884
rect 476206 152872 476212 152884
rect 476264 152872 476270 152924
rect 492674 152872 492680 152924
rect 492732 152912 492738 152924
rect 496078 152912 496084 152924
rect 492732 152884 496084 152912
rect 492732 152872 492738 152884
rect 496078 152872 496084 152884
rect 496136 152872 496142 152924
rect 33134 152804 33140 152856
rect 33192 152844 33198 152856
rect 137278 152844 137284 152856
rect 33192 152816 137284 152844
rect 33192 152804 33198 152816
rect 137278 152804 137284 152816
rect 137336 152804 137342 152856
rect 139394 152804 139400 152856
rect 139452 152844 139458 152856
rect 141694 152844 141700 152856
rect 139452 152816 141700 152844
rect 139452 152804 139458 152816
rect 141694 152804 141700 152816
rect 141752 152804 141758 152856
rect 141786 152804 141792 152856
rect 141844 152844 141850 152856
rect 146938 152844 146944 152856
rect 141844 152816 146944 152844
rect 141844 152804 141850 152816
rect 146938 152804 146944 152816
rect 146996 152804 147002 152856
rect 149054 152804 149060 152856
rect 149112 152844 149118 152856
rect 164878 152844 164884 152856
rect 149112 152816 164884 152844
rect 149112 152804 149118 152816
rect 164878 152804 164884 152816
rect 164936 152804 164942 152856
rect 170030 152804 170036 152856
rect 170088 152844 170094 152856
rect 249518 152844 249524 152856
rect 170088 152816 249524 152844
rect 170088 152804 170094 152816
rect 249518 152804 249524 152816
rect 249576 152804 249582 152856
rect 255498 152804 255504 152856
rect 255556 152844 255562 152856
rect 257246 152844 257252 152856
rect 255556 152816 257252 152844
rect 255556 152804 255562 152816
rect 257246 152804 257252 152816
rect 257304 152804 257310 152856
rect 258074 152804 258080 152856
rect 258132 152844 258138 152856
rect 316310 152844 316316 152856
rect 258132 152816 316316 152844
rect 258132 152804 258138 152816
rect 316310 152804 316316 152816
rect 316368 152804 316374 152856
rect 317138 152804 317144 152856
rect 317196 152844 317202 152856
rect 318242 152844 318248 152856
rect 317196 152816 318248 152844
rect 317196 152804 317202 152816
rect 318242 152804 318248 152816
rect 318300 152804 318306 152856
rect 322934 152804 322940 152856
rect 322992 152844 322998 152856
rect 366358 152844 366364 152856
rect 322992 152816 366364 152844
rect 322992 152804 322998 152816
rect 366358 152804 366364 152816
rect 366416 152804 366422 152856
rect 367554 152804 367560 152856
rect 367612 152844 367618 152856
rect 367612 152816 388392 152844
rect 367612 152804 367618 152816
rect 26326 152736 26332 152788
rect 26384 152776 26390 152788
rect 139118 152776 139124 152788
rect 26384 152748 139124 152776
rect 26384 152736 26390 152748
rect 139118 152736 139124 152748
rect 139176 152736 139182 152788
rect 139210 152736 139216 152788
rect 139268 152776 139274 152788
rect 149422 152776 149428 152788
rect 139268 152748 149428 152776
rect 139268 152736 139274 152748
rect 149422 152736 149428 152748
rect 149480 152736 149486 152788
rect 152826 152736 152832 152788
rect 152884 152776 152890 152788
rect 234154 152776 234160 152788
rect 152884 152748 234160 152776
rect 152884 152736 152890 152748
rect 234154 152736 234160 152748
rect 234212 152736 234218 152788
rect 237374 152736 237380 152788
rect 237432 152776 237438 152788
rect 300946 152776 300952 152788
rect 237432 152748 300952 152776
rect 237432 152736 237438 152748
rect 300946 152736 300952 152748
rect 301004 152736 301010 152788
rect 303522 152736 303528 152788
rect 303580 152776 303586 152788
rect 350994 152776 351000 152788
rect 303580 152748 351000 152776
rect 303580 152736 303586 152748
rect 350994 152736 351000 152748
rect 351052 152736 351058 152788
rect 351914 152736 351920 152788
rect 351972 152776 351978 152788
rect 388254 152776 388260 152788
rect 351972 152748 388260 152776
rect 351972 152736 351978 152748
rect 388254 152736 388260 152748
rect 388312 152736 388318 152788
rect 388364 152776 388392 152816
rect 395890 152804 395896 152856
rect 395948 152844 395954 152856
rect 395948 152816 402974 152844
rect 395948 152804 395954 152816
rect 400398 152776 400404 152788
rect 388364 152748 400404 152776
rect 400398 152736 400404 152748
rect 400456 152736 400462 152788
rect 402946 152776 402974 152816
rect 405918 152804 405924 152856
rect 405976 152844 405982 152856
rect 429286 152844 429292 152856
rect 405976 152816 429292 152844
rect 405976 152804 405982 152816
rect 429286 152804 429292 152816
rect 429344 152804 429350 152856
rect 429562 152804 429568 152856
rect 429620 152844 429626 152856
rect 441062 152844 441068 152856
rect 429620 152816 441068 152844
rect 429620 152804 429626 152816
rect 441062 152804 441068 152816
rect 441120 152804 441126 152856
rect 446674 152844 446680 152856
rect 441172 152816 446680 152844
rect 421650 152776 421656 152788
rect 402946 152748 421656 152776
rect 421650 152736 421656 152748
rect 421708 152736 421714 152788
rect 428642 152736 428648 152788
rect 428700 152776 428706 152788
rect 441172 152776 441200 152816
rect 446674 152804 446680 152816
rect 446732 152804 446738 152856
rect 447686 152804 447692 152856
rect 447744 152844 447750 152856
rect 461394 152844 461400 152856
rect 447744 152816 461400 152844
rect 447744 152804 447750 152816
rect 461394 152804 461400 152816
rect 461452 152804 461458 152856
rect 466546 152804 466552 152856
rect 466604 152844 466610 152856
rect 470410 152844 470416 152856
rect 466604 152816 470416 152844
rect 466604 152804 466610 152816
rect 470410 152804 470416 152816
rect 470468 152804 470474 152856
rect 491754 152804 491760 152856
rect 491812 152844 491818 152856
rect 495434 152844 495440 152856
rect 491812 152816 495440 152844
rect 491812 152804 491818 152816
rect 495434 152804 495440 152816
rect 495492 152804 495498 152856
rect 428700 152748 441200 152776
rect 428700 152736 428706 152748
rect 441246 152736 441252 152788
rect 441304 152776 441310 152788
rect 444834 152776 444840 152788
rect 441304 152748 444840 152776
rect 441304 152736 441310 152748
rect 444834 152736 444840 152748
rect 444892 152736 444898 152788
rect 448882 152736 448888 152788
rect 448940 152776 448946 152788
rect 462682 152776 462688 152788
rect 448940 152748 462688 152776
rect 448940 152736 448946 152748
rect 462682 152736 462688 152748
rect 462740 152736 462746 152788
rect 86126 152668 86132 152720
rect 86184 152708 86190 152720
rect 185302 152708 185308 152720
rect 86184 152680 185308 152708
rect 86184 152668 86190 152680
rect 185302 152668 185308 152680
rect 185360 152668 185366 152720
rect 190546 152668 190552 152720
rect 190604 152708 190610 152720
rect 264974 152708 264980 152720
rect 190604 152680 264980 152708
rect 190604 152668 190610 152680
rect 264974 152668 264980 152680
rect 265032 152668 265038 152720
rect 270862 152668 270868 152720
rect 270920 152708 270926 152720
rect 326614 152708 326620 152720
rect 270920 152680 326620 152708
rect 270920 152668 270926 152680
rect 326614 152668 326620 152680
rect 326672 152668 326678 152720
rect 329834 152668 329840 152720
rect 329892 152708 329898 152720
rect 361758 152708 361764 152720
rect 329892 152680 361764 152708
rect 329892 152668 329898 152680
rect 361758 152668 361764 152680
rect 361816 152668 361822 152720
rect 367002 152708 367008 152720
rect 364628 152680 367008 152708
rect 31754 152600 31760 152652
rect 31812 152640 31818 152652
rect 143626 152640 143632 152652
rect 31812 152612 143632 152640
rect 31812 152600 31818 152612
rect 143626 152600 143632 152612
rect 143684 152600 143690 152652
rect 144454 152600 144460 152652
rect 144512 152640 144518 152652
rect 159634 152640 159640 152652
rect 144512 152612 159640 152640
rect 144512 152600 144518 152612
rect 159634 152600 159640 152612
rect 159692 152600 159698 152652
rect 163498 152600 163504 152652
rect 163556 152640 163562 152652
rect 244366 152640 244372 152652
rect 163556 152612 244372 152640
rect 163556 152600 163562 152612
rect 244366 152600 244372 152612
rect 244424 152600 244430 152652
rect 245746 152600 245752 152652
rect 245804 152640 245810 152652
rect 306006 152640 306012 152652
rect 245804 152612 306012 152640
rect 245804 152600 245810 152612
rect 306006 152600 306012 152612
rect 306064 152600 306070 152652
rect 310606 152600 310612 152652
rect 310664 152640 310670 152652
rect 356790 152640 356796 152652
rect 310664 152612 356796 152640
rect 310664 152600 310670 152612
rect 356790 152600 356796 152612
rect 356848 152600 356854 152652
rect 357526 152600 357532 152652
rect 357584 152640 357590 152652
rect 359366 152640 359372 152652
rect 357584 152612 359372 152640
rect 357584 152600 357590 152612
rect 359366 152600 359372 152612
rect 359424 152600 359430 152652
rect 363230 152600 363236 152652
rect 363288 152640 363294 152652
rect 364518 152640 364524 152652
rect 363288 152612 364524 152640
rect 363288 152600 363294 152612
rect 364518 152600 364524 152612
rect 364576 152600 364582 152652
rect 18046 152532 18052 152584
rect 18104 152572 18110 152584
rect 133322 152572 133328 152584
rect 18104 152544 133328 152572
rect 18104 152532 18110 152544
rect 133322 152532 133328 152544
rect 133380 152532 133386 152584
rect 137278 152532 137284 152584
rect 137336 152572 137342 152584
rect 144270 152572 144276 152584
rect 137336 152544 144276 152572
rect 137336 152532 137342 152544
rect 144270 152532 144276 152544
rect 144328 152532 144334 152584
rect 146938 152532 146944 152584
rect 146996 152572 147002 152584
rect 157058 152572 157064 152584
rect 146996 152544 157064 152572
rect 146996 152532 147002 152544
rect 157058 152532 157064 152544
rect 157116 152532 157122 152584
rect 157334 152532 157340 152584
rect 157392 152572 157398 152584
rect 239306 152572 239312 152584
rect 157392 152544 239312 152572
rect 157392 152532 157398 152544
rect 239306 152532 239312 152544
rect 239364 152532 239370 152584
rect 240318 152532 240324 152584
rect 240376 152572 240382 152584
rect 241882 152572 241888 152584
rect 240376 152544 241888 152572
rect 240376 152532 240382 152544
rect 241882 152532 241888 152544
rect 241940 152532 241946 152584
rect 242986 152532 242992 152584
rect 243044 152572 243050 152584
rect 246942 152572 246948 152584
rect 243044 152544 246948 152572
rect 243044 152532 243050 152544
rect 246942 152532 246948 152544
rect 247000 152532 247006 152584
rect 249978 152532 249984 152584
rect 250036 152572 250042 152584
rect 310514 152572 310520 152584
rect 250036 152544 310520 152572
rect 250036 152532 250042 152544
rect 310514 152532 310520 152544
rect 310572 152532 310578 152584
rect 311894 152532 311900 152584
rect 311952 152572 311958 152584
rect 357434 152572 357440 152584
rect 311952 152544 357440 152572
rect 311952 152532 311958 152544
rect 357434 152532 357440 152544
rect 357492 152532 357498 152584
rect 359458 152532 359464 152584
rect 359516 152572 359522 152584
rect 364628 152572 364656 152680
rect 367002 152668 367008 152680
rect 367060 152668 367066 152720
rect 379054 152668 379060 152720
rect 379112 152708 379118 152720
rect 388438 152708 388444 152720
rect 379112 152680 388444 152708
rect 379112 152668 379118 152680
rect 388438 152668 388444 152680
rect 388496 152668 388502 152720
rect 388530 152668 388536 152720
rect 388588 152708 388594 152720
rect 407482 152708 407488 152720
rect 388588 152680 407488 152708
rect 388588 152668 388594 152680
rect 407482 152668 407488 152680
rect 407540 152668 407546 152720
rect 409046 152668 409052 152720
rect 409104 152708 409110 152720
rect 431862 152708 431868 152720
rect 409104 152680 431868 152708
rect 409104 152668 409110 152680
rect 431862 152668 431868 152680
rect 431920 152668 431926 152720
rect 431954 152668 431960 152720
rect 432012 152708 432018 152720
rect 434438 152708 434444 152720
rect 432012 152680 434444 152708
rect 432012 152668 432018 152680
rect 434438 152668 434444 152680
rect 434496 152668 434502 152720
rect 434530 152668 434536 152720
rect 434588 152708 434594 152720
rect 446950 152708 446956 152720
rect 434588 152680 446956 152708
rect 434588 152668 434594 152680
rect 446950 152668 446956 152680
rect 447008 152668 447014 152720
rect 447042 152668 447048 152720
rect 447100 152708 447106 152720
rect 452470 152708 452476 152720
rect 447100 152680 452476 152708
rect 447100 152668 447106 152680
rect 452470 152668 452476 152680
rect 452528 152668 452534 152720
rect 365070 152600 365076 152652
rect 365128 152640 365134 152652
rect 393406 152640 393412 152652
rect 365128 152612 393412 152640
rect 365128 152600 365134 152612
rect 393406 152600 393412 152612
rect 393464 152600 393470 152652
rect 401870 152600 401876 152652
rect 401928 152640 401934 152652
rect 426802 152640 426808 152652
rect 401928 152612 426808 152640
rect 401928 152600 401934 152612
rect 426802 152600 426808 152612
rect 426860 152600 426866 152652
rect 429194 152600 429200 152652
rect 429252 152640 429258 152652
rect 447318 152640 447324 152652
rect 429252 152612 447324 152640
rect 429252 152600 429258 152612
rect 447318 152600 447324 152612
rect 447376 152600 447382 152652
rect 447410 152600 447416 152652
rect 447468 152640 447474 152652
rect 451182 152640 451188 152652
rect 447468 152612 451188 152640
rect 447468 152600 447474 152612
rect 451182 152600 451188 152612
rect 451240 152600 451246 152652
rect 359516 152544 364656 152572
rect 359516 152532 359522 152544
rect 367094 152532 367100 152584
rect 367152 152572 367158 152584
rect 394694 152572 394700 152584
rect 367152 152544 394700 152572
rect 367152 152532 367158 152544
rect 394694 152532 394700 152544
rect 394752 152532 394758 152584
rect 397546 152532 397552 152584
rect 397604 152572 397610 152584
rect 422846 152572 422852 152584
rect 397604 152544 422852 152572
rect 397604 152532 397610 152544
rect 422846 152532 422852 152544
rect 422904 152532 422910 152584
rect 430574 152532 430580 152584
rect 430632 152572 430638 152584
rect 430632 152544 442212 152572
rect 430632 152532 430638 152544
rect 12434 152464 12440 152516
rect 12492 152504 12498 152516
rect 128814 152504 128820 152516
rect 12492 152476 128820 152504
rect 12492 152464 12498 152476
rect 128814 152464 128820 152476
rect 128872 152464 128878 152516
rect 129734 152464 129740 152516
rect 129792 152504 129798 152516
rect 218698 152504 218704 152516
rect 129792 152476 218704 152504
rect 129792 152464 129798 152476
rect 218698 152464 218704 152476
rect 218756 152464 218762 152516
rect 223758 152464 223764 152516
rect 223816 152504 223822 152516
rect 289998 152504 290004 152516
rect 223816 152476 290004 152504
rect 223816 152464 223822 152476
rect 289998 152464 290004 152476
rect 290056 152464 290062 152516
rect 297634 152464 297640 152516
rect 297692 152504 297698 152516
rect 346486 152504 346492 152516
rect 297692 152476 346492 152504
rect 297692 152464 297698 152476
rect 346486 152464 346492 152476
rect 346544 152464 346550 152516
rect 347774 152464 347780 152516
rect 347832 152504 347838 152516
rect 385034 152504 385040 152516
rect 347832 152476 385040 152504
rect 347832 152464 347838 152476
rect 385034 152464 385040 152476
rect 385092 152464 385098 152516
rect 394234 152464 394240 152516
rect 394292 152504 394298 152516
rect 420362 152504 420368 152516
rect 394292 152476 420368 152504
rect 394292 152464 394298 152476
rect 420362 152464 420368 152476
rect 420420 152464 420426 152516
rect 423398 152464 423404 152516
rect 423456 152504 423462 152516
rect 427078 152504 427084 152516
rect 423456 152476 427084 152504
rect 423456 152464 423462 152476
rect 427078 152464 427084 152476
rect 427136 152464 427142 152516
rect 433794 152504 433800 152516
rect 427786 152476 433800 152504
rect 81434 152396 81440 152448
rect 81492 152436 81498 152448
rect 175090 152436 175096 152448
rect 81492 152408 175096 152436
rect 81492 152396 81498 152408
rect 175090 152396 175096 152408
rect 175148 152396 175154 152448
rect 176746 152396 176752 152448
rect 176804 152436 176810 152448
rect 254670 152436 254676 152448
rect 176804 152408 254676 152436
rect 176804 152396 176810 152408
rect 254670 152396 254676 152408
rect 254728 152396 254734 152448
rect 256694 152396 256700 152448
rect 256752 152436 256758 152448
rect 315666 152436 315672 152448
rect 256752 152408 315672 152436
rect 256752 152396 256758 152408
rect 315666 152396 315672 152408
rect 315724 152396 315730 152448
rect 317046 152396 317052 152448
rect 317104 152436 317110 152448
rect 361298 152436 361304 152448
rect 317104 152408 361304 152436
rect 317104 152396 317110 152408
rect 361298 152396 361304 152408
rect 361356 152396 361362 152448
rect 361758 152396 361764 152448
rect 361816 152436 361822 152448
rect 371510 152436 371516 152448
rect 361816 152408 371516 152436
rect 361816 152396 361822 152408
rect 371510 152396 371516 152408
rect 371568 152396 371574 152448
rect 398466 152436 398472 152448
rect 371620 152408 398472 152436
rect 89714 152328 89720 152380
rect 89772 152368 89778 152380
rect 180242 152368 180248 152380
rect 89772 152340 180248 152368
rect 89772 152328 89778 152340
rect 180242 152328 180248 152340
rect 180300 152328 180306 152380
rect 185026 152328 185032 152380
rect 185084 152368 185090 152380
rect 259822 152368 259828 152380
rect 185084 152340 259828 152368
rect 185084 152328 185090 152340
rect 259822 152328 259828 152340
rect 259880 152328 259886 152380
rect 263594 152328 263600 152380
rect 263652 152368 263658 152380
rect 320818 152368 320824 152380
rect 263652 152340 320824 152368
rect 263652 152328 263658 152340
rect 320818 152328 320824 152340
rect 320876 152328 320882 152380
rect 321554 152328 321560 152380
rect 321612 152368 321618 152380
rect 323394 152368 323400 152380
rect 321612 152340 323400 152368
rect 321612 152328 321618 152340
rect 323394 152328 323400 152340
rect 323452 152328 323458 152380
rect 324590 152328 324596 152380
rect 324648 152368 324654 152380
rect 367646 152368 367652 152380
rect 324648 152340 367652 152368
rect 324648 152328 324654 152340
rect 367646 152328 367652 152340
rect 367704 152328 367710 152380
rect 367738 152328 367744 152380
rect 367796 152368 367802 152380
rect 371620 152368 371648 152408
rect 398466 152396 398472 152408
rect 398524 152396 398530 152448
rect 398834 152396 398840 152448
rect 398892 152436 398898 152448
rect 410702 152436 410708 152448
rect 398892 152408 410708 152436
rect 398892 152396 398898 152408
rect 410702 152396 410708 152408
rect 410760 152396 410766 152448
rect 413738 152396 413744 152448
rect 413796 152436 413802 152448
rect 427786 152436 427814 152476
rect 433794 152464 433800 152476
rect 433852 152464 433858 152516
rect 434438 152464 434444 152516
rect 434496 152504 434502 152516
rect 435726 152504 435732 152516
rect 434496 152476 435732 152504
rect 434496 152464 434502 152476
rect 435726 152464 435732 152476
rect 435784 152464 435790 152516
rect 442074 152504 442080 152516
rect 437446 152476 442080 152504
rect 413796 152408 427814 152436
rect 413796 152396 413802 152408
rect 429470 152396 429476 152448
rect 429528 152436 429534 152448
rect 437446 152436 437474 152476
rect 442074 152464 442080 152476
rect 442132 152464 442138 152516
rect 429528 152408 437474 152436
rect 429528 152396 429534 152408
rect 367796 152340 371648 152368
rect 367796 152328 367802 152340
rect 371786 152328 371792 152380
rect 371844 152368 371850 152380
rect 403618 152368 403624 152380
rect 371844 152340 403624 152368
rect 371844 152328 371850 152340
rect 403618 152328 403624 152340
rect 403676 152328 403682 152380
rect 403894 152328 403900 152380
rect 403952 152368 403958 152380
rect 418430 152368 418436 152380
rect 403952 152340 418436 152368
rect 403952 152328 403958 152340
rect 418430 152328 418436 152340
rect 418488 152328 418494 152380
rect 421926 152328 421932 152380
rect 421984 152368 421990 152380
rect 429746 152368 429752 152380
rect 421984 152340 429752 152368
rect 421984 152328 421990 152340
rect 429746 152328 429752 152340
rect 429804 152328 429810 152380
rect 441522 152368 441528 152380
rect 429948 152340 441528 152368
rect 76466 152260 76472 152312
rect 76524 152300 76530 152312
rect 162210 152300 162216 152312
rect 76524 152272 162216 152300
rect 76524 152260 76530 152272
rect 162210 152260 162216 152272
rect 162268 152260 162274 152312
rect 166994 152260 167000 152312
rect 167052 152300 167058 152312
rect 182818 152300 182824 152312
rect 167052 152272 182824 152300
rect 167052 152260 167058 152272
rect 182818 152260 182824 152272
rect 182876 152260 182882 152312
rect 186406 152260 186412 152312
rect 186464 152300 186470 152312
rect 205910 152300 205916 152312
rect 186464 152272 205916 152300
rect 186464 152260 186470 152272
rect 205910 152260 205916 152272
rect 205968 152260 205974 152312
rect 230750 152260 230756 152312
rect 230808 152300 230814 152312
rect 290642 152300 290648 152312
rect 230808 152272 290648 152300
rect 230808 152260 230814 152272
rect 290642 152260 290648 152272
rect 290700 152260 290706 152312
rect 293954 152260 293960 152312
rect 294012 152300 294018 152312
rect 341978 152300 341984 152312
rect 294012 152272 341984 152300
rect 294012 152260 294018 152272
rect 341978 152260 341984 152272
rect 342036 152260 342042 152312
rect 345014 152260 345020 152312
rect 345072 152300 345078 152312
rect 383102 152300 383108 152312
rect 345072 152272 367692 152300
rect 345072 152260 345078 152272
rect 33594 152192 33600 152244
rect 33652 152232 33658 152244
rect 109586 152232 109592 152244
rect 33652 152204 109592 152232
rect 33652 152192 33658 152204
rect 109586 152192 109592 152204
rect 109644 152192 109650 152244
rect 109678 152192 109684 152244
rect 109736 152232 109742 152244
rect 130746 152232 130752 152244
rect 109736 152204 130752 152232
rect 109736 152192 109742 152204
rect 130746 152192 130752 152204
rect 130804 152192 130810 152244
rect 135162 152192 135168 152244
rect 135220 152232 135226 152244
rect 139210 152232 139216 152244
rect 135220 152204 139216 152232
rect 135220 152192 135226 152204
rect 139210 152192 139216 152204
rect 139268 152192 139274 152244
rect 139302 152192 139308 152244
rect 139360 152232 139366 152244
rect 141786 152232 141792 152244
rect 139360 152204 141792 152232
rect 139360 152192 139366 152204
rect 141786 152192 141792 152204
rect 141844 152192 141850 152244
rect 143534 152192 143540 152244
rect 143592 152232 143598 152244
rect 229002 152232 229008 152244
rect 143592 152204 229008 152232
rect 143592 152192 143598 152204
rect 229002 152192 229008 152204
rect 229060 152192 229066 152244
rect 246114 152192 246120 152244
rect 246172 152232 246178 152244
rect 305362 152232 305368 152244
rect 246172 152204 305368 152232
rect 246172 152192 246178 152204
rect 305362 152192 305368 152204
rect 305420 152192 305426 152244
rect 319162 152192 319168 152244
rect 319220 152232 319226 152244
rect 362586 152232 362592 152244
rect 319220 152204 362592 152232
rect 319220 152192 319226 152204
rect 362586 152192 362592 152204
rect 362644 152192 362650 152244
rect 367664 152232 367692 152272
rect 369826 152272 383108 152300
rect 369826 152232 369854 152272
rect 383102 152260 383108 152272
rect 383160 152260 383166 152312
rect 383194 152260 383200 152312
rect 383252 152300 383258 152312
rect 389542 152300 389548 152312
rect 383252 152272 389548 152300
rect 383252 152260 383258 152272
rect 389542 152260 389548 152272
rect 389600 152260 389606 152312
rect 390554 152260 390560 152312
rect 390612 152300 390618 152312
rect 415210 152300 415216 152312
rect 390612 152272 415216 152300
rect 390612 152260 390618 152272
rect 415210 152260 415216 152272
rect 415268 152260 415274 152312
rect 415670 152260 415676 152312
rect 415728 152300 415734 152312
rect 419074 152300 419080 152312
rect 415728 152272 419080 152300
rect 415728 152260 415734 152272
rect 419074 152260 419080 152272
rect 419132 152260 419138 152312
rect 367664 152204 369854 152232
rect 370682 152192 370688 152244
rect 370740 152232 370746 152244
rect 402330 152232 402336 152244
rect 370740 152204 402336 152232
rect 370740 152192 370746 152204
rect 402330 152192 402336 152204
rect 402388 152192 402394 152244
rect 408862 152192 408868 152244
rect 408920 152232 408926 152244
rect 428642 152232 428648 152244
rect 408920 152204 428648 152232
rect 408920 152192 408926 152204
rect 428642 152192 428648 152204
rect 428700 152192 428706 152244
rect 429746 152192 429752 152244
rect 429804 152232 429810 152244
rect 429948 152232 429976 152340
rect 441522 152328 441528 152340
rect 441580 152328 441586 152380
rect 442184 152368 442212 152544
rect 445386 152532 445392 152584
rect 445444 152572 445450 152584
rect 459462 152572 459468 152584
rect 445444 152544 459468 152572
rect 445444 152532 445450 152544
rect 459462 152532 459468 152544
rect 459520 152532 459526 152584
rect 442350 152464 442356 152516
rect 442408 152504 442414 152516
rect 453114 152504 453120 152516
rect 442408 152476 453120 152504
rect 442408 152464 442414 152476
rect 453114 152464 453120 152476
rect 453172 152464 453178 152516
rect 488534 152464 488540 152516
rect 488592 152504 488598 152516
rect 492858 152504 492864 152516
rect 488592 152476 492864 152504
rect 488592 152464 488598 152476
rect 492858 152464 492864 152476
rect 492916 152464 492922 152516
rect 442258 152396 442264 152448
rect 442316 152436 442322 152448
rect 444742 152436 444748 152448
rect 442316 152408 444748 152436
rect 442316 152396 442322 152408
rect 444742 152396 444748 152408
rect 444800 152396 444806 152448
rect 444834 152396 444840 152448
rect 444892 152436 444898 152448
rect 456334 152436 456340 152448
rect 444892 152408 456340 152436
rect 444892 152396 444898 152408
rect 456334 152396 456340 152408
rect 456392 152396 456398 152448
rect 448606 152368 448612 152380
rect 442184 152340 448612 152368
rect 448606 152328 448612 152340
rect 448664 152328 448670 152380
rect 432690 152260 432696 152312
rect 432748 152300 432754 152312
rect 444098 152300 444104 152312
rect 432748 152272 444104 152300
rect 432748 152260 432754 152272
rect 444098 152260 444104 152272
rect 444156 152260 444162 152312
rect 444558 152260 444564 152312
rect 444616 152300 444622 152312
rect 458910 152300 458916 152312
rect 444616 152272 458916 152300
rect 444616 152260 444622 152272
rect 458910 152260 458916 152272
rect 458968 152260 458974 152312
rect 429804 152204 429976 152232
rect 429804 152192 429810 152204
rect 432782 152192 432788 152244
rect 432840 152232 432846 152244
rect 449250 152232 449256 152244
rect 432840 152204 449256 152232
rect 432840 152192 432846 152204
rect 449250 152192 449256 152204
rect 449308 152192 449314 152244
rect 69658 152124 69664 152176
rect 69716 152164 69722 152176
rect 154482 152164 154488 152176
rect 69716 152136 154488 152164
rect 69716 152124 69722 152136
rect 154482 152124 154488 152136
rect 154540 152124 154546 152176
rect 154574 152124 154580 152176
rect 154632 152164 154638 152176
rect 169938 152164 169944 152176
rect 154632 152136 169944 152164
rect 154632 152124 154638 152136
rect 169938 152124 169944 152136
rect 169996 152124 170002 152176
rect 173986 152124 173992 152176
rect 174044 152164 174050 152176
rect 193030 152164 193036 152176
rect 174044 152136 193036 152164
rect 174044 152124 174050 152136
rect 193030 152124 193036 152136
rect 193088 152124 193094 152176
rect 229370 152124 229376 152176
rect 229428 152164 229434 152176
rect 287422 152164 287428 152176
rect 229428 152136 287428 152164
rect 229428 152124 229434 152136
rect 287422 152124 287428 152136
rect 287480 152124 287486 152176
rect 295334 152124 295340 152176
rect 295392 152164 295398 152176
rect 297726 152164 297732 152176
rect 295392 152136 297732 152164
rect 295392 152124 295398 152136
rect 297726 152124 297732 152136
rect 297784 152124 297790 152176
rect 299474 152124 299480 152176
rect 299532 152164 299538 152176
rect 347130 152164 347136 152176
rect 299532 152136 347136 152164
rect 299532 152124 299538 152136
rect 347130 152124 347136 152136
rect 347188 152124 347194 152176
rect 350534 152124 350540 152176
rect 350592 152164 350598 152176
rect 386966 152164 386972 152176
rect 350592 152136 386972 152164
rect 350592 152124 350598 152136
rect 386966 152124 386972 152136
rect 387024 152124 387030 152176
rect 388530 152164 388536 152176
rect 388364 152136 388536 152164
rect 19794 152056 19800 152108
rect 19852 152096 19858 152108
rect 99926 152096 99932 152108
rect 19852 152068 99932 152096
rect 19852 152056 19858 152068
rect 99926 152056 99932 152068
rect 99984 152056 99990 152108
rect 109034 152056 109040 152108
rect 109092 152096 109098 152108
rect 128170 152096 128176 152108
rect 109092 152068 128176 152096
rect 109092 152056 109098 152068
rect 128170 152056 128176 152068
rect 128228 152056 128234 152108
rect 128446 152056 128452 152108
rect 128504 152096 128510 152108
rect 213546 152096 213552 152108
rect 128504 152068 213552 152096
rect 128504 152056 128510 152068
rect 213546 152056 213552 152068
rect 213604 152056 213610 152108
rect 252922 152056 252928 152108
rect 252980 152096 252986 152108
rect 311158 152096 311164 152108
rect 252980 152068 311164 152096
rect 252980 152056 252986 152068
rect 311158 152056 311164 152068
rect 311216 152056 311222 152108
rect 318886 152056 318892 152108
rect 318944 152096 318950 152108
rect 361942 152096 361948 152108
rect 318944 152068 361948 152096
rect 318944 152056 318950 152068
rect 361942 152056 361948 152068
rect 362000 152056 362006 152108
rect 364794 152056 364800 152108
rect 364852 152096 364858 152108
rect 367738 152096 367744 152108
rect 364852 152068 367744 152096
rect 364852 152056 364858 152068
rect 367738 152056 367744 152068
rect 367796 152056 367802 152108
rect 377766 152056 377772 152108
rect 377824 152096 377830 152108
rect 381814 152096 381820 152108
rect 377824 152068 381820 152096
rect 377824 152056 377830 152068
rect 381814 152056 381820 152068
rect 381872 152056 381878 152108
rect 388364 152096 388392 152136
rect 388530 152124 388536 152136
rect 388588 152124 388594 152176
rect 388622 152124 388628 152176
rect 388680 152164 388686 152176
rect 410058 152164 410064 152176
rect 388680 152136 410064 152164
rect 388680 152124 388686 152136
rect 410058 152124 410064 152136
rect 410116 152124 410122 152176
rect 411254 152124 411260 152176
rect 411312 152164 411318 152176
rect 431218 152164 431224 152176
rect 411312 152136 431224 152164
rect 411312 152124 411318 152136
rect 431218 152124 431224 152136
rect 431276 152124 431282 152176
rect 433426 152124 433432 152176
rect 433484 152164 433490 152176
rect 450538 152164 450544 152176
rect 433484 152136 450544 152164
rect 433484 152124 433490 152136
rect 450538 152124 450544 152136
rect 450596 152124 450602 152176
rect 408126 152096 408132 152108
rect 382016 152068 388392 152096
rect 388456 152068 408132 152096
rect 63494 151988 63500 152040
rect 63552 152028 63558 152040
rect 146846 152028 146852 152040
rect 63552 152000 146852 152028
rect 63552 151988 63558 152000
rect 146846 151988 146852 152000
rect 146904 151988 146910 152040
rect 158806 151988 158812 152040
rect 158864 152028 158870 152040
rect 172514 152028 172520 152040
rect 158864 152000 172520 152028
rect 158864 151988 158870 152000
rect 172514 151988 172520 152000
rect 172572 151988 172578 152040
rect 183094 151988 183100 152040
rect 183152 152028 183158 152040
rect 198182 152028 198188 152040
rect 183152 152000 198188 152028
rect 183152 151988 183158 152000
rect 198182 151988 198188 152000
rect 198240 151988 198246 152040
rect 264146 151988 264152 152040
rect 264204 152028 264210 152040
rect 321462 152028 321468 152040
rect 264204 152000 321468 152028
rect 264204 151988 264210 152000
rect 321462 151988 321468 152000
rect 321520 151988 321526 152040
rect 331306 151988 331312 152040
rect 331364 152028 331370 152040
rect 334342 152028 334348 152040
rect 331364 152000 334348 152028
rect 331364 151988 331370 152000
rect 334342 151988 334348 152000
rect 334400 151988 334406 152040
rect 359458 152028 359464 152040
rect 334452 152000 359464 152028
rect 75822 151920 75828 151972
rect 75880 151960 75886 151972
rect 75880 151932 84194 151960
rect 75880 151920 75886 151932
rect 74810 151852 74816 151904
rect 74868 151892 74874 151904
rect 82078 151892 82084 151904
rect 74868 151864 82084 151892
rect 74868 151852 74874 151864
rect 82078 151852 82084 151864
rect 82136 151852 82142 151904
rect 84166 151892 84194 151932
rect 105814 151920 105820 151972
rect 105872 151960 105878 151972
rect 110322 151960 110328 151972
rect 105872 151932 110328 151960
rect 105872 151920 105878 151932
rect 110322 151920 110328 151932
rect 110380 151920 110386 151972
rect 127250 151920 127256 151972
rect 127308 151960 127314 151972
rect 135898 151960 135904 151972
rect 127308 151932 135904 151960
rect 127308 151920 127314 151932
rect 135898 151920 135904 151932
rect 135956 151920 135962 151972
rect 142890 151920 142896 151972
rect 142948 151960 142954 151972
rect 223850 151960 223856 151972
rect 142948 151932 223856 151960
rect 142948 151920 142954 151932
rect 223850 151920 223856 151932
rect 223908 151920 223914 151972
rect 278038 151920 278044 151972
rect 278096 151960 278102 151972
rect 331766 151960 331772 151972
rect 278096 151932 331772 151960
rect 278096 151920 278102 151932
rect 331766 151920 331772 151932
rect 331824 151920 331830 151972
rect 151906 151892 151912 151904
rect 84166 151864 151912 151892
rect 151906 151852 151912 151864
rect 151964 151852 151970 151904
rect 164510 151852 164516 151904
rect 164568 151892 164574 151904
rect 164568 151864 171134 151892
rect 164568 151852 164574 151864
rect 71406 151784 71412 151836
rect 71464 151824 71470 151836
rect 91002 151824 91008 151836
rect 71464 151796 91008 151824
rect 71464 151784 71470 151796
rect 91002 151784 91008 151796
rect 91060 151784 91066 151836
rect 102134 151784 102140 151836
rect 102192 151824 102198 151836
rect 167362 151824 167368 151836
rect 102192 151796 167368 151824
rect 102192 151784 102198 151796
rect 167362 151784 167368 151796
rect 167420 151784 167426 151836
rect 171106 151824 171134 151864
rect 173250 151852 173256 151904
rect 173308 151892 173314 151904
rect 187878 151892 187884 151904
rect 173308 151864 187884 151892
rect 173308 151852 173314 151864
rect 187878 151852 187884 151864
rect 187936 151852 187942 151904
rect 219894 151852 219900 151904
rect 219952 151892 219958 151904
rect 275186 151892 275192 151904
rect 219952 151864 275192 151892
rect 219952 151852 219958 151864
rect 275186 151852 275192 151864
rect 275244 151852 275250 151904
rect 276106 151852 276112 151904
rect 276164 151892 276170 151904
rect 277762 151892 277768 151904
rect 276164 151864 277768 151892
rect 276164 151852 276170 151864
rect 277762 151852 277768 151864
rect 277820 151852 277826 151904
rect 280154 151852 280160 151904
rect 280212 151892 280218 151904
rect 331122 151892 331128 151904
rect 280212 151864 331128 151892
rect 280212 151852 280218 151864
rect 331122 151852 331128 151864
rect 331180 151852 331186 151904
rect 334452 151892 334480 152000
rect 359458 151988 359464 152000
rect 359516 151988 359522 152040
rect 360194 151988 360200 152040
rect 360252 152028 360258 152040
rect 367094 152028 367100 152040
rect 360252 152000 367100 152028
rect 360252 151988 360258 152000
rect 367094 151988 367100 152000
rect 367152 151988 367158 152040
rect 372798 151960 372804 151972
rect 335326 151932 372804 151960
rect 331232 151864 334480 151892
rect 177666 151824 177672 151836
rect 171106 151796 177672 151824
rect 177666 151784 177672 151796
rect 177724 151784 177730 151836
rect 215386 151784 215392 151836
rect 215444 151824 215450 151836
rect 270126 151824 270132 151836
rect 215444 151796 270132 151824
rect 215444 151784 215450 151796
rect 270126 151784 270132 151796
rect 270184 151784 270190 151836
rect 273346 151784 273352 151836
rect 273404 151824 273410 151836
rect 325970 151824 325976 151836
rect 273404 151796 325976 151824
rect 273404 151784 273410 151796
rect 325970 151784 325976 151796
rect 326028 151784 326034 151836
rect 328362 151784 328368 151836
rect 328420 151824 328426 151836
rect 331232 151824 331260 151864
rect 334526 151852 334532 151904
rect 334584 151892 334590 151904
rect 335326 151892 335354 151932
rect 372798 151920 372804 151932
rect 372856 151920 372862 151972
rect 376754 151920 376760 151972
rect 376812 151960 376818 151972
rect 382016 151960 382044 152068
rect 388456 152028 388484 152068
rect 408126 152056 408132 152068
rect 408184 152056 408190 152108
rect 418246 152056 418252 152108
rect 418304 152096 418310 152108
rect 424226 152096 424232 152108
rect 418304 152068 424232 152096
rect 418304 152056 418310 152068
rect 424226 152056 424232 152068
rect 424284 152056 424290 152108
rect 442166 152096 442172 152108
rect 434686 152068 442172 152096
rect 376812 151932 382044 151960
rect 383626 152000 388484 152028
rect 376812 151920 376818 151932
rect 334584 151864 335354 151892
rect 334584 151852 334590 151864
rect 339494 151852 339500 151904
rect 339552 151892 339558 151904
rect 377306 151892 377312 151904
rect 339552 151864 377312 151892
rect 339552 151852 339558 151864
rect 377306 151852 377312 151864
rect 377364 151852 377370 151904
rect 378226 151852 378232 151904
rect 378284 151892 378290 151904
rect 383626 151892 383654 152000
rect 388714 151988 388720 152040
rect 388772 152028 388778 152040
rect 404906 152028 404912 152040
rect 388772 152000 404912 152028
rect 388772 151988 388778 152000
rect 404906 151988 404912 152000
rect 404964 151988 404970 152040
rect 407574 151988 407580 152040
rect 407632 152028 407638 152040
rect 426158 152028 426164 152040
rect 407632 152000 426164 152028
rect 407632 151988 407638 152000
rect 426158 151988 426164 152000
rect 426216 151988 426222 152040
rect 434686 152028 434714 152068
rect 442166 152056 442172 152068
rect 442224 152056 442230 152108
rect 442994 152056 443000 152108
rect 443052 152096 443058 152108
rect 458174 152096 458180 152108
rect 443052 152068 458180 152096
rect 443052 152056 443058 152068
rect 458174 152056 458180 152068
rect 458232 152056 458238 152108
rect 485866 152056 485872 152108
rect 485924 152096 485930 152108
rect 490926 152096 490932 152108
rect 485924 152068 490932 152096
rect 485924 152056 485930 152068
rect 490926 152056 490932 152068
rect 490984 152056 490990 152108
rect 426912 152000 434714 152028
rect 386046 151920 386052 151972
rect 386104 151960 386110 151972
rect 399754 151960 399760 151972
rect 386104 151932 399760 151960
rect 386104 151920 386110 151932
rect 399754 151920 399760 151932
rect 399812 151920 399818 151972
rect 404630 151920 404636 151972
rect 404688 151960 404694 151972
rect 423582 151960 423588 151972
rect 404688 151932 423588 151960
rect 404688 151920 404694 151932
rect 423582 151920 423588 151932
rect 423640 151920 423646 151972
rect 424962 151920 424968 151972
rect 425020 151960 425026 151972
rect 426912 151960 426940 152000
rect 436186 151988 436192 152040
rect 436244 152028 436250 152040
rect 446950 152028 446956 152040
rect 436244 152000 446956 152028
rect 436244 151988 436250 152000
rect 446950 151988 446956 152000
rect 447008 151988 447014 152040
rect 447042 151988 447048 152040
rect 447100 152028 447106 152040
rect 453758 152028 453764 152040
rect 447100 152000 453764 152028
rect 447100 151988 447106 152000
rect 453758 151988 453764 152000
rect 453816 151988 453822 152040
rect 456794 151988 456800 152040
rect 456852 152028 456858 152040
rect 463326 152028 463332 152040
rect 456852 152000 463332 152028
rect 456852 151988 456858 152000
rect 463326 151988 463332 152000
rect 463384 151988 463390 152040
rect 467926 151988 467932 152040
rect 467984 152028 467990 152040
rect 472342 152028 472348 152040
rect 467984 152000 472348 152028
rect 467984 151988 467990 152000
rect 472342 151988 472348 152000
rect 472400 151988 472406 152040
rect 487522 151988 487528 152040
rect 487580 152028 487586 152040
rect 492214 152028 492220 152040
rect 487580 152000 492220 152028
rect 487580 151988 487586 152000
rect 492214 151988 492220 152000
rect 492272 151988 492278 152040
rect 499206 151988 499212 152040
rect 499264 152028 499270 152040
rect 500586 152028 500592 152040
rect 499264 152000 500592 152028
rect 499264 151988 499270 152000
rect 500586 151988 500592 152000
rect 500644 151988 500650 152040
rect 439590 151960 439596 151972
rect 425020 151932 426940 151960
rect 427004 151932 439596 151960
rect 425020 151920 425026 151932
rect 378284 151864 383654 151892
rect 378284 151852 378290 151864
rect 385862 151852 385868 151904
rect 385920 151892 385926 151904
rect 397178 151892 397184 151904
rect 385920 151864 397184 151892
rect 385920 151852 385926 151864
rect 397178 151852 397184 151864
rect 397236 151852 397242 151904
rect 397914 151852 397920 151904
rect 397972 151892 397978 151904
rect 405550 151892 405556 151904
rect 397972 151864 405556 151892
rect 397972 151852 397978 151864
rect 405550 151852 405556 151864
rect 405608 151852 405614 151904
rect 405642 151852 405648 151904
rect 405700 151892 405706 151904
rect 421006 151892 421012 151904
rect 405700 151864 421012 151892
rect 405700 151852 405706 151864
rect 421006 151852 421012 151864
rect 421064 151852 421070 151904
rect 422266 151864 422892 151892
rect 328420 151796 331260 151824
rect 328420 151784 328426 151796
rect 334066 151784 334072 151836
rect 334124 151824 334130 151836
rect 372154 151824 372160 151836
rect 334124 151796 372160 151824
rect 334124 151784 334130 151796
rect 372154 151784 372160 151796
rect 372212 151784 372218 151836
rect 380986 151784 380992 151836
rect 381044 151824 381050 151836
rect 392118 151824 392124 151836
rect 381044 151796 392124 151824
rect 381044 151784 381050 151796
rect 392118 151784 392124 151796
rect 392176 151784 392182 151836
rect 397362 151784 397368 151836
rect 397420 151824 397426 151836
rect 402974 151824 402980 151836
rect 397420 151796 402980 151824
rect 397420 151784 397426 151796
rect 402974 151784 402980 151796
rect 403032 151784 403038 151836
rect 419534 151784 419540 151836
rect 419592 151824 419598 151836
rect 422266 151824 422294 151864
rect 419592 151796 422294 151824
rect 419592 151784 419598 151796
rect 81710 151716 81716 151768
rect 81768 151756 81774 151768
rect 112806 151756 112812 151768
rect 81768 151728 112812 151756
rect 81768 151716 81774 151728
rect 112806 151716 112812 151728
rect 112864 151716 112870 151768
rect 422864 151756 422892 151864
rect 423490 151852 423496 151904
rect 423548 151892 423554 151904
rect 427004 151892 427032 151932
rect 439590 151920 439596 151932
rect 439648 151920 439654 151972
rect 441706 151920 441712 151972
rect 441764 151960 441770 151972
rect 446582 151960 446588 151972
rect 441764 151932 446588 151960
rect 441764 151920 441770 151932
rect 446582 151920 446588 151932
rect 446640 151920 446646 151972
rect 446692 151932 446996 151960
rect 423548 151864 427032 151892
rect 423548 151852 423554 151864
rect 427078 151852 427084 151904
rect 427136 151892 427142 151904
rect 437014 151892 437020 151904
rect 427136 151864 437020 151892
rect 427136 151852 427142 151864
rect 437014 151852 437020 151864
rect 437072 151852 437078 151904
rect 437474 151852 437480 151904
rect 437532 151892 437538 151904
rect 445662 151892 445668 151904
rect 437532 151864 445668 151892
rect 437532 151852 437538 151864
rect 445662 151852 445668 151864
rect 445720 151852 445726 151904
rect 445754 151852 445760 151904
rect 445812 151892 445818 151904
rect 446692 151892 446720 151932
rect 445812 151864 446720 151892
rect 446968 151892 446996 151932
rect 448054 151920 448060 151972
rect 448112 151960 448118 151972
rect 456978 151960 456984 151972
rect 448112 151932 456984 151960
rect 448112 151920 448118 151932
rect 456978 151920 456984 151932
rect 457036 151920 457042 151972
rect 468018 151920 468024 151972
rect 468076 151960 468082 151972
rect 471698 151960 471704 151972
rect 468076 151932 471704 151960
rect 468076 151920 468082 151932
rect 471698 151920 471704 151932
rect 471756 151920 471762 151972
rect 487154 151920 487160 151972
rect 487212 151960 487218 151972
rect 491570 151960 491576 151972
rect 487212 151932 491576 151960
rect 487212 151920 487218 151932
rect 491570 151920 491576 151932
rect 491628 151920 491634 151972
rect 498378 151920 498384 151972
rect 498436 151960 498442 151972
rect 499942 151960 499948 151972
rect 498436 151932 499948 151960
rect 498436 151920 498442 151932
rect 499942 151920 499948 151932
rect 500000 151920 500006 151972
rect 516042 151920 516048 151972
rect 516100 151960 516106 151972
rect 518986 151960 518992 151972
rect 516100 151932 518992 151960
rect 516100 151920 516106 151932
rect 518986 151920 518992 151932
rect 519044 151920 519050 151972
rect 460106 151892 460112 151904
rect 446968 151864 460112 151892
rect 445812 151852 445818 151864
rect 460106 151852 460112 151864
rect 460164 151852 460170 151904
rect 460198 151852 460204 151904
rect 460256 151892 460262 151904
rect 462038 151892 462044 151904
rect 460256 151864 462044 151892
rect 460256 151852 460262 151864
rect 462038 151852 462044 151864
rect 462096 151852 462102 151904
rect 469214 151852 469220 151904
rect 469272 151892 469278 151904
rect 472986 151892 472992 151904
rect 469272 151864 472992 151892
rect 469272 151852 469278 151864
rect 472986 151852 472992 151864
rect 473044 151852 473050 151904
rect 478874 151852 478880 151904
rect 478932 151892 478938 151904
rect 480714 151892 480720 151904
rect 478932 151864 480720 151892
rect 478932 151852 478938 151864
rect 480714 151852 480720 151864
rect 480772 151852 480778 151904
rect 517422 151852 517428 151904
rect 517480 151892 517486 151904
rect 520274 151892 520280 151904
rect 517480 151864 520280 151892
rect 517480 151852 517486 151864
rect 520274 151852 520280 151864
rect 520332 151852 520338 151904
rect 434438 151824 434444 151836
rect 423784 151796 434444 151824
rect 423784 151756 423812 151796
rect 434438 151784 434444 151796
rect 434496 151784 434502 151836
rect 441062 151784 441068 151836
rect 441120 151824 441126 151836
rect 446582 151824 446588 151836
rect 441120 151796 446588 151824
rect 441120 151784 441126 151796
rect 446582 151784 446588 151796
rect 446640 151784 446646 151836
rect 446950 151784 446956 151836
rect 447008 151824 447014 151836
rect 455046 151824 455052 151836
rect 447008 151796 455052 151824
rect 447008 151784 447014 151796
rect 455046 151784 455052 151796
rect 455104 151784 455110 151836
rect 466454 151784 466460 151836
rect 466512 151824 466518 151836
rect 471054 151824 471060 151836
rect 466512 151796 471060 151824
rect 466512 151784 466518 151796
rect 471054 151784 471060 151796
rect 471112 151784 471118 151836
rect 485774 151784 485780 151836
rect 485832 151824 485838 151836
rect 490282 151824 490288 151836
rect 485832 151796 490288 151824
rect 485832 151784 485838 151796
rect 490282 151784 490288 151796
rect 490340 151784 490346 151836
rect 422864 151728 423812 151756
rect 98914 151648 98920 151700
rect 98972 151688 98978 151700
rect 116026 151688 116032 151700
rect 98972 151660 116032 151688
rect 98972 151648 98978 151660
rect 116026 151648 116032 151660
rect 116084 151648 116090 151700
rect 95510 151580 95516 151632
rect 95568 151620 95574 151632
rect 115290 151620 115296 151632
rect 95568 151592 115296 151620
rect 95568 151580 95574 151592
rect 115290 151580 115296 151592
rect 115348 151580 115354 151632
rect 92014 151512 92020 151564
rect 92072 151552 92078 151564
rect 113082 151552 113088 151564
rect 92072 151524 113088 151552
rect 92072 151512 92078 151524
rect 113082 151512 113088 151524
rect 113140 151512 113146 151564
rect 26694 151444 26700 151496
rect 26752 151484 26758 151496
rect 116946 151484 116952 151496
rect 26752 151456 116952 151484
rect 26752 151444 26758 151456
rect 116946 151444 116952 151456
rect 117004 151444 117010 151496
rect 16390 151376 16396 151428
rect 16448 151416 16454 151428
rect 116762 151416 116768 151428
rect 16448 151388 116768 151416
rect 16448 151376 16454 151388
rect 116762 151376 116768 151388
rect 116820 151376 116826 151428
rect 12986 151308 12992 151360
rect 13044 151348 13050 151360
rect 116670 151348 116676 151360
rect 13044 151320 116676 151348
rect 13044 151308 13050 151320
rect 116670 151308 116676 151320
rect 116728 151308 116734 151360
rect 68002 151240 68008 151292
rect 68060 151280 68066 151292
rect 112714 151280 112720 151292
rect 68060 151252 112720 151280
rect 68060 151240 68066 151252
rect 112714 151240 112720 151252
rect 112772 151240 112778 151292
rect 64506 151172 64512 151224
rect 64564 151212 64570 151224
rect 112622 151212 112628 151224
rect 64564 151184 112628 151212
rect 64564 151172 64570 151184
rect 112622 151172 112628 151184
rect 112680 151172 112686 151224
rect 61102 151104 61108 151156
rect 61160 151144 61166 151156
rect 112530 151144 112536 151156
rect 61160 151116 112536 151144
rect 61160 151104 61166 151116
rect 112530 151104 112536 151116
rect 112588 151104 112594 151156
rect 57698 151036 57704 151088
rect 57756 151076 57762 151088
rect 110966 151076 110972 151088
rect 57756 151048 110972 151076
rect 57756 151036 57762 151048
rect 110966 151036 110972 151048
rect 111024 151036 111030 151088
rect 54202 150968 54208 151020
rect 54260 151008 54266 151020
rect 112438 151008 112444 151020
rect 54260 150980 112444 151008
rect 54260 150968 54266 150980
rect 112438 150968 112444 150980
rect 112496 150968 112502 151020
rect 50798 150900 50804 150952
rect 50856 150940 50862 150952
rect 111702 150940 111708 150952
rect 50856 150912 111708 150940
rect 50856 150900 50862 150912
rect 111702 150900 111708 150912
rect 111760 150900 111766 150952
rect 47302 150832 47308 150884
rect 47360 150872 47366 150884
rect 111610 150872 111616 150884
rect 47360 150844 111616 150872
rect 47360 150832 47366 150844
rect 111610 150832 111616 150844
rect 111668 150832 111674 150884
rect 43898 150764 43904 150816
rect 43956 150804 43962 150816
rect 111518 150804 111524 150816
rect 43956 150776 111524 150804
rect 43956 150764 43962 150776
rect 111518 150764 111524 150776
rect 111576 150764 111582 150816
rect 40494 150696 40500 150748
rect 40552 150736 40558 150748
rect 111426 150736 111432 150748
rect 40552 150708 111432 150736
rect 40552 150696 40558 150708
rect 111426 150696 111432 150708
rect 111484 150696 111490 150748
rect 36998 150628 37004 150680
rect 37056 150668 37062 150680
rect 111242 150668 111248 150680
rect 37056 150640 111248 150668
rect 37056 150628 37062 150640
rect 111242 150628 111248 150640
rect 111300 150628 111306 150680
rect 88610 150560 88616 150612
rect 88668 150600 88674 150612
rect 112990 150600 112996 150612
rect 88668 150572 112996 150600
rect 88668 150560 88674 150572
rect 112990 150560 112996 150572
rect 113048 150560 113054 150612
rect 85206 150492 85212 150544
rect 85264 150532 85270 150544
rect 115198 150532 115204 150544
rect 85264 150504 115204 150532
rect 85264 150492 85270 150504
rect 115198 150492 115204 150504
rect 115256 150492 115262 150544
rect 102318 150424 102324 150476
rect 102376 150464 102382 150476
rect 116118 150464 116124 150476
rect 102376 150436 116124 150464
rect 102376 150424 102382 150436
rect 116118 150424 116124 150436
rect 116176 150424 116182 150476
rect 78306 150288 78312 150340
rect 78364 150328 78370 150340
rect 112898 150328 112904 150340
rect 78364 150300 112904 150328
rect 78364 150288 78370 150300
rect 112898 150288 112904 150300
rect 112956 150288 112962 150340
rect 109586 150220 109592 150272
rect 109644 150260 109650 150272
rect 117222 150260 117228 150272
rect 109644 150232 117228 150260
rect 109644 150220 109650 150232
rect 117222 150220 117228 150232
rect 117280 150220 117286 150272
rect 108022 150152 108028 150204
rect 108080 150192 108086 150204
rect 117038 150192 117044 150204
rect 108080 150164 117044 150192
rect 108080 150152 108086 150164
rect 117038 150152 117044 150164
rect 117096 150152 117102 150204
rect 145098 150152 145104 150204
rect 145156 150192 145162 150204
rect 146248 150192 146254 150204
rect 145156 150164 146254 150192
rect 145156 150152 145162 150164
rect 146248 150152 146254 150164
rect 146306 150152 146312 150204
rect 146386 150152 146392 150204
rect 146444 150192 146450 150204
rect 147536 150192 147542 150204
rect 146444 150164 147542 150192
rect 146444 150152 146450 150164
rect 147536 150152 147542 150164
rect 147594 150152 147600 150204
rect 163314 150152 163320 150204
rect 163372 150192 163378 150204
rect 164188 150192 164194 150204
rect 163372 150164 164194 150192
rect 163372 150152 163378 150164
rect 164188 150152 164194 150164
rect 164246 150152 164252 150204
rect 164326 150152 164332 150204
rect 164384 150192 164390 150204
rect 165476 150192 165482 150204
rect 164384 150164 165482 150192
rect 164384 150152 164390 150164
rect 165476 150152 165482 150164
rect 165534 150152 165540 150204
rect 171134 150152 171140 150204
rect 171192 150192 171198 150204
rect 171916 150192 171922 150204
rect 171192 150164 171922 150192
rect 171192 150152 171198 150164
rect 171916 150152 171922 150164
rect 171974 150152 171980 150204
rect 181254 150152 181260 150204
rect 181312 150192 181318 150204
rect 182128 150192 182134 150204
rect 181312 150164 182134 150192
rect 181312 150152 181318 150164
rect 182128 150152 182134 150164
rect 182186 150152 182192 150204
rect 182358 150152 182364 150204
rect 182416 150192 182422 150204
rect 183416 150192 183422 150204
rect 182416 150164 183422 150192
rect 182416 150152 182422 150164
rect 183416 150152 183422 150164
rect 183474 150152 183480 150204
rect 183554 150152 183560 150204
rect 183612 150192 183618 150204
rect 184704 150192 184710 150204
rect 183612 150164 184710 150192
rect 183612 150152 183618 150164
rect 184704 150152 184710 150164
rect 184762 150152 184768 150204
rect 200206 150152 200212 150204
rect 200264 150192 200270 150204
rect 201448 150192 201454 150204
rect 200264 150164 201454 150192
rect 200264 150152 200270 150164
rect 201448 150152 201454 150164
rect 201506 150152 201512 150204
rect 213914 150152 213920 150204
rect 213972 150192 213978 150204
rect 214880 150192 214886 150204
rect 213972 150164 214886 150192
rect 213972 150152 213978 150164
rect 214880 150152 214886 150164
rect 214938 150152 214944 150204
rect 218238 150152 218244 150204
rect 218296 150192 218302 150204
rect 219388 150192 219394 150204
rect 218296 150164 219394 150192
rect 218296 150152 218302 150164
rect 219388 150152 219394 150164
rect 219446 150152 219452 150204
rect 238846 150152 238852 150204
rect 238904 150192 238910 150204
rect 239996 150192 240002 150204
rect 238904 150164 240002 150192
rect 238904 150152 238910 150164
rect 239996 150152 240002 150164
rect 240054 150152 240060 150204
rect 242894 150152 242900 150204
rect 242952 150192 242958 150204
rect 243768 150192 243774 150204
rect 242952 150164 243774 150192
rect 242952 150152 242958 150164
rect 243768 150152 243774 150164
rect 243826 150152 243832 150204
rect 247126 150152 247132 150204
rect 247184 150192 247190 150204
rect 248276 150192 248282 150204
rect 247184 150164 248282 150192
rect 247184 150152 247190 150164
rect 248276 150152 248282 150164
rect 248334 150152 248340 150204
rect 251174 150152 251180 150204
rect 251232 150192 251238 150204
rect 252140 150192 252146 150204
rect 251232 150164 252146 150192
rect 251232 150152 251238 150164
rect 252140 150152 252146 150164
rect 252198 150152 252204 150204
rect 256786 150152 256792 150204
rect 256844 150192 256850 150204
rect 257936 150192 257942 150204
rect 256844 150164 257942 150192
rect 256844 150152 256850 150164
rect 257936 150152 257942 150164
rect 257994 150152 258000 150204
rect 258166 150152 258172 150204
rect 258224 150192 258230 150204
rect 259224 150192 259230 150204
rect 258224 150164 259230 150192
rect 258224 150152 258230 150164
rect 259224 150152 259230 150164
rect 259282 150152 259288 150204
rect 260834 150152 260840 150204
rect 260892 150192 260898 150204
rect 261800 150192 261806 150204
rect 260892 150164 261806 150192
rect 260892 150152 260898 150164
rect 261800 150152 261806 150164
rect 261858 150152 261864 150204
rect 271874 150152 271880 150204
rect 271932 150192 271938 150204
rect 272748 150192 272754 150204
rect 271932 150164 272754 150192
rect 271932 150152 271938 150164
rect 272748 150152 272754 150164
rect 272806 150152 272812 150204
rect 311986 150152 311992 150204
rect 312044 150192 312050 150204
rect 313136 150192 313142 150204
rect 312044 150164 313142 150192
rect 312044 150152 312050 150164
rect 313136 150152 313142 150164
rect 313194 150152 313200 150204
rect 328454 150152 328460 150204
rect 328512 150192 328518 150204
rect 329236 150192 329242 150204
rect 328512 150164 329242 150192
rect 328512 150152 328518 150164
rect 329236 150152 329242 150164
rect 329294 150152 329300 150204
rect 332594 150152 332600 150204
rect 332652 150192 332658 150204
rect 333744 150192 333750 150204
rect 332652 150164 333750 150192
rect 332652 150152 332658 150164
rect 333744 150152 333750 150164
rect 333802 150152 333808 150204
rect 339678 150152 339684 150204
rect 339736 150192 339742 150204
rect 340736 150192 340742 150204
rect 339736 150164 340742 150192
rect 339736 150152 339742 150164
rect 340736 150152 340742 150164
rect 340794 150152 340800 150204
rect 349338 150152 349344 150204
rect 349396 150192 349402 150204
rect 350396 150192 350402 150204
rect 349396 150164 350402 150192
rect 349396 150152 349402 150164
rect 350396 150152 350402 150164
rect 350454 150152 350460 150204
rect 357618 150152 357624 150204
rect 357676 150192 357682 150204
rect 358768 150192 358774 150204
rect 357676 150164 358774 150192
rect 357676 150152 357682 150164
rect 358768 150152 358774 150164
rect 358826 150152 358832 150204
rect 358906 150152 358912 150204
rect 358964 150192 358970 150204
rect 360056 150192 360062 150204
rect 358964 150164 360062 150192
rect 358964 150152 358970 150164
rect 360056 150152 360062 150164
rect 360114 150152 360120 150204
rect 363046 150152 363052 150204
rect 363104 150192 363110 150204
rect 363920 150192 363926 150204
rect 363104 150164 363926 150192
rect 363104 150152 363110 150164
rect 363920 150152 363926 150164
rect 363978 150152 363984 150204
rect 368474 150152 368480 150204
rect 368532 150192 368538 150204
rect 369624 150192 369630 150204
rect 368532 150164 369630 150192
rect 368532 150152 368538 150164
rect 369624 150152 369630 150164
rect 369682 150152 369688 150204
rect 403158 150152 403164 150204
rect 403216 150192 403222 150204
rect 404308 150192 404314 150204
rect 403216 150164 404314 150192
rect 403216 150152 403222 150164
rect 404308 150152 404314 150164
rect 404366 150152 404372 150204
rect 446582 150152 446588 150204
rect 446640 150192 446646 150204
rect 448008 150192 448014 150204
rect 446640 150164 448014 150192
rect 446640 150152 446646 150164
rect 448008 150152 448014 150164
rect 448066 150152 448072 150204
rect 465074 150152 465080 150204
rect 465132 150192 465138 150204
rect 465948 150192 465954 150204
rect 465132 150164 465954 150192
rect 465132 150152 465138 150164
rect 465948 150152 465954 150164
rect 466006 150152 466012 150204
rect 477678 150152 477684 150204
rect 477736 150192 477742 150204
rect 478828 150192 478834 150204
rect 477736 150164 478834 150192
rect 477736 150152 477742 150164
rect 478828 150152 478834 150164
rect 478886 150152 478892 150204
rect 483106 150152 483112 150204
rect 483164 150192 483170 150204
rect 483980 150192 483986 150204
rect 483164 150164 483986 150192
rect 483164 150152 483170 150164
rect 483980 150152 483986 150164
rect 484038 150152 484044 150204
rect 505278 150152 505284 150204
rect 505336 150192 505342 150204
rect 506428 150192 506434 150204
rect 505336 150164 506434 150192
rect 505336 150152 505342 150164
rect 506428 150152 506434 150164
rect 506486 150152 506492 150204
rect 506566 150152 506572 150204
rect 506624 150192 506630 150204
rect 507716 150192 507722 150204
rect 506624 150164 507722 150192
rect 506624 150152 506630 150164
rect 507716 150152 507722 150164
rect 507774 150152 507780 150204
rect 507946 150152 507952 150204
rect 508004 150192 508010 150204
rect 509004 150192 509010 150204
rect 508004 150164 509010 150192
rect 508004 150152 508010 150164
rect 509004 150152 509010 150164
rect 509062 150152 509068 150204
rect 509326 150152 509332 150204
rect 509384 150192 509390 150204
rect 510292 150192 510298 150204
rect 509384 150164 510298 150192
rect 509384 150152 509390 150164
rect 510292 150152 510298 150164
rect 510350 150152 510356 150204
rect 518020 150152 518026 150204
rect 518078 150192 518084 150204
rect 518802 150192 518808 150204
rect 518078 150164 518808 150192
rect 518078 150152 518084 150164
rect 518802 150152 518808 150164
rect 518860 150152 518866 150204
rect 82078 150084 82084 150136
rect 82136 150124 82142 150136
rect 82136 150096 84194 150124
rect 82136 150084 82142 150096
rect 84166 150056 84194 150096
rect 91002 150084 91008 150136
rect 91060 150124 91066 150136
rect 116486 150124 116492 150136
rect 91060 150096 116492 150124
rect 91060 150084 91066 150096
rect 116486 150084 116492 150096
rect 116544 150084 116550 150136
rect 146570 150084 146576 150136
rect 146628 150124 146634 150136
rect 150664 150124 150670 150136
rect 146628 150096 150670 150124
rect 146628 150084 146634 150096
rect 150664 150084 150670 150096
rect 150722 150084 150728 150136
rect 116394 150056 116400 150068
rect 84166 150028 116400 150056
rect 116394 150016 116400 150028
rect 116452 150016 116458 150068
rect 111150 148316 111156 148368
rect 111208 148356 111214 148368
rect 117130 148356 117136 148368
rect 111208 148328 117136 148356
rect 111208 148316 111214 148328
rect 117130 148316 117136 148328
rect 117188 148316 117194 148368
rect 113082 140700 113088 140752
rect 113140 140740 113146 140752
rect 116118 140740 116124 140752
rect 113140 140712 116124 140740
rect 113140 140700 113146 140712
rect 116118 140700 116124 140712
rect 116176 140700 116182 140752
rect 112990 137912 112996 137964
rect 113048 137952 113054 137964
rect 116118 137952 116124 137964
rect 113048 137924 116124 137952
rect 113048 137912 113054 137924
rect 116118 137912 116124 137924
rect 116176 137912 116182 137964
rect 116302 137300 116308 137352
rect 116360 137340 116366 137352
rect 116486 137340 116492 137352
rect 116360 137312 116492 137340
rect 116360 137300 116366 137312
rect 116486 137300 116492 137312
rect 116544 137300 116550 137352
rect 112806 133832 112812 133884
rect 112864 133872 112870 133884
rect 116026 133872 116032 133884
rect 112864 133844 116032 133872
rect 112864 133832 112870 133844
rect 116026 133832 116032 133844
rect 116084 133832 116090 133884
rect 114186 132608 114192 132660
rect 114244 132648 114250 132660
rect 115198 132648 115204 132660
rect 114244 132620 115204 132648
rect 114244 132608 114250 132620
rect 115198 132608 115204 132620
rect 115256 132608 115262 132660
rect 112898 132404 112904 132456
rect 112956 132444 112962 132456
rect 116118 132444 116124 132456
rect 112956 132416 116124 132444
rect 112956 132404 112962 132416
rect 116118 132404 116124 132416
rect 116176 132404 116182 132456
rect 112714 126896 112720 126948
rect 112772 126936 112778 126948
rect 116026 126936 116032 126948
rect 112772 126908 116032 126936
rect 112772 126896 112778 126908
rect 116026 126896 116032 126908
rect 116084 126896 116090 126948
rect 112622 124108 112628 124160
rect 112680 124148 112686 124160
rect 116118 124148 116124 124160
rect 112680 124120 116124 124148
rect 112680 124108 112686 124120
rect 116118 124108 116124 124120
rect 116176 124108 116182 124160
rect 112530 122748 112536 122800
rect 112588 122788 112594 122800
rect 115934 122788 115940 122800
rect 112588 122760 115940 122788
rect 112588 122748 112594 122760
rect 115934 122748 115940 122760
rect 115992 122748 115998 122800
rect 111702 121388 111708 121440
rect 111760 121428 111766 121440
rect 116118 121428 116124 121440
rect 111760 121400 116124 121428
rect 111760 121388 111766 121400
rect 116118 121388 116124 121400
rect 116176 121388 116182 121440
rect 112438 118600 112444 118652
rect 112496 118640 112502 118652
rect 116118 118640 116124 118652
rect 112496 118612 116124 118640
rect 112496 118600 112502 118612
rect 116118 118600 116124 118612
rect 116176 118600 116182 118652
rect 116486 117988 116492 118040
rect 116544 118028 116550 118040
rect 117222 118028 117228 118040
rect 116544 118000 117228 118028
rect 116544 117988 116550 118000
rect 117222 117988 117228 118000
rect 117280 117988 117286 118040
rect 111610 117240 111616 117292
rect 111668 117280 111674 117292
rect 116118 117280 116124 117292
rect 111668 117252 116124 117280
rect 111668 117240 111674 117252
rect 116118 117240 116124 117252
rect 116176 117240 116182 117292
rect 111518 114452 111524 114504
rect 111576 114492 111582 114504
rect 116118 114492 116124 114504
rect 111576 114464 116124 114492
rect 111576 114452 111582 114464
rect 116118 114452 116124 114464
rect 116176 114452 116182 114504
rect 111426 113092 111432 113144
rect 111484 113132 111490 113144
rect 115934 113132 115940 113144
rect 111484 113104 115940 113132
rect 111484 113092 111490 113104
rect 115934 113092 115940 113104
rect 115992 113092 115998 113144
rect 111334 111732 111340 111784
rect 111392 111772 111398 111784
rect 116118 111772 116124 111784
rect 111392 111744 116124 111772
rect 111392 111732 111398 111744
rect 116118 111732 116124 111744
rect 116176 111732 116182 111784
rect 111150 108944 111156 108996
rect 111208 108984 111214 108996
rect 116118 108984 116124 108996
rect 111208 108956 116124 108984
rect 111208 108944 111214 108956
rect 116118 108944 116124 108956
rect 116176 108944 116182 108996
rect 111242 92420 111248 92472
rect 111300 92460 111306 92472
rect 116118 92460 116124 92472
rect 111300 92432 116124 92460
rect 111300 92420 111306 92432
rect 116118 92420 116124 92432
rect 116176 92420 116182 92472
rect 111058 89632 111064 89684
rect 111116 89672 111122 89684
rect 116118 89672 116124 89684
rect 111116 89644 116124 89672
rect 111116 89632 111122 89644
rect 116118 89632 116124 89644
rect 116176 89632 116182 89684
rect 113818 88272 113824 88324
rect 113876 88312 113882 88324
rect 116026 88312 116032 88324
rect 113876 88284 116032 88312
rect 113876 88272 113882 88284
rect 116026 88272 116032 88284
rect 116084 88272 116090 88324
rect 113910 83920 113916 83972
rect 113968 83960 113974 83972
rect 116578 83960 116584 83972
rect 113968 83932 116584 83960
rect 113968 83920 113974 83932
rect 116578 83920 116584 83932
rect 116636 83920 116642 83972
rect 114002 82764 114008 82816
rect 114060 82804 114066 82816
rect 116210 82804 116216 82816
rect 114060 82776 116216 82804
rect 114060 82764 114066 82776
rect 116210 82764 116216 82776
rect 116268 82764 116274 82816
rect 114094 79976 114100 80028
rect 114152 80016 114158 80028
rect 115934 80016 115940 80028
rect 114152 79988 115940 80016
rect 114152 79976 114158 79988
rect 115934 79976 115940 79988
rect 115992 79976 115998 80028
rect 114186 78616 114192 78668
rect 114244 78656 114250 78668
rect 116118 78656 116124 78668
rect 114244 78628 116124 78656
rect 114244 78616 114250 78628
rect 116118 78616 116124 78628
rect 116176 78616 116182 78668
rect 114186 71748 114192 71800
rect 114244 71788 114250 71800
rect 116578 71788 116584 71800
rect 114244 71760 116584 71788
rect 114244 71748 114250 71760
rect 116578 71748 116584 71760
rect 116636 71748 116642 71800
rect 114094 69028 114100 69080
rect 114152 69068 114158 69080
rect 116302 69068 116308 69080
rect 114152 69040 116308 69068
rect 114152 69028 114158 69040
rect 116302 69028 116308 69040
rect 116360 69028 116366 69080
rect 114002 67600 114008 67652
rect 114060 67640 114066 67652
rect 116118 67640 116124 67652
rect 114060 67612 116124 67640
rect 114060 67600 114066 67612
rect 116118 67600 116124 67612
rect 116176 67600 116182 67652
rect 113910 66240 113916 66292
rect 113968 66280 113974 66292
rect 116578 66280 116584 66292
rect 113968 66252 116584 66280
rect 113968 66240 113974 66252
rect 116578 66240 116584 66252
rect 116636 66240 116642 66292
rect 113358 64676 113364 64728
rect 113416 64716 113422 64728
rect 116578 64716 116584 64728
rect 113416 64688 116584 64716
rect 113416 64676 113422 64688
rect 116578 64676 116584 64688
rect 116636 64676 116642 64728
rect 113818 63520 113824 63572
rect 113876 63560 113882 63572
rect 116210 63560 116216 63572
rect 113876 63532 116216 63560
rect 113876 63520 113882 63532
rect 116210 63520 116216 63532
rect 116268 63520 116274 63572
rect 112438 62092 112444 62144
rect 112496 62132 112502 62144
rect 116118 62132 116124 62144
rect 112496 62104 116124 62132
rect 112496 62092 112502 62104
rect 116118 62092 116124 62104
rect 116176 62092 116182 62144
rect 112530 42780 112536 42832
rect 112588 42820 112594 42832
rect 116118 42820 116124 42832
rect 112588 42792 116124 42820
rect 112588 42780 112594 42792
rect 116118 42780 116124 42792
rect 116176 42780 116182 42832
rect 115842 7896 115848 7948
rect 115900 7936 115906 7948
rect 116762 7936 116768 7948
rect 115900 7908 116768 7936
rect 115900 7896 115906 7908
rect 116762 7896 116768 7908
rect 116820 7896 116826 7948
rect 117222 7868 117228 7880
rect 116688 7840 117228 7868
rect 116688 7744 116716 7840
rect 117222 7828 117228 7840
rect 117280 7828 117286 7880
rect 116946 7760 116952 7812
rect 117004 7760 117010 7812
rect 117038 7760 117044 7812
rect 117096 7800 117102 7812
rect 117314 7800 117320 7812
rect 117096 7772 117320 7800
rect 117096 7760 117102 7772
rect 117314 7760 117320 7772
rect 117372 7760 117378 7812
rect 116670 7692 116676 7744
rect 116728 7692 116734 7744
rect 116964 7460 116992 7760
rect 117038 7460 117044 7472
rect 116964 7432 117044 7460
rect 117038 7420 117044 7432
rect 117096 7420 117102 7472
rect 170140 3012 179414 3040
rect 111702 2864 111708 2916
rect 111760 2904 111766 2916
rect 111760 2876 170076 2904
rect 111760 2864 111766 2876
rect 111794 2796 111800 2848
rect 111852 2836 111858 2848
rect 111852 2808 168374 2836
rect 111852 2796 111858 2808
rect 168346 2360 168374 2808
rect 170048 2774 170076 2876
rect 169956 2746 170076 2774
rect 169956 2700 169984 2746
rect 169680 2672 169984 2700
rect 170140 2700 170168 3012
rect 179386 2972 179414 3012
rect 180766 3012 183554 3040
rect 180766 2972 180794 3012
rect 179386 2944 180794 2972
rect 183526 2972 183554 3012
rect 183526 2944 200114 2972
rect 183526 2876 186452 2904
rect 183526 2768 183554 2876
rect 186424 2836 186452 2876
rect 200086 2836 200114 2944
rect 186424 2808 193444 2836
rect 200086 2808 293954 2836
rect 182146 2740 183554 2768
rect 182146 2700 182174 2740
rect 170140 2672 170352 2700
rect 169680 2428 169708 2672
rect 170324 2508 170352 2672
rect 178006 2672 182174 2700
rect 178006 2632 178034 2672
rect 176626 2604 178034 2632
rect 170306 2456 170312 2508
rect 170364 2456 170370 2508
rect 176626 2428 176654 2604
rect 193416 2496 193444 2808
rect 193582 2496 193588 2508
rect 193416 2468 193588 2496
rect 193582 2456 193588 2468
rect 193640 2456 193646 2508
rect 293926 2496 293954 2808
rect 425808 2808 443684 2836
rect 425808 2508 425836 2808
rect 443656 2508 443684 2808
rect 294782 2496 294788 2508
rect 293926 2468 294788 2496
rect 294782 2456 294788 2468
rect 294840 2456 294846 2508
rect 425790 2456 425796 2508
rect 425848 2456 425854 2508
rect 443638 2456 443644 2508
rect 443696 2456 443702 2508
rect 169680 2400 176654 2428
rect 170306 2360 170312 2372
rect 168346 2332 170312 2360
rect 170306 2320 170312 2332
rect 170364 2320 170370 2372
rect 111058 1952 111064 1964
rect 93826 1924 100984 1952
rect 62390 1844 62396 1896
rect 62448 1884 62454 1896
rect 65334 1884 65340 1896
rect 62448 1856 65340 1884
rect 62448 1844 62454 1856
rect 65334 1844 65340 1856
rect 65392 1844 65398 1896
rect 68002 1844 68008 1896
rect 68060 1884 68066 1896
rect 77110 1884 77116 1896
rect 68060 1856 77116 1884
rect 68060 1844 68066 1856
rect 77110 1844 77116 1856
rect 77168 1844 77174 1896
rect 77754 1844 77760 1896
rect 77812 1884 77818 1896
rect 88334 1884 88340 1896
rect 77812 1856 88340 1884
rect 77812 1844 77818 1856
rect 88334 1844 88340 1856
rect 88392 1844 88398 1896
rect 89346 1844 89352 1896
rect 89404 1884 89410 1896
rect 93826 1884 93854 1924
rect 89404 1856 93854 1884
rect 89404 1844 89410 1856
rect 94866 1844 94872 1896
rect 94924 1884 94930 1896
rect 100754 1884 100760 1896
rect 94924 1856 100760 1884
rect 94924 1844 94930 1856
rect 100754 1844 100760 1856
rect 100812 1844 100818 1896
rect 64138 1776 64144 1828
rect 64196 1816 64202 1828
rect 69382 1816 69388 1828
rect 64196 1788 69388 1816
rect 64196 1776 64202 1788
rect 69382 1776 69388 1788
rect 69440 1776 69446 1828
rect 77018 1776 77024 1828
rect 77076 1816 77082 1828
rect 85942 1816 85948 1828
rect 77076 1788 85948 1816
rect 77076 1776 77082 1788
rect 85942 1776 85948 1788
rect 86000 1776 86006 1828
rect 86034 1776 86040 1828
rect 86092 1816 86098 1828
rect 100956 1816 100984 1924
rect 102704 1924 111064 1952
rect 102704 1896 102732 1924
rect 111058 1912 111064 1924
rect 111116 1912 111122 1964
rect 102686 1844 102692 1896
rect 102744 1844 102750 1896
rect 104158 1844 104164 1896
rect 104216 1884 104222 1896
rect 109218 1884 109224 1896
rect 104216 1856 109224 1884
rect 104216 1844 104222 1856
rect 109218 1844 109224 1856
rect 109276 1844 109282 1896
rect 109310 1844 109316 1896
rect 109368 1884 109374 1896
rect 109368 1856 110184 1884
rect 109368 1844 109374 1856
rect 109586 1816 109592 1828
rect 86092 1788 100892 1816
rect 100956 1788 109592 1816
rect 86092 1776 86098 1788
rect 62666 1708 62672 1760
rect 62724 1748 62730 1760
rect 68830 1748 68836 1760
rect 62724 1720 68836 1748
rect 62724 1708 62730 1720
rect 68830 1708 68836 1720
rect 68888 1708 68894 1760
rect 77938 1708 77944 1760
rect 77996 1748 78002 1760
rect 78306 1748 78312 1760
rect 77996 1720 78312 1748
rect 77996 1708 78002 1720
rect 78306 1708 78312 1720
rect 78364 1708 78370 1760
rect 82630 1708 82636 1760
rect 82688 1748 82694 1760
rect 100708 1748 100714 1760
rect 82688 1720 100714 1748
rect 82688 1708 82694 1720
rect 100708 1708 100714 1720
rect 100766 1708 100772 1760
rect 100864 1748 100892 1788
rect 109586 1776 109592 1788
rect 109644 1776 109650 1828
rect 109954 1748 109960 1760
rect 100864 1720 109960 1748
rect 109954 1708 109960 1720
rect 110012 1708 110018 1760
rect 110156 1748 110184 1856
rect 112438 1748 112444 1760
rect 110156 1720 112444 1748
rect 112438 1708 112444 1720
rect 112496 1708 112502 1760
rect 69290 1640 69296 1692
rect 69348 1680 69354 1692
rect 101030 1680 101036 1692
rect 69348 1652 101036 1680
rect 69348 1640 69354 1652
rect 101030 1640 101036 1652
rect 101088 1640 101094 1692
rect 104158 1680 104164 1692
rect 101140 1652 104164 1680
rect 59354 1572 59360 1624
rect 59412 1612 59418 1624
rect 68554 1612 68560 1624
rect 59412 1584 68560 1612
rect 59412 1572 59418 1584
rect 68554 1572 68560 1584
rect 68612 1572 68618 1624
rect 79318 1572 79324 1624
rect 79376 1612 79382 1624
rect 97258 1612 97264 1624
rect 79376 1584 97264 1612
rect 79376 1572 79382 1584
rect 97258 1572 97264 1584
rect 97316 1572 97322 1624
rect 99374 1572 99380 1624
rect 99432 1612 99438 1624
rect 100708 1612 100714 1624
rect 99432 1584 100714 1612
rect 99432 1572 99438 1584
rect 100708 1572 100714 1584
rect 100766 1572 100772 1624
rect 100938 1572 100944 1624
rect 100996 1612 101002 1624
rect 101140 1612 101168 1652
rect 104158 1640 104164 1652
rect 104216 1640 104222 1692
rect 105998 1640 106004 1692
rect 106056 1680 106062 1692
rect 116578 1680 116584 1692
rect 106056 1652 116584 1680
rect 106056 1640 106062 1652
rect 116578 1640 116584 1652
rect 116636 1640 116642 1692
rect 100996 1584 101168 1612
rect 100996 1572 101002 1584
rect 101214 1572 101220 1624
rect 101272 1612 101278 1624
rect 110138 1612 110144 1624
rect 101272 1584 110144 1612
rect 101272 1572 101278 1584
rect 110138 1572 110144 1584
rect 110196 1572 110202 1624
rect 72694 1504 72700 1556
rect 72752 1544 72758 1556
rect 110414 1544 110420 1556
rect 72752 1516 110420 1544
rect 72752 1504 72758 1516
rect 110414 1504 110420 1516
rect 110472 1504 110478 1556
rect 42610 1436 42616 1488
rect 42668 1476 42674 1488
rect 78122 1476 78128 1488
rect 42668 1448 78128 1476
rect 42668 1436 42674 1448
rect 78122 1436 78128 1448
rect 78180 1436 78186 1488
rect 97258 1436 97264 1488
rect 97316 1476 97322 1488
rect 104158 1476 104164 1488
rect 97316 1448 104164 1476
rect 97316 1436 97322 1448
rect 104158 1436 104164 1448
rect 104216 1436 104222 1488
rect 104250 1436 104256 1488
rect 104308 1476 104314 1488
rect 106274 1476 106280 1488
rect 104308 1448 106280 1476
rect 104308 1436 104314 1448
rect 106274 1436 106280 1448
rect 106332 1436 106338 1488
rect 106366 1436 106372 1488
rect 106424 1476 106430 1488
rect 109310 1476 109316 1488
rect 106424 1448 109316 1476
rect 106424 1436 106430 1448
rect 109310 1436 109316 1448
rect 109368 1436 109374 1488
rect 109402 1436 109408 1488
rect 109460 1476 109466 1488
rect 143626 1476 143632 1488
rect 109460 1448 143632 1476
rect 109460 1436 109466 1448
rect 143626 1436 143632 1448
rect 143684 1436 143690 1488
rect 46014 1368 46020 1420
rect 46072 1408 46078 1420
rect 116486 1408 116492 1420
rect 46072 1380 116492 1408
rect 46072 1368 46078 1380
rect 116486 1368 116492 1380
rect 116544 1368 116550 1420
rect 294782 1368 294788 1420
rect 294840 1408 294846 1420
rect 343634 1408 343640 1420
rect 294840 1380 343640 1408
rect 294840 1368 294846 1380
rect 343634 1368 343640 1380
rect 343692 1368 343698 1420
rect 491294 1368 491300 1420
rect 491352 1408 491358 1420
rect 493594 1408 493600 1420
rect 491352 1380 493600 1408
rect 491352 1368 491358 1380
rect 493594 1368 493600 1380
rect 493652 1368 493658 1420
rect 2682 1300 2688 1352
rect 2740 1340 2746 1352
rect 116302 1340 116308 1352
rect 2740 1312 116308 1340
rect 2740 1300 2746 1312
rect 116302 1300 116308 1312
rect 116360 1300 116366 1352
rect 39298 1232 39304 1284
rect 39356 1272 39362 1284
rect 116394 1272 116400 1284
rect 39356 1244 116400 1272
rect 39356 1232 39362 1244
rect 116394 1232 116400 1244
rect 116452 1232 116458 1284
rect 49326 1164 49332 1216
rect 49384 1204 49390 1216
rect 116670 1204 116676 1216
rect 49384 1176 116676 1204
rect 49384 1164 49390 1176
rect 116670 1164 116676 1176
rect 116728 1164 116734 1216
rect 52638 1096 52644 1148
rect 52696 1136 52702 1148
rect 117222 1136 117228 1148
rect 52696 1108 117228 1136
rect 52696 1096 52702 1108
rect 117222 1096 117228 1108
rect 117280 1096 117286 1148
rect 55950 1028 55956 1080
rect 56008 1068 56014 1080
rect 111794 1068 111800 1080
rect 56008 1040 111800 1068
rect 56008 1028 56014 1040
rect 111794 1028 111800 1040
rect 111852 1028 111858 1080
rect 65978 960 65984 1012
rect 66036 1000 66042 1012
rect 116854 1000 116860 1012
rect 66036 972 116860 1000
rect 66036 960 66042 972
rect 116854 960 116860 972
rect 116912 960 116918 1012
rect 76006 892 76012 944
rect 76064 932 76070 944
rect 112530 932 112536 944
rect 76064 904 112536 932
rect 76064 892 76070 904
rect 112530 892 112536 904
rect 112588 892 112594 944
rect 98362 824 98368 876
rect 98420 864 98426 876
rect 105078 864 105084 876
rect 98420 836 105084 864
rect 98420 824 98426 836
rect 105078 824 105084 836
rect 105136 824 105142 876
rect 92658 756 92664 808
rect 92716 796 92722 808
rect 110046 796 110052 808
rect 92716 768 110052 796
rect 92716 756 92722 768
rect 110046 756 110052 768
rect 110104 756 110110 808
rect 103698 688 103704 740
rect 103756 728 103762 740
rect 106366 728 106372 740
rect 103756 700 106372 728
rect 103756 688 103762 700
rect 106366 688 106372 700
rect 106424 688 106430 740
<< via1 >>
rect 126336 160080 126388 160132
rect 128360 160080 128412 160132
rect 153016 160080 153068 160132
rect 66720 160012 66772 160064
rect 142804 160012 142856 160064
rect 142896 160012 142948 160064
rect 154488 160012 154540 160064
rect 158812 160012 158864 160064
rect 159916 160012 159968 160064
rect 196164 160012 196216 160064
rect 207756 160012 207808 160064
rect 276112 160012 276164 160064
rect 277492 160012 277544 160064
rect 280160 160012 280212 160064
rect 280804 160012 280856 160064
rect 76748 159944 76800 159996
rect 164516 159944 164568 159996
rect 166632 159944 166684 159996
rect 197636 159944 197688 159996
rect 201040 159944 201092 159996
rect 271880 159944 271932 159996
rect 274916 159944 274968 159996
rect 324412 159944 324464 159996
rect 324504 159944 324556 159996
rect 328368 159944 328420 159996
rect 328460 159944 328512 159996
rect 331312 159944 331364 159996
rect 331496 160012 331548 160064
rect 334072 160012 334124 160064
rect 334624 160012 334676 160064
rect 374736 160012 374788 160064
rect 381636 160012 381688 160064
rect 398840 160012 398892 160064
rect 401784 160012 401836 160064
rect 407580 160012 407632 160064
rect 426992 160012 427044 160064
rect 445300 160012 445352 160064
rect 332600 159944 332652 159996
rect 333704 159944 333756 159996
rect 374000 159944 374052 159996
rect 374920 159944 374972 159996
rect 397920 159944 397972 159996
rect 399208 159944 399260 159996
rect 418252 159944 418304 159996
rect 424416 159944 424468 159996
rect 443460 159944 443512 159996
rect 457996 159944 458048 159996
rect 464896 159944 464948 159996
rect 466460 159944 466512 159996
rect 473360 159944 473412 159996
rect 479064 159944 479116 159996
rect 485228 159944 485280 159996
rect 49884 159876 49936 159928
rect 133604 159876 133656 159928
rect 133696 159876 133748 159928
rect 137100 159876 137152 159928
rect 137284 159876 137336 159928
rect 142712 159876 142764 159928
rect 142804 159876 142856 159928
rect 70032 159808 70084 159860
rect 153016 159808 153068 159860
rect 153200 159876 153252 159928
rect 189724 159876 189776 159928
rect 194324 159876 194376 159928
rect 267556 159876 267608 159928
rect 270776 159876 270828 159928
rect 273352 159876 273404 159928
rect 274088 159876 274140 159928
rect 328552 159876 328604 159928
rect 328736 159876 328788 159928
rect 370044 159876 370096 159928
rect 374092 159876 374144 159928
rect 380716 159876 380768 159928
rect 380808 159876 380860 159928
rect 388628 159876 388680 159928
rect 389180 159876 389232 159928
rect 415952 159876 416004 159928
rect 416044 159876 416096 159928
rect 423404 159876 423456 159928
rect 423588 159876 423640 159928
rect 442816 159876 442868 159928
rect 154396 159808 154448 159860
rect 156512 159808 156564 159860
rect 172428 159808 172480 159860
rect 176660 159808 176712 159860
rect 181996 159808 182048 159860
rect 184296 159808 184348 159860
rect 185032 159808 185084 159860
rect 60004 159740 60056 159792
rect 149060 159740 149112 159792
rect 149796 159740 149848 159792
rect 180800 159740 180852 159792
rect 180892 159740 180944 159792
rect 255504 159808 255556 159860
rect 260656 159808 260708 159860
rect 317144 159808 317196 159860
rect 187608 159740 187660 159792
rect 262220 159740 262272 159792
rect 267372 159740 267424 159792
rect 317788 159740 317840 159792
rect 318892 159740 318944 159792
rect 321100 159808 321152 159860
rect 363236 159808 363288 159860
rect 364800 159808 364852 159860
rect 395528 159808 395580 159860
rect 410156 159808 410208 159860
rect 432512 159808 432564 159860
rect 450452 159808 450504 159860
rect 456800 159808 456852 159860
rect 458916 159808 458968 159860
rect 465356 159808 465408 159860
rect 467288 159808 467340 159860
rect 473452 159808 473504 159860
rect 482376 159808 482428 159860
rect 487344 159808 487396 159860
rect 321560 159740 321612 159792
rect 326988 159740 327040 159792
rect 368940 159740 368992 159792
rect 375748 159740 375800 159792
rect 405832 159740 405884 159792
rect 406844 159740 406896 159792
rect 429936 159740 429988 159792
rect 448796 159740 448848 159792
rect 460204 159740 460256 159792
rect 53288 159672 53340 159724
rect 137284 159672 137336 159724
rect 137376 159672 137428 159724
rect 139308 159672 139360 159724
rect 139768 159672 139820 159724
rect 158720 159672 158772 159724
rect 39856 159604 39908 159656
rect 124036 159604 124088 159656
rect 127164 159604 127216 159656
rect 136272 159604 136324 159656
rect 136364 159604 136416 159656
rect 164148 159672 164200 159724
rect 167460 159672 167512 159724
rect 242992 159672 243044 159724
rect 248052 159672 248104 159724
rect 308496 159672 308548 159724
rect 315304 159672 315356 159724
rect 351276 159672 351328 159724
rect 351368 159672 351420 159724
rect 357808 159672 357860 159724
rect 369032 159672 369084 159724
rect 401048 159672 401100 159724
rect 403440 159672 403492 159724
rect 427360 159672 427412 159724
rect 447140 159672 447192 159724
rect 458180 159672 458232 159724
rect 459744 159672 459796 159724
rect 466552 159672 466604 159724
rect 472348 159672 472400 159724
rect 479432 159672 479484 159724
rect 479892 159672 479944 159724
rect 485964 159672 486016 159724
rect 163228 159604 163280 159656
rect 174084 159604 174136 159656
rect 174176 159604 174228 159656
rect 251180 159604 251232 159656
rect 254768 159604 254820 159656
rect 313740 159604 313792 159656
rect 314384 159604 314436 159656
rect 357532 159604 357584 159656
rect 357624 159604 357676 159656
rect 358820 159604 358872 159656
rect 362316 159604 362368 159656
rect 395252 159604 395304 159656
rect 407672 159604 407724 159656
rect 430672 159604 430724 159656
rect 453856 159604 453908 159656
rect 465080 159604 465132 159656
rect 470600 159604 470652 159656
rect 477684 159604 477736 159656
rect 480720 159604 480772 159656
rect 486516 159604 486568 159656
rect 22192 159536 22244 159588
rect 127256 159536 127308 159588
rect 127624 159536 127676 159588
rect 133696 159536 133748 159588
rect 133788 159536 133840 159588
rect 139492 159536 139544 159588
rect 140596 159536 140648 159588
rect 218152 159536 218204 159588
rect 221188 159536 221240 159588
rect 28908 159468 28960 159520
rect 132868 159468 132920 159520
rect 23020 159400 23072 159452
rect 136548 159468 136600 159520
rect 137192 159468 137244 159520
rect 142804 159468 142856 159520
rect 142988 159468 143040 159520
rect 144460 159468 144512 159520
rect 147312 159468 147364 159520
rect 226340 159468 226392 159520
rect 227904 159468 227956 159520
rect 287336 159468 287388 159520
rect 287520 159536 287572 159588
rect 337016 159536 337068 159588
rect 288072 159468 288124 159520
rect 291660 159468 291712 159520
rect 295064 159468 295116 159520
rect 295156 159468 295208 159520
rect 337936 159468 337988 159520
rect 339500 159468 339552 159520
rect 342168 159536 342220 159588
rect 380532 159536 380584 159588
rect 380716 159536 380768 159588
rect 344560 159468 344612 159520
rect 344652 159468 344704 159520
rect 382556 159468 382608 159520
rect 385776 159536 385828 159588
rect 413192 159536 413244 159588
rect 416872 159536 416924 159588
rect 437664 159536 437716 159588
rect 451280 159536 451332 159588
rect 463700 159536 463752 159588
rect 469772 159536 469824 159588
rect 476120 159536 476172 159588
rect 478144 159536 478196 159588
rect 484584 159536 484636 159588
rect 388720 159468 388772 159520
rect 413560 159468 413612 159520
rect 435088 159468 435140 159520
rect 454684 159468 454736 159520
rect 466644 159468 466696 159520
rect 484032 159468 484084 159520
rect 489000 159468 489052 159520
rect 133052 159400 133104 159452
rect 156604 159400 156656 159452
rect 160744 159400 160796 159452
rect 240324 159400 240376 159452
rect 247224 159400 247276 159452
rect 307760 159400 307812 159452
rect 308588 159400 308640 159452
rect 349804 159400 349856 159452
rect 349896 159400 349948 159452
rect 354220 159400 354272 159452
rect 2872 159332 2924 159384
rect 116124 159332 116176 159384
rect 116216 159332 116268 159384
rect 127624 159332 127676 159384
rect 129648 159332 129700 159384
rect 142896 159332 142948 159384
rect 142988 159332 143040 159384
rect 147128 159332 147180 159384
rect 150624 159332 150676 159384
rect 152740 159332 152792 159384
rect 154028 159332 154080 159384
rect 236736 159332 236788 159384
rect 241336 159332 241388 159384
rect 303436 159332 303488 159384
rect 307668 159332 307720 159384
rect 348792 159332 348844 159384
rect 348884 159332 348936 159384
rect 83464 159264 83516 159316
rect 167000 159264 167052 159316
rect 169944 159264 169996 159316
rect 195336 159264 195388 159316
rect 197728 159264 197780 159316
rect 214380 159264 214432 159316
rect 214472 159264 214524 159316
rect 282828 159264 282880 159316
rect 287336 159264 287388 159316
rect 293224 159264 293276 159316
rect 294236 159264 294288 159316
rect 343640 159264 343692 159316
rect 343824 159264 343876 159316
rect 349988 159264 350040 159316
rect 351276 159332 351328 159384
rect 357624 159400 357676 159452
rect 358084 159400 358136 159452
rect 392400 159400 392452 159452
rect 395068 159400 395120 159452
rect 405648 159400 405700 159452
rect 420276 159400 420328 159452
rect 440332 159400 440384 159452
rect 452108 159400 452160 159452
rect 464252 159400 464304 159452
rect 468944 159400 468996 159452
rect 475016 159400 475068 159452
rect 476488 159400 476540 159452
rect 483296 159400 483348 159452
rect 518808 159400 518860 159452
rect 521844 159400 521896 159452
rect 355600 159332 355652 159384
rect 390744 159332 390796 159384
rect 404268 159332 404320 159384
rect 428004 159332 428056 159384
rect 385592 159264 385644 159316
rect 388352 159264 388404 159316
rect 401600 159264 401652 159316
rect 427820 159264 427872 159316
rect 446036 159332 446088 159384
rect 453028 159332 453080 159384
rect 465264 159332 465316 159384
rect 468116 159332 468168 159384
rect 474740 159332 474792 159384
rect 477316 159332 477368 159384
rect 483112 159332 483164 159384
rect 518716 159332 518768 159384
rect 522672 159332 522724 159384
rect 90180 159196 90232 159248
rect 173256 159196 173308 159248
rect 173348 159196 173400 159248
rect 195244 159196 195296 159248
rect 196900 159196 196952 159248
rect 211804 159196 211856 159248
rect 213644 159196 213696 159248
rect 279792 159196 279844 159248
rect 281632 159196 281684 159248
rect 328460 159196 328512 159248
rect 332048 159196 332100 159248
rect 334532 159196 334584 159248
rect 335452 159196 335504 159248
rect 375380 159196 375432 159248
rect 391664 159196 391716 159248
rect 403900 159196 403952 159248
rect 457168 159196 457220 159248
rect 464620 159196 464672 159248
rect 63316 159128 63368 159180
rect 102140 159128 102192 159180
rect 103612 159128 103664 159180
rect 183100 159128 183152 159180
rect 193496 159128 193548 159180
rect 223580 159128 223632 159180
rect 234620 159128 234672 159180
rect 298376 159128 298428 159180
rect 301872 159128 301924 159180
rect 349712 159128 349764 159180
rect 80152 159060 80204 159112
rect 89720 159060 89772 159112
rect 96896 159060 96948 159112
rect 173992 159060 174044 159112
rect 174084 159060 174136 159112
rect 179052 159060 179104 159112
rect 180800 159060 180852 159112
rect 181628 159060 181680 159112
rect 186780 159060 186832 159112
rect 214564 159060 214616 159112
rect 220360 159060 220412 159112
rect 229376 159060 229428 159112
rect 230480 159060 230532 159112
rect 294512 159060 294564 159112
rect 300952 159060 301004 159112
rect 349068 159060 349120 159112
rect 92756 158992 92808 159044
rect 116032 158992 116084 159044
rect 116124 158992 116176 159044
rect 118700 158992 118752 159044
rect 119620 158992 119672 159044
rect 133788 158992 133840 159044
rect 133880 158992 133932 159044
rect 210240 158992 210292 159044
rect 210332 158992 210384 159044
rect 214012 158992 214064 159044
rect 214380 158992 214432 159044
rect 215392 158992 215444 159044
rect 224224 158992 224276 159044
rect 227720 158992 227772 159044
rect 233792 158992 233844 159044
rect 291660 158992 291712 159044
rect 291752 158992 291804 159044
rect 293960 158992 294012 159044
rect 298468 158992 298520 159044
rect 299480 158992 299532 159044
rect 306840 158992 306892 159044
rect 353300 159128 353352 159180
rect 353852 159128 353904 159180
rect 357716 159128 357768 159180
rect 357808 159128 357860 159180
rect 387616 159128 387668 159180
rect 392492 159128 392544 159180
rect 415676 159128 415728 159180
rect 461400 159128 461452 159180
rect 468024 159128 468076 159180
rect 349988 159060 350040 159112
rect 377772 159060 377824 159112
rect 350080 158992 350132 159044
rect 354864 158992 354916 159044
rect 113640 158924 113692 158976
rect 120080 158924 120132 158976
rect 120448 158924 120500 158976
rect 106188 158856 106240 158908
rect 122564 158856 122616 158908
rect 122748 158924 122800 158976
rect 186412 158924 186464 158976
rect 195244 158924 195296 158976
rect 194508 158856 194560 158908
rect 195336 158856 195388 158908
rect 198740 158856 198792 158908
rect 203616 158924 203668 158976
rect 233148 158924 233200 158976
rect 240508 158924 240560 158976
rect 300860 158924 300912 158976
rect 310244 158924 310296 158976
rect 310704 158924 310756 158976
rect 313556 158924 313608 158976
rect 357624 158992 357676 159044
rect 357716 158992 357768 159044
rect 380900 159060 380952 159112
rect 390836 159060 390888 159112
rect 391940 159060 391992 159112
rect 422760 159060 422812 159112
rect 424968 159060 425020 159112
rect 460572 159060 460624 159112
rect 466460 159060 466512 159112
rect 473176 159060 473228 159112
rect 478880 159060 478932 159112
rect 481548 159060 481600 159112
rect 487252 159060 487304 159112
rect 204076 158856 204128 158908
rect 206928 158856 206980 158908
rect 233884 158856 233936 158908
rect 253940 158856 253992 158908
rect 311992 158856 312044 158908
rect 318616 158856 318668 158908
rect 319168 158856 319220 158908
rect 102784 158788 102836 158840
rect 123944 158788 123996 158840
rect 124036 158788 124088 158840
rect 135168 158788 135220 158840
rect 136272 158788 136324 158840
rect 196072 158788 196124 158840
rect 200212 158788 200264 158840
rect 224224 158788 224276 158840
rect 224592 158788 224644 158840
rect 230756 158788 230808 158840
rect 243912 158788 243964 158840
rect 246120 158788 246172 158840
rect 261484 158788 261536 158840
rect 318708 158788 318760 158840
rect 99472 158720 99524 158772
rect 113640 158720 113692 158772
rect 113732 158720 113784 158772
rect 122748 158720 122800 158772
rect 122932 158720 122984 158772
rect 142988 158720 143040 158772
rect 143080 158720 143132 158772
rect 176476 158720 176528 158772
rect 180064 158720 180116 158772
rect 202880 158720 202932 158772
rect 204444 158720 204496 158772
rect 219900 158720 219952 158772
rect 227076 158720 227128 158772
rect 241428 158720 241480 158772
rect 244740 158720 244792 158772
rect 245752 158720 245804 158772
rect 251456 158720 251508 158772
rect 252928 158720 252980 158772
rect 268200 158720 268252 158772
rect 324044 158856 324096 158908
rect 324412 158856 324464 158908
rect 328460 158856 328512 158908
rect 328644 158856 328696 158908
rect 365168 158924 365220 158976
rect 371516 158924 371568 158976
rect 382464 158992 382516 159044
rect 411352 158992 411404 159044
rect 463056 158992 463108 159044
rect 469220 158992 469272 159044
rect 471428 158992 471480 159044
rect 477592 158992 477644 159044
rect 397368 158924 397420 158976
rect 419356 158924 419408 158976
rect 423496 158924 423548 158976
rect 465632 158924 465684 158976
rect 472532 158924 472584 158976
rect 474832 158924 474884 158976
rect 481640 158924 481692 158976
rect 506572 158924 506624 158976
rect 508412 158924 508464 158976
rect 516692 158924 516744 158976
rect 520188 158924 520240 158976
rect 363052 158856 363104 158908
rect 363972 158856 364024 158908
rect 385868 158856 385920 158908
rect 411812 158856 411864 158908
rect 413744 158856 413796 158908
rect 455512 158856 455564 158908
rect 463608 158856 463660 158908
rect 464712 158856 464764 158908
rect 471428 158856 471480 158908
rect 474004 158856 474056 158908
rect 481364 158856 481416 158908
rect 508320 158856 508372 158908
rect 509240 158856 509292 158908
rect 509332 158856 509384 158908
rect 511816 158856 511868 158908
rect 515036 158856 515088 158908
rect 518532 158856 518584 158908
rect 320272 158720 320324 158772
rect 357256 158788 357308 158840
rect 380992 158788 381044 158840
rect 398380 158788 398432 158840
rect 404636 158788 404688 158840
rect 408500 158788 408552 158840
rect 411260 158788 411312 158840
rect 456340 158788 456392 158840
rect 463516 158788 463568 158840
rect 463884 158788 463936 158840
rect 471520 158788 471572 158840
rect 507952 158788 508004 158840
rect 510068 158788 510120 158840
rect 512184 158788 512236 158840
rect 514300 158788 514352 158840
rect 514852 158788 514904 158840
rect 517612 158788 517664 158840
rect 322020 158720 322072 158772
rect 80980 158652 81032 158704
rect 180800 158652 180852 158704
rect 181720 158652 181772 158704
rect 256792 158652 256844 158704
rect 327908 158720 327960 158772
rect 328644 158652 328696 158704
rect 367376 158720 367428 158772
rect 386052 158720 386104 158772
rect 387524 158720 387576 158772
rect 390560 158720 390612 158772
rect 405096 158720 405148 158772
rect 408868 158720 408920 158772
rect 412640 158720 412692 158772
rect 419540 158720 419592 158772
rect 462228 158720 462280 158772
rect 467932 158720 467984 158772
rect 475660 158720 475712 158772
rect 482652 158720 482704 158772
rect 505284 158720 505336 158772
rect 506756 158720 506808 158772
rect 509608 158720 509660 158772
rect 510896 158720 510948 158772
rect 510988 158720 511040 158772
rect 512644 158720 512696 158772
rect 513564 158720 513616 158772
rect 515956 158720 516008 158772
rect 368480 158652 368532 158704
rect 70860 158584 70912 158636
rect 172704 158584 172756 158636
rect 175004 158584 175056 158636
rect 252744 158584 252796 158636
rect 74264 158516 74316 158568
rect 175372 158516 175424 158568
rect 178408 158516 178460 158568
rect 255412 158516 255464 158568
rect 60832 158448 60884 158500
rect 164332 158448 164384 158500
rect 164424 158448 164476 158500
rect 242440 158448 242492 158500
rect 64144 158380 64196 158432
rect 162124 158380 162176 158432
rect 67548 158312 67600 158364
rect 162308 158312 162360 158364
rect 167552 158312 167604 158364
rect 168288 158380 168340 158432
rect 247592 158380 247644 158432
rect 170588 158312 170640 158364
rect 171692 158312 171744 158364
rect 249892 158312 249944 158364
rect 54116 158244 54168 158296
rect 153016 158244 153068 158296
rect 47400 158176 47452 158228
rect 153108 158176 153160 158228
rect 157432 158244 157484 158296
rect 158260 158244 158312 158296
rect 161940 158244 161992 158296
rect 162216 158244 162268 158296
rect 164884 158244 164936 158296
rect 164976 158244 165028 158296
rect 245016 158244 245068 158296
rect 50712 158108 50764 158160
rect 154856 158176 154908 158228
rect 164608 158176 164660 158228
rect 164792 158176 164844 158228
rect 237472 158176 237524 158228
rect 249800 158176 249852 158228
rect 309876 158176 309928 158228
rect 153476 158108 153528 158160
rect 155132 158108 155184 158160
rect 155224 158108 155276 158160
rect 160100 158108 160152 158160
rect 161572 158108 161624 158160
rect 164424 158108 164476 158160
rect 164884 158108 164936 158160
rect 238852 158108 238904 158160
rect 246396 158108 246448 158160
rect 307300 158108 307352 158160
rect 37280 158040 37332 158092
rect 146300 158040 146352 158092
rect 148140 158040 148192 158092
rect 231952 158040 232004 158092
rect 239680 158040 239732 158092
rect 302332 158040 302384 158092
rect 388 157972 440 158024
rect 118884 157972 118936 158024
rect 134708 157972 134760 158024
rect 221924 157972 221976 158024
rect 236368 157972 236420 158024
rect 299664 157972 299716 158024
rect 77576 157904 77628 157956
rect 178040 157904 178092 157956
rect 87696 157836 87748 157888
rect 185308 157904 185360 157956
rect 188436 157904 188488 157956
rect 263048 157904 263100 157956
rect 91008 157768 91060 157820
rect 188528 157836 188580 157888
rect 190092 157836 190144 157888
rect 264336 157836 264388 157888
rect 181536 157768 181588 157820
rect 191104 157768 191156 157820
rect 195152 157768 195204 157820
rect 267740 157768 267792 157820
rect 84292 157700 84344 157752
rect 182364 157700 182416 157752
rect 185124 157700 185176 157752
rect 260472 157700 260524 157752
rect 94412 157632 94464 157684
rect 181536 157632 181588 157684
rect 181628 157632 181680 157684
rect 200304 157632 200356 157684
rect 202880 157632 202932 157684
rect 255872 157632 255924 157684
rect 111156 157564 111208 157616
rect 200580 157564 200632 157616
rect 200764 157564 200816 157616
rect 203984 157564 204036 157616
rect 204076 157564 204128 157616
rect 251456 157564 251508 157616
rect 107844 157496 107896 157548
rect 200212 157496 200264 157548
rect 200304 157496 200356 157548
rect 233516 157496 233568 157548
rect 117872 157428 117924 157480
rect 209136 157428 209188 157480
rect 233148 157428 233200 157480
rect 273812 157428 273864 157480
rect 107016 157360 107068 157412
rect 107752 157360 107804 157412
rect 141424 157360 141476 157412
rect 226892 157360 226944 157412
rect 45652 157292 45704 157344
rect 153844 157292 153896 157344
rect 191840 157292 191892 157344
rect 265164 157292 265216 157344
rect 49056 157224 49108 157276
rect 156420 157224 156472 157276
rect 156604 157224 156656 157276
rect 219992 157224 220044 157276
rect 283380 157224 283432 157276
rect 335544 157224 335596 157276
rect 38936 157156 38988 157208
rect 148784 157156 148836 157208
rect 151820 157156 151872 157208
rect 152924 157156 152976 157208
rect 158720 157156 158772 157208
rect 166172 157156 166224 157208
rect 166264 157156 166316 157208
rect 171140 157156 171192 157208
rect 172428 157156 172480 157208
rect 179696 157156 179748 157208
rect 183376 157156 183428 157208
rect 258172 157156 258224 157208
rect 273260 157156 273312 157208
rect 327632 157156 327684 157208
rect 31392 157088 31444 157140
rect 142988 157088 143040 157140
rect 151544 157088 151596 157140
rect 234804 157088 234856 157140
rect 279976 157088 280028 157140
rect 333060 157088 333112 157140
rect 28080 157020 28132 157072
rect 139952 157020 140004 157072
rect 142252 157020 142304 157072
rect 227812 157020 227864 157072
rect 276664 157020 276716 157072
rect 330484 157020 330536 157072
rect 24676 156952 24728 157004
rect 137192 156952 137244 157004
rect 144828 156952 144880 157004
rect 229560 156952 229612 157004
rect 232964 156952 233016 157004
rect 297088 156952 297140 157004
rect 17960 156884 18012 156936
rect 132684 156884 132736 156936
rect 138112 156884 138164 156936
rect 224500 156884 224552 156936
rect 229652 156884 229704 156936
rect 294052 156884 294104 156936
rect 296812 156884 296864 156936
rect 345848 156884 345900 156936
rect 21364 156816 21416 156868
rect 135260 156816 135312 156868
rect 135536 156816 135588 156868
rect 222568 156816 222620 156868
rect 222844 156816 222896 156868
rect 289360 156816 289412 156868
rect 300124 156816 300176 156868
rect 348056 156816 348108 156868
rect 127992 156748 128044 156800
rect 216864 156748 216916 156800
rect 219532 156748 219584 156800
rect 286784 156748 286836 156800
rect 290096 156748 290148 156800
rect 339684 156748 339736 156800
rect 14648 156680 14700 156732
rect 130108 156680 130160 156732
rect 138940 156680 138992 156732
rect 225144 156680 225196 156732
rect 293408 156680 293460 156732
rect 343272 156680 343324 156732
rect 2044 156612 2096 156664
rect 120448 156612 120500 156664
rect 121276 156612 121328 156664
rect 211344 156612 211396 156664
rect 216128 156612 216180 156664
rect 284208 156612 284260 156664
rect 286692 156612 286744 156664
rect 338212 156612 338264 156664
rect 521844 156612 521896 156664
rect 523500 156612 523552 156664
rect 69204 156544 69256 156596
rect 166264 156544 166316 156596
rect 166356 156544 166408 156596
rect 175924 156544 175976 156596
rect 79324 156476 79376 156528
rect 179604 156544 179656 156596
rect 179696 156544 179748 156596
rect 191012 156544 191064 156596
rect 191196 156544 191248 156596
rect 176200 156476 176252 156528
rect 12072 156408 12124 156460
rect 109040 156408 109092 156460
rect 115388 156408 115440 156460
rect 187884 156408 187936 156460
rect 89352 156340 89404 156392
rect 187240 156340 187292 156392
rect 97724 156272 97776 156324
rect 193680 156340 193732 156392
rect 200672 156544 200724 156596
rect 198556 156476 198608 156528
rect 200856 156476 200908 156528
rect 201868 156544 201920 156596
rect 273260 156544 273312 156596
rect 202696 156476 202748 156528
rect 206100 156476 206152 156528
rect 276020 156476 276072 156528
rect 207204 156408 207256 156460
rect 209412 156408 209464 156460
rect 279056 156408 279108 156460
rect 225788 156340 225840 156392
rect 226248 156340 226300 156392
rect 291936 156340 291988 156392
rect 191012 156272 191064 156324
rect 238668 156272 238720 156324
rect 15476 156204 15528 156256
rect 109684 156204 109736 156256
rect 114560 156204 114612 156256
rect 206560 156204 206612 156256
rect 211804 156204 211856 156256
rect 269488 156204 269540 156256
rect 109500 156136 109552 156188
rect 200672 156136 200724 156188
rect 200764 156136 200816 156188
rect 213920 156136 213972 156188
rect 124588 156068 124640 156120
rect 214196 156068 214248 156120
rect 214564 156068 214616 156120
rect 260840 156136 260892 156188
rect 223580 156068 223632 156120
rect 266452 156068 266504 156120
rect 125508 156000 125560 156052
rect 200764 156000 200816 156052
rect 200856 156000 200908 156052
rect 270592 156000 270644 156052
rect 11244 155932 11296 155984
rect 127440 155932 127492 155984
rect 131396 155932 131448 155984
rect 218244 155932 218296 155984
rect 75920 155864 75972 155916
rect 177028 155864 177080 155916
rect 179236 155864 179288 155916
rect 255688 155864 255740 155916
rect 292580 155864 292632 155916
rect 342352 155864 342404 155916
rect 75092 155796 75144 155848
rect 176384 155796 176436 155848
rect 176476 155796 176528 155848
rect 185676 155796 185728 155848
rect 185952 155796 186004 155848
rect 261116 155796 261168 155848
rect 299296 155796 299348 155848
rect 347872 155796 347924 155848
rect 43168 155728 43220 155780
rect 75828 155728 75880 155780
rect 78404 155728 78456 155780
rect 178960 155728 179012 155780
rect 179052 155728 179104 155780
rect 185768 155728 185820 155780
rect 185860 155728 185912 155780
rect 258540 155728 258592 155780
rect 295984 155728 296036 155780
rect 345204 155728 345256 155780
rect 46572 155660 46624 155712
rect 69664 155660 69716 155712
rect 71688 155660 71740 155712
rect 173072 155660 173124 155712
rect 173164 155660 173216 155712
rect 250812 155660 250864 155712
rect 289268 155660 289320 155712
rect 340052 155660 340104 155712
rect 36452 155592 36504 155644
rect 63500 155592 63552 155644
rect 64972 155592 65024 155644
rect 168656 155592 168708 155644
rect 169116 155592 169168 155644
rect 247132 155592 247184 155644
rect 269948 155592 270000 155644
rect 325332 155592 325384 155644
rect 51540 155524 51592 155576
rect 158352 155524 158404 155576
rect 159088 155524 159140 155576
rect 240600 155524 240652 155576
rect 266544 155524 266596 155576
rect 321836 155524 321888 155576
rect 340420 155524 340472 155576
rect 379244 155524 379296 155576
rect 54944 155456 54996 155508
rect 160928 155456 160980 155508
rect 162400 155456 162452 155508
rect 243084 155456 243136 155508
rect 263232 155456 263284 155508
rect 320180 155456 320232 155508
rect 337108 155456 337160 155508
rect 376668 155456 376720 155508
rect 48228 155388 48280 155440
rect 151728 155388 151780 155440
rect 152740 155388 152792 155440
rect 155592 155388 155644 155440
rect 155684 155388 155736 155440
rect 237564 155388 237616 155440
rect 259828 155388 259880 155440
rect 317604 155388 317656 155440
rect 332876 155388 332928 155440
rect 373448 155388 373500 155440
rect 4528 155320 4580 155372
rect 122012 155320 122064 155372
rect 123760 155320 123812 155372
rect 128452 155320 128504 155372
rect 148968 155320 149020 155372
rect 232872 155320 232924 155372
rect 256516 155320 256568 155372
rect 315028 155320 315080 155372
rect 329564 155320 329616 155372
rect 370872 155320 370924 155372
rect 376576 155320 376628 155372
rect 406844 155320 406896 155372
rect 8760 155252 8812 155304
rect 125600 155252 125652 155304
rect 132224 155252 132276 155304
rect 219532 155252 219584 155304
rect 243176 155252 243228 155304
rect 5356 155184 5408 155236
rect 123024 155184 123076 155236
rect 128820 155184 128872 155236
rect 217416 155184 217468 155236
rect 233884 155184 233936 155236
rect 243544 155184 243596 155236
rect 253112 155252 253164 155304
rect 312452 155252 312504 155304
rect 373172 155252 373224 155304
rect 403164 155252 403216 155304
rect 304724 155184 304776 155236
rect 306012 155184 306064 155236
rect 352932 155184 352984 155236
rect 369860 155184 369912 155236
rect 401692 155184 401744 155236
rect 56600 155116 56652 155168
rect 76472 155116 76524 155168
rect 81808 155116 81860 155168
rect 181352 155116 181404 155168
rect 182548 155116 182600 155168
rect 185400 155116 185452 155168
rect 185492 155116 185544 155168
rect 73436 155048 73488 155100
rect 81440 155048 81492 155100
rect 88524 155048 88576 155100
rect 186596 155048 186648 155100
rect 189264 155116 189316 155168
rect 263784 155116 263836 155168
rect 302700 155116 302752 155168
rect 349344 155116 349396 155168
rect 192392 155048 192444 155100
rect 192668 155048 192720 155100
rect 266268 155048 266320 155100
rect 312728 155048 312780 155100
rect 357900 155048 357952 155100
rect 91836 154980 91888 155032
rect 189172 154980 189224 155032
rect 195980 154980 196032 155032
rect 268844 154980 268896 155032
rect 86040 154912 86092 154964
rect 183560 154912 183612 154964
rect 185584 154912 185636 154964
rect 191748 154912 191800 154964
rect 199384 154912 199436 154964
rect 271420 154912 271472 154964
rect 96068 154844 96120 154896
rect 185492 154844 185544 154896
rect 185676 154844 185728 154896
rect 98644 154776 98696 154828
rect 194324 154776 194376 154828
rect 202788 154844 202840 154896
rect 273444 154844 273496 154896
rect 228364 154776 228416 154828
rect 95240 154708 95292 154760
rect 185584 154708 185636 154760
rect 185768 154708 185820 154760
rect 229652 154708 229704 154760
rect 118792 154640 118844 154692
rect 209780 154640 209832 154692
rect 212816 154640 212868 154692
rect 281632 154776 281684 154828
rect 229836 154708 229888 154760
rect 242900 154708 242952 154760
rect 243544 154708 243596 154760
rect 276480 154708 276532 154760
rect 241428 154640 241480 154692
rect 292580 154640 292632 154692
rect 122104 154572 122156 154624
rect 212264 154572 212316 154624
rect 227720 154572 227772 154624
rect 272064 154572 272116 154624
rect 58348 154504 58400 154556
rect 44180 154436 44232 154488
rect 146760 154436 146812 154488
rect 147036 154436 147088 154488
rect 148324 154436 148376 154488
rect 41512 154368 41564 154420
rect 146576 154368 146628 154420
rect 146944 154368 146996 154420
rect 152372 154368 152424 154420
rect 152740 154504 152792 154556
rect 210516 154504 210568 154556
rect 215300 154504 215352 154556
rect 283196 154504 283248 154556
rect 285864 154504 285916 154556
rect 337476 154504 337528 154556
rect 352288 154504 352340 154556
rect 388904 154504 388956 154556
rect 153016 154436 153068 154488
rect 207848 154436 207900 154488
rect 211252 154436 211304 154488
rect 280988 154436 281040 154488
rect 281724 154436 281776 154488
rect 334900 154436 334952 154488
rect 349252 154436 349304 154488
rect 386328 154436 386380 154488
rect 163320 154368 163372 154420
rect 164148 154368 164200 154420
rect 165712 154368 165764 154420
rect 165804 154368 165856 154420
rect 175924 154368 175976 154420
rect 176016 154368 176068 154420
rect 181260 154368 181312 154420
rect 181996 154368 182048 154420
rect 254032 154368 254084 154420
rect 258264 154368 258316 154420
rect 316960 154368 317012 154420
rect 345572 154368 345624 154420
rect 383844 154368 383896 154420
rect 116032 154300 116084 154352
rect 121920 154300 121972 154352
rect 123944 154300 123996 154352
rect 127348 154300 127400 154352
rect 127532 154300 127584 154352
rect 189816 154300 189868 154352
rect 191196 154300 191248 154352
rect 202052 154300 202104 154352
rect 208584 154300 208636 154352
rect 278412 154300 278464 154352
rect 278780 154300 278832 154352
rect 332416 154300 332468 154352
rect 342260 154300 342312 154352
rect 381176 154300 381228 154352
rect 400312 154300 400364 154352
rect 425520 154300 425572 154352
rect 30564 154232 30616 154284
rect 137284 154232 137336 154284
rect 26884 154164 26936 154216
rect 136088 154164 136140 154216
rect 189540 154232 189592 154284
rect 191012 154232 191064 154284
rect 199476 154232 199528 154284
rect 204536 154232 204588 154284
rect 274640 154232 274692 154284
rect 275100 154232 275152 154284
rect 329932 154232 329984 154284
rect 339592 154232 339644 154284
rect 378600 154232 378652 154284
rect 393412 154232 393464 154284
rect 419724 154232 419776 154284
rect 23480 154096 23532 154148
rect 137100 154096 137152 154148
rect 13820 154028 13872 154080
rect 129464 154028 129516 154080
rect 129556 154028 129608 154080
rect 139492 154164 139544 154216
rect 146944 154164 146996 154216
rect 147128 154164 147180 154216
rect 137560 154096 137612 154148
rect 146852 154096 146904 154148
rect 148232 154164 148284 154216
rect 153200 154164 153252 154216
rect 154488 154164 154540 154216
rect 175832 154164 175884 154216
rect 176108 154164 176160 154216
rect 253388 154164 253440 154216
rect 255320 154164 255372 154216
rect 314384 154164 314436 154216
rect 335636 154164 335688 154216
rect 376024 154164 376076 154216
rect 386604 154164 386656 154216
rect 414572 154164 414624 154216
rect 166264 154096 166316 154148
rect 166356 154096 166408 154148
rect 175740 154096 175792 154148
rect 175924 154096 175976 154148
rect 245660 154096 245712 154148
rect 248420 154096 248472 154148
rect 309232 154096 309284 154148
rect 325700 154096 325752 154148
rect 368296 154096 368348 154148
rect 389732 154096 389784 154148
rect 417148 154096 417200 154148
rect 137284 154028 137336 154080
rect 142344 154028 142396 154080
rect 144920 154028 144972 154080
rect 16580 153960 16632 154012
rect 132040 153960 132092 154012
rect 136088 153960 136140 154012
rect 139768 153960 139820 154012
rect 480 153892 532 153944
rect 119804 153892 119856 153944
rect 120080 153892 120132 153944
rect 2964 153824 3016 153876
rect 121736 153824 121788 153876
rect 121920 153892 121972 153944
rect 127532 153892 127584 153944
rect 146668 153892 146720 153944
rect 146760 153892 146812 153944
rect 147772 153892 147824 153944
rect 152924 154028 152976 154080
rect 235448 154028 235500 154080
rect 245568 154028 245620 154080
rect 306656 154028 306708 154080
rect 316132 154028 316184 154080
rect 360660 154028 360712 154080
rect 363144 154028 363196 154080
rect 396540 154028 396592 154080
rect 400128 154028 400180 154080
rect 424876 154028 424928 154080
rect 148324 153960 148376 154012
rect 230940 153960 230992 154012
rect 231860 153960 231912 154012
rect 296444 153960 296496 154012
rect 322848 153960 322900 154012
rect 365812 153960 365864 154012
rect 379612 153960 379664 154012
rect 409420 153960 409472 154012
rect 230296 153892 230348 153944
rect 234712 153892 234764 153944
rect 299020 153892 299072 153944
rect 318800 153892 318852 153944
rect 363144 153892 363196 153944
rect 383292 153892 383344 153944
rect 411996 153892 412048 153944
rect 421104 153892 421156 153944
rect 440884 153892 440936 153944
rect 128360 153824 128412 153876
rect 215484 153824 215536 153876
rect 218060 153824 218112 153876
rect 286140 153824 286192 153876
rect 309140 153824 309192 153876
rect 355508 153824 355560 153876
rect 356060 153824 356112 153876
rect 391480 153824 391532 153876
rect 396080 153824 396132 153876
rect 422300 153824 422352 153876
rect 62120 153756 62172 153808
rect 166172 153756 166224 153808
rect 166264 153756 166316 153808
rect 212908 153756 212960 153808
rect 224960 153756 225012 153808
rect 291292 153756 291344 153808
rect 359004 153756 359056 153808
rect 394056 153756 394108 153808
rect 425244 153756 425296 153808
rect 432696 153756 432748 153808
rect 71780 153688 71832 153740
rect 173900 153688 173952 153740
rect 175832 153688 175884 153740
rect 218060 153688 218112 153740
rect 227996 153688 228048 153740
rect 293868 153688 293920 153740
rect 365720 153688 365772 153740
rect 399116 153688 399168 153740
rect 81900 153620 81952 153672
rect 175648 153620 175700 153672
rect 175740 153620 175792 153672
rect 223212 153620 223264 153672
rect 241520 153620 241572 153672
rect 304080 153620 304132 153672
rect 101312 153552 101364 153604
rect 104900 153484 104952 153536
rect 191012 153484 191064 153536
rect 191288 153552 191340 153604
rect 236092 153552 236144 153604
rect 238944 153552 238996 153604
rect 301596 153552 301648 153604
rect 196900 153484 196952 153536
rect 198740 153484 198792 153536
rect 248880 153484 248932 153536
rect 251548 153484 251600 153536
rect 311808 153484 311860 153536
rect 107936 153416 107988 153468
rect 191196 153416 191248 153468
rect 191288 153416 191340 153468
rect 194968 153416 195020 153468
rect 196164 153416 196216 153468
rect 241244 153416 241296 153468
rect 264980 153416 265032 153468
rect 321744 153416 321796 153468
rect 426164 153416 426216 153468
rect 429476 153416 429528 153468
rect 111800 153348 111852 153400
rect 204628 153348 204680 153400
rect 262404 153348 262456 153400
rect 319536 153348 319588 153400
rect 112260 153280 112312 153332
rect 205272 153280 205324 153332
rect 269120 153280 269172 153332
rect 274548 153280 274600 153332
rect 274640 153280 274692 153332
rect 275836 153280 275888 153332
rect 275928 153280 275980 153332
rect 324688 153280 324740 153332
rect 34520 153212 34572 153264
rect 145564 153212 145616 153264
rect 146668 153212 146720 153264
rect 189448 153212 189500 153264
rect 189540 153212 189592 153264
rect 197544 153212 197596 153264
rect 197636 153212 197688 153264
rect 246304 153212 246356 153264
rect 271972 153212 272024 153264
rect 327264 153212 327316 153264
rect 360844 153212 360896 153264
rect 107752 153144 107804 153196
rect 200764 153144 200816 153196
rect 218152 153144 218204 153196
rect 226248 153144 226300 153196
rect 226340 153144 226392 153196
rect 231584 153144 231636 153196
rect 237196 153144 237248 153196
rect 300308 153144 300360 153196
rect 300860 153144 300912 153196
rect 302884 153144 302936 153196
rect 303620 153144 303672 153196
rect 351644 153144 351696 153196
rect 354772 153144 354824 153196
rect 364984 153144 365036 153196
rect 395160 153144 395212 153196
rect 395528 153144 395580 153196
rect 397828 153144 397880 153196
rect 401600 153144 401652 153196
rect 415860 153144 415912 153196
rect 416964 153144 417016 153196
rect 438308 153144 438360 153196
rect 438860 153144 438912 153196
rect 442448 153144 442500 153196
rect 442908 153144 442960 153196
rect 457628 153144 457680 153196
rect 458180 153144 458232 153196
rect 460756 153144 460808 153196
rect 463608 153144 463660 153196
rect 467196 153144 467248 153196
rect 471520 153144 471572 153196
rect 473636 153144 473688 153196
rect 474740 153144 474792 153196
rect 476856 153144 476908 153196
rect 477592 153144 477644 153196
rect 479340 153144 479392 153196
rect 483204 153144 483256 153196
rect 488448 153144 488500 153196
rect 489920 153144 489972 153196
rect 493508 153144 493560 153196
rect 494152 153144 494204 153196
rect 496728 153144 496780 153196
rect 496820 153144 496872 153196
rect 499304 153144 499356 153196
rect 500868 153144 500920 153196
rect 501880 153144 501932 153196
rect 503352 153144 503404 153196
rect 503812 153144 503864 153196
rect 511632 153144 511684 153196
rect 513472 153144 513524 153196
rect 514208 153144 514260 153196
rect 516140 153144 516192 153196
rect 30196 153076 30248 153128
rect 110972 153076 111024 153128
rect 116400 153076 116452 153128
rect 208492 153076 208544 153128
rect 214012 153076 214064 153128
rect 279332 153076 279384 153128
rect 279792 153076 279844 153128
rect 282276 153076 282328 153128
rect 284300 153076 284352 153128
rect 336832 153076 336884 153128
rect 337016 153076 337068 153128
rect 338764 153076 338816 153128
rect 340880 153076 340932 153128
rect 379888 153076 379940 153128
rect 384948 153076 385000 153128
rect 413100 153076 413152 153128
rect 414112 153076 414164 153128
rect 431868 153076 431920 153128
rect 431960 153076 432012 153128
rect 432788 153076 432840 153128
rect 437940 153076 437992 153128
rect 454408 153076 454460 153128
rect 463516 153076 463568 153128
rect 467840 153076 467892 153128
rect 471428 153076 471480 153128
rect 474280 153076 474332 153128
rect 475016 153076 475068 153128
rect 477500 153076 477552 153128
rect 484400 153076 484452 153128
rect 489644 153076 489696 153128
rect 491300 153076 491352 153128
rect 494796 153076 494848 153128
rect 495440 153076 495492 153128
rect 498016 153076 498068 153128
rect 500960 153076 501012 153128
rect 502524 153076 502576 153128
rect 512920 153076 512972 153128
rect 515128 153076 515180 153128
rect 23296 153008 23348 153060
rect 108028 153008 108080 153060
rect 110328 153008 110380 153060
rect 203340 153008 203392 153060
rect 210240 153008 210292 153060
rect 221280 153008 221332 153060
rect 230572 153008 230624 153060
rect 295800 153008 295852 153060
rect 305184 153008 305236 153060
rect 352288 153008 352340 153060
rect 358912 153008 358964 153060
rect 364892 153008 364944 153060
rect 364984 153008 365036 153060
rect 390192 153008 390244 153060
rect 391940 153008 391992 153060
rect 417792 153008 417844 153060
rect 418160 153008 418212 153060
rect 438952 153008 439004 153060
rect 440424 153008 440476 153060
rect 455696 153008 455748 153060
rect 464620 153008 464672 153060
rect 468392 153008 468444 153060
rect 472532 153008 472584 153060
rect 474924 153008 474976 153060
rect 476120 153008 476172 153060
rect 478236 153008 478288 153060
rect 490012 153008 490064 153060
rect 494152 153008 494204 153060
rect 495992 153008 496044 153060
rect 498660 153008 498712 153060
rect 499672 153008 499724 153060
rect 501236 153008 501288 153060
rect 9496 152940 9548 152992
rect 92572 152940 92624 152992
rect 99564 152940 99616 152992
rect 195612 152940 195664 152992
rect 196072 152940 196124 152992
rect 216128 152940 216180 152992
rect 216680 152940 216732 152992
rect 284852 152940 284904 152992
rect 290188 152940 290240 152992
rect 341340 152940 341392 152992
rect 346400 152940 346452 152992
rect 93308 152872 93360 152924
rect 190460 152872 190512 152924
rect 194508 152872 194560 152924
rect 211068 152872 211120 152924
rect 211160 152872 211212 152924
rect 280344 152872 280396 152924
rect 284116 152872 284168 152924
rect 336188 152872 336240 152924
rect 338120 152872 338172 152924
rect 377956 152872 378008 152924
rect 380900 152872 380952 152924
rect 383200 152872 383252 152924
rect 383752 152940 383804 152992
rect 412640 152940 412692 152992
rect 415216 152940 415268 152992
rect 436376 152940 436428 152992
rect 436468 152940 436520 152992
rect 442356 152940 442408 152992
rect 442448 152940 442500 152992
rect 446772 152940 446824 152992
rect 464896 152940 464948 152992
rect 469128 152940 469180 152992
rect 473360 152940 473412 152992
rect 475568 152940 475620 152992
rect 494244 152940 494296 152992
rect 497372 152940 497424 152992
rect 384396 152872 384448 152924
rect 388444 152872 388496 152924
rect 408776 152872 408828 152924
rect 410708 152872 410760 152924
rect 433156 152872 433208 152924
rect 434720 152872 434772 152924
rect 451832 152872 451884 152924
rect 465356 152872 465408 152924
rect 469772 152872 469824 152924
rect 473452 152872 473504 152924
rect 476212 152872 476264 152924
rect 492680 152872 492732 152924
rect 496084 152872 496136 152924
rect 33140 152804 33192 152856
rect 137284 152804 137336 152856
rect 139400 152804 139452 152856
rect 141700 152804 141752 152856
rect 141792 152804 141844 152856
rect 146944 152804 146996 152856
rect 149060 152804 149112 152856
rect 164884 152804 164936 152856
rect 170036 152804 170088 152856
rect 249524 152804 249576 152856
rect 255504 152804 255556 152856
rect 257252 152804 257304 152856
rect 258080 152804 258132 152856
rect 316316 152804 316368 152856
rect 317144 152804 317196 152856
rect 318248 152804 318300 152856
rect 322940 152804 322992 152856
rect 366364 152804 366416 152856
rect 367560 152804 367612 152856
rect 26332 152736 26384 152788
rect 139124 152736 139176 152788
rect 139216 152736 139268 152788
rect 149428 152736 149480 152788
rect 152832 152736 152884 152788
rect 234160 152736 234212 152788
rect 237380 152736 237432 152788
rect 300952 152736 301004 152788
rect 303528 152736 303580 152788
rect 351000 152736 351052 152788
rect 351920 152736 351972 152788
rect 388260 152736 388312 152788
rect 395896 152804 395948 152856
rect 400404 152736 400456 152788
rect 405924 152804 405976 152856
rect 429292 152804 429344 152856
rect 429568 152804 429620 152856
rect 441068 152804 441120 152856
rect 421656 152736 421708 152788
rect 428648 152736 428700 152788
rect 446680 152804 446732 152856
rect 447692 152804 447744 152856
rect 461400 152804 461452 152856
rect 466552 152804 466604 152856
rect 470416 152804 470468 152856
rect 491760 152804 491812 152856
rect 495440 152804 495492 152856
rect 441252 152736 441304 152788
rect 444840 152736 444892 152788
rect 448888 152736 448940 152788
rect 462688 152736 462740 152788
rect 86132 152668 86184 152720
rect 185308 152668 185360 152720
rect 190552 152668 190604 152720
rect 264980 152668 265032 152720
rect 270868 152668 270920 152720
rect 326620 152668 326672 152720
rect 329840 152668 329892 152720
rect 361764 152668 361816 152720
rect 31760 152600 31812 152652
rect 143632 152600 143684 152652
rect 144460 152600 144512 152652
rect 159640 152600 159692 152652
rect 163504 152600 163556 152652
rect 244372 152600 244424 152652
rect 245752 152600 245804 152652
rect 306012 152600 306064 152652
rect 310612 152600 310664 152652
rect 356796 152600 356848 152652
rect 357532 152600 357584 152652
rect 359372 152600 359424 152652
rect 363236 152600 363288 152652
rect 364524 152600 364576 152652
rect 18052 152532 18104 152584
rect 133328 152532 133380 152584
rect 137284 152532 137336 152584
rect 144276 152532 144328 152584
rect 146944 152532 146996 152584
rect 157064 152532 157116 152584
rect 157340 152532 157392 152584
rect 239312 152532 239364 152584
rect 240324 152532 240376 152584
rect 241888 152532 241940 152584
rect 242992 152532 243044 152584
rect 246948 152532 247000 152584
rect 249984 152532 250036 152584
rect 310520 152532 310572 152584
rect 311900 152532 311952 152584
rect 357440 152532 357492 152584
rect 359464 152532 359516 152584
rect 367008 152668 367060 152720
rect 379060 152668 379112 152720
rect 388444 152668 388496 152720
rect 388536 152668 388588 152720
rect 407488 152668 407540 152720
rect 409052 152668 409104 152720
rect 431868 152668 431920 152720
rect 431960 152668 432012 152720
rect 434444 152668 434496 152720
rect 434536 152668 434588 152720
rect 446956 152668 447008 152720
rect 447048 152668 447100 152720
rect 452476 152668 452528 152720
rect 365076 152600 365128 152652
rect 393412 152600 393464 152652
rect 401876 152600 401928 152652
rect 426808 152600 426860 152652
rect 429200 152600 429252 152652
rect 447324 152600 447376 152652
rect 447416 152600 447468 152652
rect 451188 152600 451240 152652
rect 367100 152532 367152 152584
rect 394700 152532 394752 152584
rect 397552 152532 397604 152584
rect 422852 152532 422904 152584
rect 430580 152532 430632 152584
rect 12440 152464 12492 152516
rect 128820 152464 128872 152516
rect 129740 152464 129792 152516
rect 218704 152464 218756 152516
rect 223764 152464 223816 152516
rect 290004 152464 290056 152516
rect 297640 152464 297692 152516
rect 346492 152464 346544 152516
rect 347780 152464 347832 152516
rect 385040 152464 385092 152516
rect 394240 152464 394292 152516
rect 420368 152464 420420 152516
rect 423404 152464 423456 152516
rect 427084 152464 427136 152516
rect 81440 152396 81492 152448
rect 175096 152396 175148 152448
rect 176752 152396 176804 152448
rect 254676 152396 254728 152448
rect 256700 152396 256752 152448
rect 315672 152396 315724 152448
rect 317052 152396 317104 152448
rect 361304 152396 361356 152448
rect 361764 152396 361816 152448
rect 371516 152396 371568 152448
rect 89720 152328 89772 152380
rect 180248 152328 180300 152380
rect 185032 152328 185084 152380
rect 259828 152328 259880 152380
rect 263600 152328 263652 152380
rect 320824 152328 320876 152380
rect 321560 152328 321612 152380
rect 323400 152328 323452 152380
rect 324596 152328 324648 152380
rect 367652 152328 367704 152380
rect 367744 152328 367796 152380
rect 398472 152396 398524 152448
rect 398840 152396 398892 152448
rect 410708 152396 410760 152448
rect 413744 152396 413796 152448
rect 433800 152464 433852 152516
rect 434444 152464 434496 152516
rect 435732 152464 435784 152516
rect 429476 152396 429528 152448
rect 442080 152464 442132 152516
rect 371792 152328 371844 152380
rect 403624 152328 403676 152380
rect 403900 152328 403952 152380
rect 418436 152328 418488 152380
rect 421932 152328 421984 152380
rect 429752 152328 429804 152380
rect 76472 152260 76524 152312
rect 162216 152260 162268 152312
rect 167000 152260 167052 152312
rect 182824 152260 182876 152312
rect 186412 152260 186464 152312
rect 205916 152260 205968 152312
rect 230756 152260 230808 152312
rect 290648 152260 290700 152312
rect 293960 152260 294012 152312
rect 341984 152260 342036 152312
rect 345020 152260 345072 152312
rect 33600 152192 33652 152244
rect 109592 152192 109644 152244
rect 109684 152192 109736 152244
rect 130752 152192 130804 152244
rect 135168 152192 135220 152244
rect 139216 152192 139268 152244
rect 139308 152192 139360 152244
rect 141792 152192 141844 152244
rect 143540 152192 143592 152244
rect 229008 152192 229060 152244
rect 246120 152192 246172 152244
rect 305368 152192 305420 152244
rect 319168 152192 319220 152244
rect 362592 152192 362644 152244
rect 383108 152260 383160 152312
rect 383200 152260 383252 152312
rect 389548 152260 389600 152312
rect 390560 152260 390612 152312
rect 415216 152260 415268 152312
rect 415676 152260 415728 152312
rect 419080 152260 419132 152312
rect 370688 152192 370740 152244
rect 402336 152192 402388 152244
rect 408868 152192 408920 152244
rect 428648 152192 428700 152244
rect 429752 152192 429804 152244
rect 441528 152328 441580 152380
rect 445392 152532 445444 152584
rect 459468 152532 459520 152584
rect 442356 152464 442408 152516
rect 453120 152464 453172 152516
rect 488540 152464 488592 152516
rect 492864 152464 492916 152516
rect 442264 152396 442316 152448
rect 444748 152396 444800 152448
rect 444840 152396 444892 152448
rect 456340 152396 456392 152448
rect 448612 152328 448664 152380
rect 432696 152260 432748 152312
rect 444104 152260 444156 152312
rect 444564 152260 444616 152312
rect 458916 152260 458968 152312
rect 432788 152192 432840 152244
rect 449256 152192 449308 152244
rect 69664 152124 69716 152176
rect 154488 152124 154540 152176
rect 154580 152124 154632 152176
rect 169944 152124 169996 152176
rect 173992 152124 174044 152176
rect 193036 152124 193088 152176
rect 229376 152124 229428 152176
rect 287428 152124 287480 152176
rect 295340 152124 295392 152176
rect 297732 152124 297784 152176
rect 299480 152124 299532 152176
rect 347136 152124 347188 152176
rect 350540 152124 350592 152176
rect 386972 152124 387024 152176
rect 19800 152056 19852 152108
rect 99932 152056 99984 152108
rect 109040 152056 109092 152108
rect 128176 152056 128228 152108
rect 128452 152056 128504 152108
rect 213552 152056 213604 152108
rect 252928 152056 252980 152108
rect 311164 152056 311216 152108
rect 318892 152056 318944 152108
rect 361948 152056 362000 152108
rect 364800 152056 364852 152108
rect 367744 152056 367796 152108
rect 377772 152056 377824 152108
rect 381820 152056 381872 152108
rect 388536 152124 388588 152176
rect 388628 152124 388680 152176
rect 410064 152124 410116 152176
rect 411260 152124 411312 152176
rect 431224 152124 431276 152176
rect 433432 152124 433484 152176
rect 450544 152124 450596 152176
rect 63500 151988 63552 152040
rect 146852 151988 146904 152040
rect 158812 151988 158864 152040
rect 172520 151988 172572 152040
rect 183100 151988 183152 152040
rect 198188 151988 198240 152040
rect 264152 151988 264204 152040
rect 321468 151988 321520 152040
rect 331312 151988 331364 152040
rect 334348 151988 334400 152040
rect 75828 151920 75880 151972
rect 74816 151852 74868 151904
rect 82084 151852 82136 151904
rect 105820 151920 105872 151972
rect 110328 151920 110380 151972
rect 127256 151920 127308 151972
rect 135904 151920 135956 151972
rect 142896 151920 142948 151972
rect 223856 151920 223908 151972
rect 278044 151920 278096 151972
rect 331772 151920 331824 151972
rect 151912 151852 151964 151904
rect 164516 151852 164568 151904
rect 71412 151784 71464 151836
rect 91008 151784 91060 151836
rect 102140 151784 102192 151836
rect 167368 151784 167420 151836
rect 173256 151852 173308 151904
rect 187884 151852 187936 151904
rect 219900 151852 219952 151904
rect 275192 151852 275244 151904
rect 276112 151852 276164 151904
rect 277768 151852 277820 151904
rect 280160 151852 280212 151904
rect 331128 151852 331180 151904
rect 359464 151988 359516 152040
rect 360200 151988 360252 152040
rect 367100 151988 367152 152040
rect 177672 151784 177724 151836
rect 215392 151784 215444 151836
rect 270132 151784 270184 151836
rect 273352 151784 273404 151836
rect 325976 151784 326028 151836
rect 328368 151784 328420 151836
rect 334532 151852 334584 151904
rect 372804 151920 372856 151972
rect 376760 151920 376812 151972
rect 408132 152056 408184 152108
rect 418252 152056 418304 152108
rect 424232 152056 424284 152108
rect 339500 151852 339552 151904
rect 377312 151852 377364 151904
rect 378232 151852 378284 151904
rect 388720 151988 388772 152040
rect 404912 151988 404964 152040
rect 407580 151988 407632 152040
rect 426164 151988 426216 152040
rect 442172 152056 442224 152108
rect 443000 152056 443052 152108
rect 458180 152056 458232 152108
rect 485872 152056 485924 152108
rect 490932 152056 490984 152108
rect 386052 151920 386104 151972
rect 399760 151920 399812 151972
rect 404636 151920 404688 151972
rect 423588 151920 423640 151972
rect 424968 151920 425020 151972
rect 436192 151988 436244 152040
rect 446956 151988 447008 152040
rect 447048 151988 447100 152040
rect 453764 151988 453816 152040
rect 456800 151988 456852 152040
rect 463332 151988 463384 152040
rect 467932 151988 467984 152040
rect 472348 151988 472400 152040
rect 487528 151988 487580 152040
rect 492220 151988 492272 152040
rect 499212 151988 499264 152040
rect 500592 151988 500644 152040
rect 385868 151852 385920 151904
rect 397184 151852 397236 151904
rect 397920 151852 397972 151904
rect 405556 151852 405608 151904
rect 405648 151852 405700 151904
rect 421012 151852 421064 151904
rect 334072 151784 334124 151836
rect 372160 151784 372212 151836
rect 380992 151784 381044 151836
rect 392124 151784 392176 151836
rect 397368 151784 397420 151836
rect 402980 151784 403032 151836
rect 419540 151784 419592 151836
rect 81716 151716 81768 151768
rect 112812 151716 112864 151768
rect 423496 151852 423548 151904
rect 439596 151920 439648 151972
rect 441712 151920 441764 151972
rect 446588 151920 446640 151972
rect 427084 151852 427136 151904
rect 437020 151852 437072 151904
rect 437480 151852 437532 151904
rect 445668 151852 445720 151904
rect 445760 151852 445812 151904
rect 448060 151920 448112 151972
rect 456984 151920 457036 151972
rect 468024 151920 468076 151972
rect 471704 151920 471756 151972
rect 487160 151920 487212 151972
rect 491576 151920 491628 151972
rect 498384 151920 498436 151972
rect 499948 151920 500000 151972
rect 516048 151920 516100 151972
rect 518992 151920 519044 151972
rect 460112 151852 460164 151904
rect 460204 151852 460256 151904
rect 462044 151852 462096 151904
rect 469220 151852 469272 151904
rect 472992 151852 473044 151904
rect 478880 151852 478932 151904
rect 480720 151852 480772 151904
rect 517428 151852 517480 151904
rect 520280 151852 520332 151904
rect 434444 151784 434496 151836
rect 441068 151784 441120 151836
rect 446588 151784 446640 151836
rect 446956 151784 447008 151836
rect 455052 151784 455104 151836
rect 466460 151784 466512 151836
rect 471060 151784 471112 151836
rect 485780 151784 485832 151836
rect 490288 151784 490340 151836
rect 98920 151648 98972 151700
rect 116032 151648 116084 151700
rect 95516 151580 95568 151632
rect 115296 151580 115348 151632
rect 92020 151512 92072 151564
rect 113088 151512 113140 151564
rect 26700 151444 26752 151496
rect 116952 151444 117004 151496
rect 16396 151376 16448 151428
rect 116768 151376 116820 151428
rect 12992 151308 13044 151360
rect 116676 151308 116728 151360
rect 68008 151240 68060 151292
rect 112720 151240 112772 151292
rect 64512 151172 64564 151224
rect 112628 151172 112680 151224
rect 61108 151104 61160 151156
rect 112536 151104 112588 151156
rect 57704 151036 57756 151088
rect 110972 151036 111024 151088
rect 54208 150968 54260 151020
rect 112444 150968 112496 151020
rect 50804 150900 50856 150952
rect 111708 150900 111760 150952
rect 47308 150832 47360 150884
rect 111616 150832 111668 150884
rect 43904 150764 43956 150816
rect 111524 150764 111576 150816
rect 40500 150696 40552 150748
rect 111432 150696 111484 150748
rect 37004 150628 37056 150680
rect 111248 150628 111300 150680
rect 88616 150560 88668 150612
rect 112996 150560 113048 150612
rect 85212 150492 85264 150544
rect 115204 150492 115256 150544
rect 102324 150424 102376 150476
rect 116124 150424 116176 150476
rect 78312 150288 78364 150340
rect 112904 150288 112956 150340
rect 109592 150220 109644 150272
rect 117228 150220 117280 150272
rect 108028 150152 108080 150204
rect 117044 150152 117096 150204
rect 145104 150152 145156 150204
rect 146254 150152 146306 150204
rect 146392 150152 146444 150204
rect 147542 150152 147594 150204
rect 163320 150152 163372 150204
rect 164194 150152 164246 150204
rect 164332 150152 164384 150204
rect 165482 150152 165534 150204
rect 171140 150152 171192 150204
rect 171922 150152 171974 150204
rect 181260 150152 181312 150204
rect 182134 150152 182186 150204
rect 182364 150152 182416 150204
rect 183422 150152 183474 150204
rect 183560 150152 183612 150204
rect 184710 150152 184762 150204
rect 200212 150152 200264 150204
rect 201454 150152 201506 150204
rect 213920 150152 213972 150204
rect 214886 150152 214938 150204
rect 218244 150152 218296 150204
rect 219394 150152 219446 150204
rect 238852 150152 238904 150204
rect 240002 150152 240054 150204
rect 242900 150152 242952 150204
rect 243774 150152 243826 150204
rect 247132 150152 247184 150204
rect 248282 150152 248334 150204
rect 251180 150152 251232 150204
rect 252146 150152 252198 150204
rect 256792 150152 256844 150204
rect 257942 150152 257994 150204
rect 258172 150152 258224 150204
rect 259230 150152 259282 150204
rect 260840 150152 260892 150204
rect 261806 150152 261858 150204
rect 271880 150152 271932 150204
rect 272754 150152 272806 150204
rect 311992 150152 312044 150204
rect 313142 150152 313194 150204
rect 328460 150152 328512 150204
rect 329242 150152 329294 150204
rect 332600 150152 332652 150204
rect 333750 150152 333802 150204
rect 339684 150152 339736 150204
rect 340742 150152 340794 150204
rect 349344 150152 349396 150204
rect 350402 150152 350454 150204
rect 357624 150152 357676 150204
rect 358774 150152 358826 150204
rect 358912 150152 358964 150204
rect 360062 150152 360114 150204
rect 363052 150152 363104 150204
rect 363926 150152 363978 150204
rect 368480 150152 368532 150204
rect 369630 150152 369682 150204
rect 403164 150152 403216 150204
rect 404314 150152 404366 150204
rect 446588 150152 446640 150204
rect 448014 150152 448066 150204
rect 465080 150152 465132 150204
rect 465954 150152 466006 150204
rect 477684 150152 477736 150204
rect 478834 150152 478886 150204
rect 483112 150152 483164 150204
rect 483986 150152 484038 150204
rect 505284 150152 505336 150204
rect 506434 150152 506486 150204
rect 506572 150152 506624 150204
rect 507722 150152 507774 150204
rect 507952 150152 508004 150204
rect 509010 150152 509062 150204
rect 509332 150152 509384 150204
rect 510298 150152 510350 150204
rect 518026 150152 518078 150204
rect 518808 150152 518860 150204
rect 82084 150084 82136 150136
rect 91008 150084 91060 150136
rect 116492 150084 116544 150136
rect 146576 150084 146628 150136
rect 150670 150084 150722 150136
rect 116400 150016 116452 150068
rect 111156 148316 111208 148368
rect 117136 148316 117188 148368
rect 113088 140700 113140 140752
rect 116124 140700 116176 140752
rect 112996 137912 113048 137964
rect 116124 137912 116176 137964
rect 116308 137300 116360 137352
rect 116492 137300 116544 137352
rect 112812 133832 112864 133884
rect 116032 133832 116084 133884
rect 114192 132608 114244 132660
rect 115204 132608 115256 132660
rect 112904 132404 112956 132456
rect 116124 132404 116176 132456
rect 112720 126896 112772 126948
rect 116032 126896 116084 126948
rect 112628 124108 112680 124160
rect 116124 124108 116176 124160
rect 112536 122748 112588 122800
rect 115940 122748 115992 122800
rect 111708 121388 111760 121440
rect 116124 121388 116176 121440
rect 112444 118600 112496 118652
rect 116124 118600 116176 118652
rect 116492 117988 116544 118040
rect 117228 117988 117280 118040
rect 111616 117240 111668 117292
rect 116124 117240 116176 117292
rect 111524 114452 111576 114504
rect 116124 114452 116176 114504
rect 111432 113092 111484 113144
rect 115940 113092 115992 113144
rect 111340 111732 111392 111784
rect 116124 111732 116176 111784
rect 111156 108944 111208 108996
rect 116124 108944 116176 108996
rect 111248 92420 111300 92472
rect 116124 92420 116176 92472
rect 111064 89632 111116 89684
rect 116124 89632 116176 89684
rect 113824 88272 113876 88324
rect 116032 88272 116084 88324
rect 113916 83920 113968 83972
rect 116584 83920 116636 83972
rect 114008 82764 114060 82816
rect 116216 82764 116268 82816
rect 114100 79976 114152 80028
rect 115940 79976 115992 80028
rect 114192 78616 114244 78668
rect 116124 78616 116176 78668
rect 114192 71748 114244 71800
rect 116584 71748 116636 71800
rect 114100 69028 114152 69080
rect 116308 69028 116360 69080
rect 114008 67600 114060 67652
rect 116124 67600 116176 67652
rect 113916 66240 113968 66292
rect 116584 66240 116636 66292
rect 113364 64676 113416 64728
rect 116584 64676 116636 64728
rect 113824 63520 113876 63572
rect 116216 63520 116268 63572
rect 112444 62092 112496 62144
rect 116124 62092 116176 62144
rect 112536 42780 112588 42832
rect 116124 42780 116176 42832
rect 115848 7896 115900 7948
rect 116768 7896 116820 7948
rect 117228 7828 117280 7880
rect 116952 7760 117004 7812
rect 117044 7760 117096 7812
rect 117320 7760 117372 7812
rect 116676 7692 116728 7744
rect 117044 7420 117096 7472
rect 111708 2864 111760 2916
rect 111800 2796 111852 2848
rect 170312 2456 170364 2508
rect 193588 2456 193640 2508
rect 294788 2456 294840 2508
rect 425796 2456 425848 2508
rect 443644 2456 443696 2508
rect 170312 2320 170364 2372
rect 62396 1844 62448 1896
rect 65340 1844 65392 1896
rect 68008 1844 68060 1896
rect 77116 1844 77168 1896
rect 77760 1844 77812 1896
rect 88340 1844 88392 1896
rect 89352 1844 89404 1896
rect 94872 1844 94924 1896
rect 100760 1844 100812 1896
rect 64144 1776 64196 1828
rect 69388 1776 69440 1828
rect 77024 1776 77076 1828
rect 85948 1776 86000 1828
rect 86040 1776 86092 1828
rect 111064 1912 111116 1964
rect 102692 1844 102744 1896
rect 104164 1844 104216 1896
rect 109224 1844 109276 1896
rect 109316 1844 109368 1896
rect 62672 1708 62724 1760
rect 68836 1708 68888 1760
rect 77944 1708 77996 1760
rect 78312 1708 78364 1760
rect 82636 1708 82688 1760
rect 100714 1708 100766 1760
rect 109592 1776 109644 1828
rect 109960 1708 110012 1760
rect 112444 1708 112496 1760
rect 69296 1640 69348 1692
rect 101036 1640 101088 1692
rect 59360 1572 59412 1624
rect 68560 1572 68612 1624
rect 79324 1572 79376 1624
rect 97264 1572 97316 1624
rect 99380 1572 99432 1624
rect 100714 1572 100766 1624
rect 100944 1572 100996 1624
rect 104164 1640 104216 1692
rect 106004 1640 106056 1692
rect 116584 1640 116636 1692
rect 101220 1572 101272 1624
rect 110144 1572 110196 1624
rect 72700 1504 72752 1556
rect 110420 1504 110472 1556
rect 42616 1436 42668 1488
rect 78128 1436 78180 1488
rect 97264 1436 97316 1488
rect 104164 1436 104216 1488
rect 104256 1436 104308 1488
rect 106280 1436 106332 1488
rect 106372 1436 106424 1488
rect 109316 1436 109368 1488
rect 109408 1436 109460 1488
rect 143632 1436 143684 1488
rect 46020 1368 46072 1420
rect 116492 1368 116544 1420
rect 294788 1368 294840 1420
rect 343640 1368 343692 1420
rect 491300 1368 491352 1420
rect 493600 1368 493652 1420
rect 2688 1300 2740 1352
rect 116308 1300 116360 1352
rect 39304 1232 39356 1284
rect 116400 1232 116452 1284
rect 49332 1164 49384 1216
rect 116676 1164 116728 1216
rect 52644 1096 52696 1148
rect 117228 1096 117280 1148
rect 55956 1028 56008 1080
rect 111800 1028 111852 1080
rect 65984 960 66036 1012
rect 116860 960 116912 1012
rect 76012 892 76064 944
rect 112536 892 112588 944
rect 98368 824 98420 876
rect 105084 824 105136 876
rect 92664 756 92716 808
rect 110052 756 110104 808
rect 103704 688 103756 740
rect 106372 688 106424 740
<< metal2 >>
rect 386 163200 442 164400
rect 492 163254 1164 163282
rect 400 158030 428 163200
rect 388 158024 440 158030
rect 388 157966 440 157972
rect 492 153950 520 163254
rect 1136 163146 1164 163254
rect 1214 163200 1270 164400
rect 2042 163200 2098 164400
rect 2870 163200 2926 164400
rect 2976 163254 3648 163282
rect 1228 163146 1256 163200
rect 1136 163118 1256 163146
rect 2056 156670 2084 163200
rect 2884 159390 2912 163200
rect 2872 159384 2924 159390
rect 2872 159326 2924 159332
rect 2044 156664 2096 156670
rect 2044 156606 2096 156612
rect 480 153944 532 153950
rect 480 153886 532 153892
rect 2976 153882 3004 163254
rect 3620 163146 3648 163254
rect 3698 163200 3754 164400
rect 4526 163200 4582 164400
rect 5354 163200 5410 164400
rect 5552 163254 6132 163282
rect 3712 163146 3740 163200
rect 3620 163118 3740 163146
rect 4540 155378 4568 163200
rect 4528 155372 4580 155378
rect 4528 155314 4580 155320
rect 5368 155242 5396 163200
rect 5356 155236 5408 155242
rect 5356 155178 5408 155184
rect 2964 153876 3016 153882
rect 2964 153818 3016 153824
rect 5552 152425 5580 163254
rect 6104 163146 6132 163254
rect 6182 163200 6238 164400
rect 7102 163200 7158 164400
rect 7576 163254 7880 163282
rect 6196 163146 6224 163200
rect 6104 163118 6224 163146
rect 7116 153785 7144 163200
rect 7576 153921 7604 163254
rect 7852 163146 7880 163254
rect 7930 163200 7986 164400
rect 8758 163200 8814 164400
rect 9586 163200 9642 164400
rect 9692 163254 10364 163282
rect 7944 163146 7972 163200
rect 7852 163118 7972 163146
rect 8772 155310 8800 163200
rect 9600 159497 9628 163200
rect 9586 159488 9642 159497
rect 9586 159423 9642 159432
rect 8760 155304 8812 155310
rect 8760 155246 8812 155252
rect 9692 154057 9720 163254
rect 10336 163146 10364 163254
rect 10414 163200 10470 164400
rect 11242 163200 11298 164400
rect 12070 163200 12126 164400
rect 12452 163254 12848 163282
rect 10428 163146 10456 163200
rect 10336 163118 10456 163146
rect 11256 155990 11284 163200
rect 12084 156466 12112 163200
rect 12072 156460 12124 156466
rect 12072 156402 12124 156408
rect 11244 155984 11296 155990
rect 11244 155926 11296 155932
rect 9678 154048 9734 154057
rect 9678 153983 9734 153992
rect 7562 153912 7618 153921
rect 7562 153847 7618 153856
rect 7102 153776 7158 153785
rect 7102 153711 7158 153720
rect 9496 152992 9548 152998
rect 9496 152934 9548 152940
rect 5538 152416 5594 152425
rect 5538 152351 5594 152360
rect 6090 150648 6146 150657
rect 6090 150583 6146 150592
rect 2686 150512 2742 150521
rect 2686 150447 2742 150456
rect 2700 149940 2728 150447
rect 6104 149940 6132 150583
rect 9508 149940 9536 152934
rect 12452 152522 12480 163254
rect 12820 163146 12848 163254
rect 12898 163200 12954 164400
rect 13818 163200 13874 164400
rect 14646 163200 14702 164400
rect 15474 163200 15530 164400
rect 16302 163200 16358 164400
rect 16592 163254 17080 163282
rect 12912 163146 12940 163200
rect 12820 163118 12940 163146
rect 13832 154086 13860 163200
rect 14660 156738 14688 163200
rect 14648 156732 14700 156738
rect 14648 156674 14700 156680
rect 15488 156262 15516 163200
rect 16316 159361 16344 163200
rect 16302 159352 16358 159361
rect 16302 159287 16358 159296
rect 15476 156256 15528 156262
rect 15476 156198 15528 156204
rect 13820 154080 13872 154086
rect 13820 154022 13872 154028
rect 16592 154018 16620 163254
rect 17052 163146 17080 163254
rect 17130 163200 17186 164400
rect 17958 163200 18014 164400
rect 18064 163254 18736 163282
rect 17144 163146 17172 163200
rect 17052 163118 17172 163146
rect 17972 156942 18000 163200
rect 17960 156936 18012 156942
rect 17960 156878 18012 156884
rect 16580 154012 16632 154018
rect 16580 153954 16632 153960
rect 18064 152590 18092 163254
rect 18708 163146 18736 163254
rect 18786 163200 18842 164400
rect 19352 163254 19564 163282
rect 18800 163146 18828 163200
rect 18708 163118 18828 163146
rect 18052 152584 18104 152590
rect 19352 152561 19380 163254
rect 19536 163146 19564 163254
rect 19614 163200 19670 164400
rect 19720 163254 20484 163282
rect 19628 163146 19656 163200
rect 19536 163118 19656 163146
rect 19720 154193 19748 163254
rect 20456 163146 20484 163254
rect 20534 163200 20590 164400
rect 21362 163200 21418 164400
rect 22190 163200 22246 164400
rect 23018 163200 23074 164400
rect 23492 163254 23796 163282
rect 20548 163146 20576 163200
rect 20456 163118 20576 163146
rect 21376 156874 21404 163200
rect 22204 159594 22232 163200
rect 22192 159588 22244 159594
rect 22192 159530 22244 159536
rect 23032 159458 23060 163200
rect 23020 159452 23072 159458
rect 23020 159394 23072 159400
rect 21364 156868 21416 156874
rect 21364 156810 21416 156816
rect 19706 154184 19762 154193
rect 23492 154154 23520 163254
rect 23768 163146 23796 163254
rect 23846 163200 23902 164400
rect 24674 163200 24730 164400
rect 24872 163254 25452 163282
rect 23860 163146 23888 163200
rect 23768 163118 23888 163146
rect 24688 157010 24716 163200
rect 24676 157004 24728 157010
rect 24676 156946 24728 156952
rect 19706 154119 19762 154128
rect 23480 154148 23532 154154
rect 23480 154090 23532 154096
rect 23296 153060 23348 153066
rect 23296 153002 23348 153008
rect 18052 152526 18104 152532
rect 19338 152552 19394 152561
rect 12440 152516 12492 152522
rect 19338 152487 19394 152496
rect 12440 152458 12492 152464
rect 19800 152108 19852 152114
rect 19800 152050 19852 152056
rect 16396 151428 16448 151434
rect 16396 151370 16448 151376
rect 12992 151360 13044 151366
rect 12992 151302 13044 151308
rect 13004 149940 13032 151302
rect 16408 149940 16436 151370
rect 19812 149940 19840 152050
rect 23308 149940 23336 153002
rect 24872 152697 24900 163254
rect 25424 163146 25452 163254
rect 25502 163200 25558 164400
rect 26330 163200 26386 164400
rect 26896 163254 27200 163282
rect 25516 163146 25544 163200
rect 25424 163118 25544 163146
rect 26344 152794 26372 163200
rect 26896 154222 26924 163254
rect 27172 163146 27200 163254
rect 27250 163200 27306 164400
rect 28078 163200 28134 164400
rect 28906 163200 28962 164400
rect 29734 163200 29790 164400
rect 30562 163200 30618 164400
rect 31390 163200 31446 164400
rect 31772 163254 32168 163282
rect 27264 163146 27292 163200
rect 27172 163118 27292 163146
rect 28092 157078 28120 163200
rect 28920 159526 28948 163200
rect 29748 159633 29776 163200
rect 29734 159624 29790 159633
rect 29734 159559 29790 159568
rect 28908 159520 28960 159526
rect 28908 159462 28960 159468
rect 28080 157072 28132 157078
rect 28080 157014 28132 157020
rect 30576 154290 30604 163200
rect 31404 157146 31432 163200
rect 31392 157140 31444 157146
rect 31392 157082 31444 157088
rect 30564 154284 30616 154290
rect 30564 154226 30616 154232
rect 26884 154216 26936 154222
rect 26884 154158 26936 154164
rect 30196 153128 30248 153134
rect 30196 153070 30248 153076
rect 26332 152788 26384 152794
rect 26332 152730 26384 152736
rect 24858 152688 24914 152697
rect 24858 152623 24914 152632
rect 26700 151496 26752 151502
rect 26700 151438 26752 151444
rect 26712 149940 26740 151438
rect 30208 149940 30236 153070
rect 31772 152658 31800 163254
rect 32140 163146 32168 163254
rect 32218 163200 32274 164400
rect 33138 163200 33194 164400
rect 33966 163200 34022 164400
rect 34532 163254 34744 163282
rect 32232 163146 32260 163200
rect 32140 163118 32260 163146
rect 33152 152862 33180 163200
rect 33980 158001 34008 163200
rect 33966 157992 34022 158001
rect 33966 157927 34022 157936
rect 34532 153270 34560 163254
rect 34716 163146 34744 163254
rect 34794 163200 34850 164400
rect 35622 163200 35678 164400
rect 36450 163200 36506 164400
rect 37278 163200 37334 164400
rect 37384 163254 38056 163282
rect 34808 163146 34836 163200
rect 34716 163118 34836 163146
rect 35636 156641 35664 163200
rect 35622 156632 35678 156641
rect 35622 156567 35678 156576
rect 36464 155650 36492 163200
rect 37292 158098 37320 163200
rect 37280 158092 37332 158098
rect 37280 158034 37332 158040
rect 36452 155644 36504 155650
rect 36452 155586 36504 155592
rect 37384 154329 37412 163254
rect 38028 163146 38056 163254
rect 38106 163200 38162 164400
rect 38934 163200 38990 164400
rect 39854 163200 39910 164400
rect 40682 163200 40738 164400
rect 41510 163200 41566 164400
rect 42338 163200 42394 164400
rect 43166 163200 43222 164400
rect 43994 163200 44050 164400
rect 44192 163254 44772 163282
rect 38120 163146 38148 163200
rect 38028 163118 38148 163146
rect 38948 157214 38976 163200
rect 39868 159662 39896 163200
rect 39856 159656 39908 159662
rect 39856 159598 39908 159604
rect 40696 158137 40724 163200
rect 40682 158128 40738 158137
rect 40682 158063 40738 158072
rect 38936 157208 38988 157214
rect 38936 157150 38988 157156
rect 41524 154426 41552 163200
rect 42352 156777 42380 163200
rect 42338 156768 42394 156777
rect 42338 156703 42394 156712
rect 43180 155786 43208 163200
rect 44008 158273 44036 163200
rect 43994 158264 44050 158273
rect 43994 158199 44050 158208
rect 43168 155780 43220 155786
rect 43168 155722 43220 155728
rect 44192 154494 44220 163254
rect 44744 163146 44772 163254
rect 44822 163200 44878 164400
rect 45650 163200 45706 164400
rect 46570 163200 46626 164400
rect 47398 163200 47454 164400
rect 48226 163200 48282 164400
rect 49054 163200 49110 164400
rect 49882 163200 49938 164400
rect 50710 163200 50766 164400
rect 51538 163200 51594 164400
rect 52366 163200 52422 164400
rect 53286 163200 53342 164400
rect 54114 163200 54170 164400
rect 54942 163200 54998 164400
rect 55770 163200 55826 164400
rect 56598 163200 56654 164400
rect 57426 163200 57482 164400
rect 58254 163200 58310 164400
rect 58360 163254 59032 163282
rect 44836 163146 44864 163200
rect 44744 163118 44864 163146
rect 45664 157350 45692 163200
rect 45652 157344 45704 157350
rect 45652 157286 45704 157292
rect 46584 155718 46612 163200
rect 47412 158234 47440 163200
rect 47400 158228 47452 158234
rect 47400 158170 47452 158176
rect 46572 155712 46624 155718
rect 46572 155654 46624 155660
rect 48240 155446 48268 163200
rect 49068 157282 49096 163200
rect 49896 159934 49924 163200
rect 49884 159928 49936 159934
rect 49884 159870 49936 159876
rect 50724 158166 50752 163200
rect 50712 158160 50764 158166
rect 50712 158102 50764 158108
rect 49056 157276 49108 157282
rect 49056 157218 49108 157224
rect 51552 155582 51580 163200
rect 52380 156913 52408 163200
rect 53300 159730 53328 163200
rect 53288 159724 53340 159730
rect 53288 159666 53340 159672
rect 54128 158302 54156 163200
rect 54116 158296 54168 158302
rect 54116 158238 54168 158244
rect 52366 156904 52422 156913
rect 52366 156839 52422 156848
rect 51540 155576 51592 155582
rect 51540 155518 51592 155524
rect 54956 155514 54984 163200
rect 55784 157049 55812 163200
rect 55770 157040 55826 157049
rect 55770 156975 55826 156984
rect 54944 155508 54996 155514
rect 54944 155450 54996 155456
rect 48228 155440 48280 155446
rect 48228 155382 48280 155388
rect 56612 155174 56640 163200
rect 57440 158409 57468 163200
rect 57426 158400 57482 158409
rect 57426 158335 57482 158344
rect 58268 155417 58296 163200
rect 58254 155408 58310 155417
rect 58254 155343 58310 155352
rect 56600 155168 56652 155174
rect 56600 155110 56652 155116
rect 58360 154562 58388 163254
rect 59004 163146 59032 163254
rect 59082 163200 59138 164400
rect 60002 163200 60058 164400
rect 60830 163200 60886 164400
rect 61658 163200 61714 164400
rect 62132 163254 62436 163282
rect 59096 163146 59124 163200
rect 59004 163118 59124 163146
rect 60016 159798 60044 163200
rect 60004 159792 60056 159798
rect 60004 159734 60056 159740
rect 60844 158506 60872 163200
rect 60832 158500 60884 158506
rect 60832 158442 60884 158448
rect 61672 155281 61700 163200
rect 61658 155272 61714 155281
rect 61658 155207 61714 155216
rect 58348 154556 58400 154562
rect 58348 154498 58400 154504
rect 44180 154488 44232 154494
rect 44180 154430 44232 154436
rect 41512 154420 41564 154426
rect 41512 154362 41564 154368
rect 37370 154320 37426 154329
rect 37370 154255 37426 154264
rect 62132 153814 62160 163254
rect 62408 163146 62436 163254
rect 62486 163200 62542 164400
rect 63314 163200 63370 164400
rect 64142 163200 64198 164400
rect 64970 163200 65026 164400
rect 65168 163254 65840 163282
rect 62500 163146 62528 163200
rect 62408 163118 62528 163146
rect 63328 159186 63356 163200
rect 63316 159180 63368 159186
rect 63316 159122 63368 159128
rect 64156 158438 64184 163200
rect 64144 158432 64196 158438
rect 64144 158374 64196 158380
rect 64984 155650 65012 163200
rect 63500 155644 63552 155650
rect 63500 155586 63552 155592
rect 64972 155644 65024 155650
rect 64972 155586 65024 155592
rect 62120 153808 62172 153814
rect 62120 153750 62172 153756
rect 34520 153264 34572 153270
rect 34520 153206 34572 153212
rect 33140 152856 33192 152862
rect 33140 152798 33192 152804
rect 31760 152652 31812 152658
rect 31760 152594 31812 152600
rect 33600 152244 33652 152250
rect 33600 152186 33652 152192
rect 33612 149940 33640 152186
rect 63512 152046 63540 155586
rect 65168 154465 65196 163254
rect 65812 163146 65840 163254
rect 65890 163200 65946 164400
rect 66718 163200 66774 164400
rect 67546 163200 67602 164400
rect 68374 163200 68430 164400
rect 69202 163200 69258 164400
rect 70030 163200 70086 164400
rect 70858 163200 70914 164400
rect 71686 163200 71742 164400
rect 71792 163254 72556 163282
rect 65904 163146 65932 163200
rect 65812 163118 65932 163146
rect 66732 160070 66760 163200
rect 66720 160064 66772 160070
rect 66720 160006 66772 160012
rect 67560 158370 67588 163200
rect 67548 158364 67600 158370
rect 67548 158306 67600 158312
rect 68388 155553 68416 163200
rect 69216 156602 69244 163200
rect 70044 159866 70072 163200
rect 70032 159860 70084 159866
rect 70032 159802 70084 159808
rect 70872 158642 70900 163200
rect 70860 158636 70912 158642
rect 70860 158578 70912 158584
rect 69204 156596 69256 156602
rect 69204 156538 69256 156544
rect 71700 155718 71728 163200
rect 69664 155712 69716 155718
rect 69664 155654 69716 155660
rect 71688 155712 71740 155718
rect 71688 155654 71740 155660
rect 68374 155544 68430 155553
rect 68374 155479 68430 155488
rect 65154 154456 65210 154465
rect 65154 154391 65210 154400
rect 69676 152182 69704 155654
rect 71792 153746 71820 163254
rect 72528 163146 72556 163254
rect 72606 163200 72662 164400
rect 73434 163200 73490 164400
rect 74262 163200 74318 164400
rect 75090 163200 75146 164400
rect 75918 163200 75974 164400
rect 76746 163200 76802 164400
rect 77574 163200 77630 164400
rect 78402 163200 78458 164400
rect 79322 163200 79378 164400
rect 80150 163200 80206 164400
rect 80978 163200 81034 164400
rect 81806 163200 81862 164400
rect 81912 163254 82584 163282
rect 72620 163146 72648 163200
rect 72528 163118 72648 163146
rect 73448 155106 73476 163200
rect 74276 158574 74304 163200
rect 74264 158568 74316 158574
rect 74264 158510 74316 158516
rect 75104 155854 75132 163200
rect 75932 155922 75960 163200
rect 76760 160002 76788 163200
rect 76748 159996 76800 160002
rect 76748 159938 76800 159944
rect 77588 157962 77616 163200
rect 77576 157956 77628 157962
rect 77576 157898 77628 157904
rect 75920 155916 75972 155922
rect 75920 155858 75972 155864
rect 75092 155848 75144 155854
rect 75092 155790 75144 155796
rect 78416 155786 78444 163200
rect 79336 156534 79364 163200
rect 80164 159118 80192 163200
rect 80152 159112 80204 159118
rect 80152 159054 80204 159060
rect 80992 158710 81020 163200
rect 80980 158704 81032 158710
rect 80980 158646 81032 158652
rect 79324 156528 79376 156534
rect 79324 156470 79376 156476
rect 75828 155780 75880 155786
rect 75828 155722 75880 155728
rect 78404 155780 78456 155786
rect 78404 155722 78456 155728
rect 73436 155100 73488 155106
rect 73436 155042 73488 155048
rect 71780 153740 71832 153746
rect 71780 153682 71832 153688
rect 69664 152176 69716 152182
rect 69664 152118 69716 152124
rect 63500 152040 63552 152046
rect 63500 151982 63552 151988
rect 75840 151978 75868 155722
rect 81820 155174 81848 163200
rect 76472 155168 76524 155174
rect 76472 155110 76524 155116
rect 81808 155168 81860 155174
rect 81808 155110 81860 155116
rect 76484 152318 76512 155110
rect 81440 155100 81492 155106
rect 81440 155042 81492 155048
rect 81452 152454 81480 155042
rect 81912 153678 81940 163254
rect 82556 163146 82584 163254
rect 82634 163200 82690 164400
rect 83462 163200 83518 164400
rect 84290 163200 84346 164400
rect 85118 163200 85174 164400
rect 86038 163200 86094 164400
rect 86144 163254 86816 163282
rect 82648 163146 82676 163200
rect 82556 163118 82676 163146
rect 83476 159322 83504 163200
rect 83464 159316 83516 159322
rect 83464 159258 83516 159264
rect 84304 157758 84332 163200
rect 84292 157752 84344 157758
rect 84292 157694 84344 157700
rect 85132 155689 85160 163200
rect 85118 155680 85174 155689
rect 85118 155615 85174 155624
rect 86052 154970 86080 163200
rect 86040 154964 86092 154970
rect 86040 154906 86092 154912
rect 81900 153672 81952 153678
rect 81900 153614 81952 153620
rect 86144 152726 86172 163254
rect 86788 163146 86816 163254
rect 86866 163200 86922 164400
rect 87694 163200 87750 164400
rect 88522 163200 88578 164400
rect 89350 163200 89406 164400
rect 90178 163200 90234 164400
rect 91006 163200 91062 164400
rect 91834 163200 91890 164400
rect 92754 163200 92810 164400
rect 93320 163254 93532 163282
rect 86880 163146 86908 163200
rect 86788 163118 86908 163146
rect 87708 157894 87736 163200
rect 87696 157888 87748 157894
rect 87696 157830 87748 157836
rect 88536 155106 88564 163200
rect 89364 156398 89392 163200
rect 90192 159254 90220 163200
rect 90180 159248 90232 159254
rect 90180 159190 90232 159196
rect 89720 159112 89772 159118
rect 89720 159054 89772 159060
rect 89352 156392 89404 156398
rect 89352 156334 89404 156340
rect 88524 155100 88576 155106
rect 88524 155042 88576 155048
rect 86132 152720 86184 152726
rect 86132 152662 86184 152668
rect 81440 152448 81492 152454
rect 81440 152390 81492 152396
rect 89732 152386 89760 159054
rect 91020 157826 91048 163200
rect 91008 157820 91060 157826
rect 91008 157762 91060 157768
rect 91848 155038 91876 163200
rect 92768 159050 92796 163200
rect 92756 159044 92808 159050
rect 92756 158986 92808 158992
rect 91836 155032 91888 155038
rect 91836 154974 91888 154980
rect 92572 152992 92624 152998
rect 92572 152934 92624 152940
rect 89720 152380 89772 152386
rect 89720 152322 89772 152328
rect 76472 152312 76524 152318
rect 76472 152254 76524 152260
rect 75828 151972 75880 151978
rect 75828 151914 75880 151920
rect 74816 151904 74868 151910
rect 74816 151846 74868 151852
rect 82084 151904 82136 151910
rect 82084 151846 82136 151852
rect 71412 151836 71464 151842
rect 71412 151778 71464 151784
rect 68008 151292 68060 151298
rect 68008 151234 68060 151240
rect 64512 151224 64564 151230
rect 64512 151166 64564 151172
rect 61108 151156 61160 151162
rect 61108 151098 61160 151104
rect 57704 151088 57756 151094
rect 57704 151030 57756 151036
rect 54208 151020 54260 151026
rect 54208 150962 54260 150968
rect 50804 150952 50856 150958
rect 50804 150894 50856 150900
rect 47308 150884 47360 150890
rect 47308 150826 47360 150832
rect 43904 150816 43956 150822
rect 43904 150758 43956 150764
rect 40500 150748 40552 150754
rect 40500 150690 40552 150696
rect 37004 150680 37056 150686
rect 37004 150622 37056 150628
rect 37016 149940 37044 150622
rect 40512 149940 40540 150690
rect 43916 149940 43944 150758
rect 47320 149940 47348 150826
rect 50816 149940 50844 150894
rect 54220 149940 54248 150962
rect 57716 149940 57744 151030
rect 61120 149940 61148 151098
rect 64524 149940 64552 151166
rect 68020 149940 68048 151234
rect 71424 149940 71452 151778
rect 74828 149940 74856 151846
rect 81716 151768 81768 151774
rect 81716 151710 81768 151716
rect 78312 150340 78364 150346
rect 78312 150282 78364 150288
rect 78324 149940 78352 150282
rect 81728 149940 81756 151710
rect 82096 150142 82124 151846
rect 91008 151836 91060 151842
rect 91008 151778 91060 151784
rect 88616 150612 88668 150618
rect 88616 150554 88668 150560
rect 85212 150544 85264 150550
rect 85212 150486 85264 150492
rect 82084 150136 82136 150142
rect 82084 150078 82136 150084
rect 85224 149940 85252 150486
rect 88628 149940 88656 150554
rect 91020 150142 91048 151778
rect 92020 151564 92072 151570
rect 92020 151506 92072 151512
rect 91008 150136 91060 150142
rect 91008 150078 91060 150084
rect 92032 149940 92060 151506
rect 92584 149705 92612 152934
rect 93320 152930 93348 163254
rect 93504 163146 93532 163254
rect 93582 163200 93638 164400
rect 94410 163200 94466 164400
rect 95238 163200 95294 164400
rect 96066 163200 96122 164400
rect 96894 163200 96950 164400
rect 97722 163200 97778 164400
rect 98642 163200 98698 164400
rect 99470 163200 99526 164400
rect 99576 163254 100248 163282
rect 93596 163146 93624 163200
rect 93504 163118 93624 163146
rect 94424 157690 94452 163200
rect 94412 157684 94464 157690
rect 94412 157626 94464 157632
rect 95252 154766 95280 163200
rect 96080 154902 96108 163200
rect 96908 159118 96936 163200
rect 96896 159112 96948 159118
rect 96896 159054 96948 159060
rect 97736 156330 97764 163200
rect 97724 156324 97776 156330
rect 97724 156266 97776 156272
rect 96068 154896 96120 154902
rect 96068 154838 96120 154844
rect 98656 154834 98684 163200
rect 99484 158778 99512 163200
rect 99472 158772 99524 158778
rect 99472 158714 99524 158720
rect 98644 154828 98696 154834
rect 98644 154770 98696 154776
rect 95240 154760 95292 154766
rect 95240 154702 95292 154708
rect 99576 152998 99604 163254
rect 100220 163146 100248 163254
rect 100298 163200 100354 164400
rect 101126 163200 101182 164400
rect 101324 163254 101904 163282
rect 100312 163146 100340 163200
rect 100220 163118 100340 163146
rect 101140 158545 101168 163200
rect 101126 158536 101182 158545
rect 101126 158471 101182 158480
rect 101324 153610 101352 163254
rect 101876 163146 101904 163254
rect 101954 163200 102010 164400
rect 102782 163200 102838 164400
rect 103610 163200 103666 164400
rect 104438 163200 104494 164400
rect 104912 163254 105308 163282
rect 101968 163146 101996 163200
rect 101876 163118 101996 163146
rect 102140 159180 102192 159186
rect 102140 159122 102192 159128
rect 101312 153604 101364 153610
rect 101312 153546 101364 153552
rect 99564 152992 99616 152998
rect 99564 152934 99616 152940
rect 93308 152924 93360 152930
rect 93308 152866 93360 152872
rect 99932 152108 99984 152114
rect 99932 152050 99984 152056
rect 98920 151700 98972 151706
rect 98920 151642 98972 151648
rect 95516 151632 95568 151638
rect 95516 151574 95568 151580
rect 95528 149940 95556 151574
rect 98932 149940 98960 151642
rect 99944 149841 99972 152050
rect 102152 151842 102180 159122
rect 102796 158846 102824 163200
rect 103624 159186 103652 163200
rect 103612 159180 103664 159186
rect 103612 159122 103664 159128
rect 102784 158840 102836 158846
rect 102784 158782 102836 158788
rect 104452 157185 104480 163200
rect 104438 157176 104494 157185
rect 104438 157111 104494 157120
rect 104912 153542 104940 163254
rect 105280 163146 105308 163254
rect 105358 163200 105414 164400
rect 106186 163200 106242 164400
rect 107014 163200 107070 164400
rect 107842 163200 107898 164400
rect 107948 163254 108620 163282
rect 105372 163146 105400 163200
rect 105280 163118 105400 163146
rect 106200 158914 106228 163200
rect 106188 158908 106240 158914
rect 106188 158850 106240 158856
rect 107028 157418 107056 163200
rect 107856 157554 107884 163200
rect 107844 157548 107896 157554
rect 107844 157490 107896 157496
rect 107016 157412 107068 157418
rect 107016 157354 107068 157360
rect 107752 157412 107804 157418
rect 107752 157354 107804 157360
rect 104900 153536 104952 153542
rect 104900 153478 104952 153484
rect 107764 153202 107792 157354
rect 107948 153474 107976 163254
rect 108592 163146 108620 163254
rect 108670 163200 108726 164400
rect 109498 163200 109554 164400
rect 110326 163200 110382 164400
rect 111154 163200 111210 164400
rect 111812 163254 112024 163282
rect 108684 163146 108712 163200
rect 108592 163118 108712 163146
rect 109040 156460 109092 156466
rect 109040 156402 109092 156408
rect 107936 153468 107988 153474
rect 107936 153410 107988 153416
rect 107752 153196 107804 153202
rect 107752 153138 107804 153144
rect 108028 153060 108080 153066
rect 108028 153002 108080 153008
rect 105820 151972 105872 151978
rect 105820 151914 105872 151920
rect 102140 151836 102192 151842
rect 102140 151778 102192 151784
rect 102324 150476 102376 150482
rect 102324 150418 102376 150424
rect 102336 149940 102364 150418
rect 105832 149940 105860 151914
rect 108040 150210 108068 153002
rect 109052 152114 109080 156402
rect 109512 156194 109540 163200
rect 109684 156256 109736 156262
rect 109684 156198 109736 156204
rect 109500 156188 109552 156194
rect 109500 156130 109552 156136
rect 109696 152250 109724 156198
rect 110340 153066 110368 163200
rect 111168 157622 111196 163200
rect 111156 157616 111208 157622
rect 111156 157558 111208 157564
rect 111812 153406 111840 163254
rect 111996 163146 112024 163254
rect 112074 163200 112130 164400
rect 112272 163254 112852 163282
rect 112088 163146 112116 163200
rect 111996 163118 112116 163146
rect 111800 153400 111852 153406
rect 111800 153342 111852 153348
rect 112272 153338 112300 163254
rect 112824 163146 112852 163254
rect 112902 163200 112958 164400
rect 113730 163200 113786 164400
rect 114558 163200 114614 164400
rect 115386 163200 115442 164400
rect 116214 163200 116270 164400
rect 116412 163254 116992 163282
rect 112916 163146 112944 163200
rect 112824 163118 112944 163146
rect 113640 158976 113692 158982
rect 113640 158918 113692 158924
rect 113652 158778 113680 158918
rect 113744 158778 113772 163200
rect 113640 158772 113692 158778
rect 113640 158714 113692 158720
rect 113732 158772 113784 158778
rect 113732 158714 113784 158720
rect 114572 156262 114600 163200
rect 115400 156466 115428 163200
rect 116228 159390 116256 163200
rect 116124 159384 116176 159390
rect 116124 159326 116176 159332
rect 116216 159384 116268 159390
rect 116216 159326 116268 159332
rect 116136 159050 116164 159326
rect 116032 159044 116084 159050
rect 116032 158986 116084 158992
rect 116124 159044 116176 159050
rect 116124 158986 116176 158992
rect 115388 156460 115440 156466
rect 115388 156402 115440 156408
rect 114560 156256 114612 156262
rect 114560 156198 114612 156204
rect 116044 154358 116072 158986
rect 116032 154352 116084 154358
rect 116032 154294 116084 154300
rect 112260 153332 112312 153338
rect 112260 153274 112312 153280
rect 116412 153134 116440 163254
rect 116964 163146 116992 163254
rect 117042 163200 117098 164400
rect 117870 163200 117926 164400
rect 118790 163200 118846 164400
rect 119618 163200 119674 164400
rect 120446 163200 120502 164400
rect 121274 163200 121330 164400
rect 122102 163200 122158 164400
rect 122930 163200 122986 164400
rect 123758 163200 123814 164400
rect 124586 163200 124642 164400
rect 125506 163200 125562 164400
rect 126334 163200 126390 164400
rect 127162 163200 127218 164400
rect 127990 163200 128046 164400
rect 128818 163200 128874 164400
rect 129646 163200 129702 164400
rect 129752 163254 130424 163282
rect 117056 163146 117084 163200
rect 116964 163118 117084 163146
rect 117884 157486 117912 163200
rect 118700 159044 118752 159050
rect 118700 158986 118752 158992
rect 117872 157480 117924 157486
rect 117872 157422 117924 157428
rect 110972 153128 111024 153134
rect 110972 153070 111024 153076
rect 116400 153128 116452 153134
rect 118712 153105 118740 158986
rect 118804 154698 118832 163200
rect 119632 159050 119660 163200
rect 119620 159044 119672 159050
rect 119620 158986 119672 158992
rect 120460 158982 120488 163200
rect 120080 158976 120132 158982
rect 120080 158918 120132 158924
rect 120448 158976 120500 158982
rect 120448 158918 120500 158924
rect 118884 158024 118936 158030
rect 118884 157966 118936 157972
rect 118792 154692 118844 154698
rect 118792 154634 118844 154640
rect 116400 153070 116452 153076
rect 118698 153096 118754 153105
rect 110328 153060 110380 153066
rect 110328 153002 110380 153008
rect 109592 152244 109644 152250
rect 109592 152186 109644 152192
rect 109684 152244 109736 152250
rect 109684 152186 109736 152192
rect 109040 152108 109092 152114
rect 109040 152050 109092 152056
rect 109604 150278 109632 152186
rect 110328 151972 110380 151978
rect 110328 151914 110380 151920
rect 109592 150272 109644 150278
rect 109592 150214 109644 150220
rect 108028 150204 108080 150210
rect 108028 150146 108080 150152
rect 99930 149832 99986 149841
rect 99930 149767 99986 149776
rect 92570 149696 92626 149705
rect 92570 149631 92626 149640
rect 109250 149382 109632 149410
rect 109604 148073 109632 149382
rect 109590 148064 109646 148073
rect 109590 147999 109646 148008
rect 110340 146441 110368 151914
rect 110984 151814 111012 153070
rect 118698 153031 118754 153040
rect 110984 151786 111196 151814
rect 110972 151088 111024 151094
rect 110972 151030 111024 151036
rect 110984 147393 111012 151030
rect 111062 150512 111118 150521
rect 111062 150447 111118 150456
rect 110970 147384 111026 147393
rect 110970 147319 111026 147328
rect 110326 146432 110382 146441
rect 110326 146367 110382 146376
rect 111076 89690 111104 150447
rect 111168 148374 111196 151786
rect 112812 151768 112864 151774
rect 112812 151710 112864 151716
rect 112720 151292 112772 151298
rect 112720 151234 112772 151240
rect 112628 151224 112680 151230
rect 112628 151166 112680 151172
rect 112536 151156 112588 151162
rect 112536 151098 112588 151104
rect 112444 151020 112496 151026
rect 112444 150962 112496 150968
rect 111708 150952 111760 150958
rect 111708 150894 111760 150900
rect 111616 150884 111668 150890
rect 111616 150826 111668 150832
rect 111524 150816 111576 150822
rect 111524 150758 111576 150764
rect 111432 150748 111484 150754
rect 111432 150690 111484 150696
rect 111248 150680 111300 150686
rect 111248 150622 111300 150628
rect 111338 150648 111394 150657
rect 111156 148368 111208 148374
rect 111156 148310 111208 148316
rect 111260 148186 111288 150622
rect 111338 150583 111394 150592
rect 111168 148158 111288 148186
rect 111168 109002 111196 148158
rect 111352 148050 111380 150583
rect 111260 148022 111380 148050
rect 111156 108996 111208 109002
rect 111156 108938 111208 108944
rect 111260 92478 111288 148022
rect 111444 147914 111472 150690
rect 111352 147886 111472 147914
rect 111352 111790 111380 147886
rect 111536 147778 111564 150758
rect 111444 147750 111564 147778
rect 111444 113150 111472 147750
rect 111628 147642 111656 150826
rect 111536 147614 111656 147642
rect 111536 114510 111564 147614
rect 111720 147506 111748 150894
rect 111628 147478 111748 147506
rect 111628 117298 111656 147478
rect 111706 147384 111762 147393
rect 111706 147319 111762 147328
rect 111720 121446 111748 147319
rect 111708 121440 111760 121446
rect 111708 121382 111760 121388
rect 112456 118658 112484 150962
rect 112548 122806 112576 151098
rect 112640 124166 112668 151166
rect 112732 126954 112760 151234
rect 112824 133890 112852 151710
rect 116032 151700 116084 151706
rect 116032 151642 116084 151648
rect 115296 151632 115348 151638
rect 115296 151574 115348 151580
rect 113088 151564 113140 151570
rect 113088 151506 113140 151512
rect 112996 150612 113048 150618
rect 112996 150554 113048 150560
rect 112904 150340 112956 150346
rect 112904 150282 112956 150288
rect 112812 133884 112864 133890
rect 112812 133826 112864 133832
rect 112916 132462 112944 150282
rect 113008 137970 113036 150554
rect 113100 140758 113128 151506
rect 115204 150544 115256 150550
rect 115204 150486 115256 150492
rect 113822 144256 113878 144265
rect 113822 144191 113878 144200
rect 113088 140752 113140 140758
rect 113088 140694 113140 140700
rect 112996 137964 113048 137970
rect 112996 137906 113048 137912
rect 112904 132456 112956 132462
rect 112904 132398 112956 132404
rect 112720 126948 112772 126954
rect 112720 126890 112772 126896
rect 112628 124160 112680 124166
rect 112628 124102 112680 124108
rect 112536 122800 112588 122806
rect 112536 122742 112588 122748
rect 112444 118652 112496 118658
rect 112444 118594 112496 118600
rect 111616 117292 111668 117298
rect 111616 117234 111668 117240
rect 111524 114504 111576 114510
rect 111524 114446 111576 114452
rect 111432 113144 111484 113150
rect 111432 113086 111484 113092
rect 111340 111784 111392 111790
rect 111340 111726 111392 111732
rect 111248 92472 111300 92478
rect 111248 92414 111300 92420
rect 111064 89684 111116 89690
rect 111064 89626 111116 89632
rect 113836 88330 113864 144191
rect 115216 135561 115244 150486
rect 115308 141409 115336 151574
rect 116044 143313 116072 151642
rect 116952 151496 117004 151502
rect 116952 151438 117004 151444
rect 116768 151428 116820 151434
rect 116768 151370 116820 151376
rect 116676 151360 116728 151366
rect 116676 151302 116728 151308
rect 116124 150476 116176 150482
rect 116124 150418 116176 150424
rect 116136 145217 116164 150418
rect 116492 150136 116544 150142
rect 116492 150078 116544 150084
rect 116400 150068 116452 150074
rect 116400 150010 116452 150016
rect 116122 145208 116178 145217
rect 116122 145143 116178 145152
rect 116030 143304 116086 143313
rect 116030 143239 116086 143248
rect 115294 141400 115350 141409
rect 115294 141335 115350 141344
rect 116124 140752 116176 140758
rect 116124 140694 116176 140700
rect 116136 139505 116164 140694
rect 116122 139496 116178 139505
rect 116122 139431 116178 139440
rect 116124 137964 116176 137970
rect 116124 137906 116176 137912
rect 116136 137601 116164 137906
rect 116122 137592 116178 137601
rect 116122 137527 116178 137536
rect 116308 137352 116360 137358
rect 116308 137294 116360 137300
rect 115202 135552 115258 135561
rect 115202 135487 115258 135496
rect 116032 133884 116084 133890
rect 116032 133826 116084 133832
rect 116044 133657 116072 133826
rect 116030 133648 116086 133657
rect 116030 133583 116086 133592
rect 114190 132832 114246 132841
rect 114190 132767 114246 132776
rect 114204 132666 114232 132767
rect 114192 132660 114244 132666
rect 114192 132602 114244 132608
rect 115204 132660 115256 132666
rect 115204 132602 115256 132608
rect 113914 121408 113970 121417
rect 113914 121343 113970 121352
rect 113824 88324 113876 88330
rect 113824 88266 113876 88272
rect 113928 83978 113956 121343
rect 114006 110120 114062 110129
rect 114006 110055 114062 110064
rect 113916 83972 113968 83978
rect 113916 83914 113968 83920
rect 114020 82822 114048 110055
rect 114098 98696 114154 98705
rect 114098 98631 114154 98640
rect 114008 82816 114060 82822
rect 114008 82758 114060 82764
rect 114112 80034 114140 98631
rect 114190 87272 114246 87281
rect 114190 87207 114246 87216
rect 114100 80028 114152 80034
rect 114100 79970 114152 79976
rect 114204 78674 114232 87207
rect 115216 85649 115244 132602
rect 116124 132456 116176 132462
rect 116124 132398 116176 132404
rect 116136 131753 116164 132398
rect 116122 131744 116178 131753
rect 116122 131679 116178 131688
rect 116320 127945 116348 137294
rect 116412 129849 116440 150010
rect 116504 137358 116532 150078
rect 116582 149696 116638 149705
rect 116582 149631 116638 149640
rect 116492 137352 116544 137358
rect 116492 137294 116544 137300
rect 116398 129840 116454 129849
rect 116398 129775 116454 129784
rect 116306 127936 116362 127945
rect 116306 127871 116362 127880
rect 116032 126948 116084 126954
rect 116032 126890 116084 126896
rect 116044 126041 116072 126890
rect 116030 126032 116086 126041
rect 116030 125967 116086 125976
rect 116124 124160 116176 124166
rect 116122 124128 116124 124137
rect 116176 124128 116178 124137
rect 116122 124063 116178 124072
rect 115940 122800 115992 122806
rect 115940 122742 115992 122748
rect 115952 122233 115980 122742
rect 115938 122224 115994 122233
rect 115938 122159 115994 122168
rect 116124 121440 116176 121446
rect 116124 121382 116176 121388
rect 116136 120193 116164 121382
rect 116122 120184 116178 120193
rect 116122 120119 116178 120128
rect 116124 118652 116176 118658
rect 116124 118594 116176 118600
rect 116136 118289 116164 118594
rect 116122 118280 116178 118289
rect 116122 118215 116178 118224
rect 116492 118040 116544 118046
rect 116492 117982 116544 117988
rect 116124 117292 116176 117298
rect 116124 117234 116176 117240
rect 116136 116385 116164 117234
rect 116122 116376 116178 116385
rect 116122 116311 116178 116320
rect 116124 114504 116176 114510
rect 116122 114472 116124 114481
rect 116176 114472 116178 114481
rect 116122 114407 116178 114416
rect 115940 113144 115992 113150
rect 115940 113086 115992 113092
rect 115952 112577 115980 113086
rect 115938 112568 115994 112577
rect 115938 112503 115994 112512
rect 116124 111784 116176 111790
rect 116124 111726 116176 111732
rect 116136 110673 116164 111726
rect 116122 110664 116178 110673
rect 116122 110599 116178 110608
rect 116124 108996 116176 109002
rect 116124 108938 116176 108944
rect 116136 108769 116164 108938
rect 116122 108760 116178 108769
rect 116122 108695 116178 108704
rect 116504 106865 116532 117982
rect 116490 106856 116546 106865
rect 116490 106791 116546 106800
rect 116596 93401 116624 149631
rect 116688 95305 116716 151302
rect 116780 97209 116808 151370
rect 116858 149832 116914 149841
rect 116858 149767 116914 149776
rect 116872 99113 116900 149767
rect 116964 102921 116992 151438
rect 117228 150272 117280 150278
rect 117228 150214 117280 150220
rect 117044 150204 117096 150210
rect 117044 150146 117096 150152
rect 116950 102912 117006 102921
rect 116950 102847 117006 102856
rect 117056 101017 117084 150146
rect 117136 148368 117188 148374
rect 117136 148310 117188 148316
rect 117148 104825 117176 148310
rect 117240 118046 117268 150214
rect 118896 149954 118924 157966
rect 120092 153950 120120 158918
rect 121288 156670 121316 163200
rect 120448 156664 120500 156670
rect 120448 156606 120500 156612
rect 121276 156664 121328 156670
rect 121276 156606 121328 156612
rect 119804 153944 119856 153950
rect 119804 153886 119856 153892
rect 120080 153944 120132 153950
rect 120080 153886 120132 153892
rect 119816 150226 119844 153886
rect 120460 150226 120488 156606
rect 122012 155372 122064 155378
rect 122012 155314 122064 155320
rect 121920 154352 121972 154358
rect 121920 154294 121972 154300
rect 121932 153950 121960 154294
rect 121920 153944 121972 153950
rect 121920 153886 121972 153892
rect 121736 153876 121788 153882
rect 121736 153818 121788 153824
rect 121090 153096 121146 153105
rect 121090 153031 121146 153040
rect 121104 150226 121132 153031
rect 121748 150226 121776 153818
rect 122024 151814 122052 155314
rect 122116 154630 122144 163200
rect 122748 158976 122800 158982
rect 122562 158944 122618 158953
rect 122748 158918 122800 158924
rect 122562 158879 122564 158888
rect 122616 158879 122618 158888
rect 122564 158850 122616 158856
rect 122760 158778 122788 158918
rect 122944 158778 122972 163200
rect 122748 158772 122800 158778
rect 122748 158714 122800 158720
rect 122932 158772 122984 158778
rect 122932 158714 122984 158720
rect 123772 155378 123800 163200
rect 124036 159656 124088 159662
rect 124036 159598 124088 159604
rect 123850 159488 123906 159497
rect 123850 159423 123906 159432
rect 123760 155372 123812 155378
rect 123760 155314 123812 155320
rect 123024 155236 123076 155242
rect 123024 155178 123076 155184
rect 122104 154624 122156 154630
rect 122104 154566 122156 154572
rect 122024 151786 122420 151814
rect 122392 150226 122420 151786
rect 123036 150226 123064 155178
rect 123864 153105 123892 159423
rect 124048 158846 124076 159598
rect 124494 158944 124550 158953
rect 124494 158879 124550 158888
rect 123944 158840 123996 158846
rect 123944 158782 123996 158788
rect 124036 158840 124088 158846
rect 124036 158782 124088 158788
rect 123956 154358 123984 158782
rect 123944 154352 123996 154358
rect 123944 154294 123996 154300
rect 124508 153785 124536 158879
rect 124600 156126 124628 163200
rect 124588 156120 124640 156126
rect 124588 156062 124640 156068
rect 125520 156058 125548 163200
rect 126348 160138 126376 163200
rect 126336 160132 126388 160138
rect 126336 160074 126388 160080
rect 127176 159662 127204 163200
rect 127164 159656 127216 159662
rect 127164 159598 127216 159604
rect 127256 159588 127308 159594
rect 127256 159530 127308 159536
rect 127624 159588 127676 159594
rect 127624 159530 127676 159536
rect 125508 156052 125560 156058
rect 125508 155994 125560 156000
rect 125600 155304 125652 155310
rect 125600 155246 125652 155252
rect 124954 153912 125010 153921
rect 124954 153847 125010 153856
rect 124310 153776 124366 153785
rect 124310 153711 124366 153720
rect 124494 153776 124550 153785
rect 124494 153711 124550 153720
rect 123850 153096 123906 153105
rect 123850 153031 123906 153040
rect 123666 152416 123722 152425
rect 123666 152351 123722 152360
rect 123680 150226 123708 152351
rect 124324 150226 124352 153711
rect 124968 150226 124996 153847
rect 125612 150226 125640 155246
rect 126886 154048 126942 154057
rect 126886 153983 126942 153992
rect 126242 153096 126298 153105
rect 126242 153031 126298 153040
rect 126256 150226 126284 153031
rect 126900 150226 126928 153983
rect 127268 151978 127296 159530
rect 127636 159390 127664 159530
rect 127624 159384 127676 159390
rect 127624 159326 127676 159332
rect 128004 156806 128032 163200
rect 128360 160132 128412 160138
rect 128360 160074 128412 160080
rect 127992 156800 128044 156806
rect 127992 156742 128044 156748
rect 127440 155984 127492 155990
rect 127440 155926 127492 155932
rect 127348 154352 127400 154358
rect 127348 154294 127400 154300
rect 127360 154057 127388 154294
rect 127346 154048 127402 154057
rect 127346 153983 127402 153992
rect 127256 151972 127308 151978
rect 127256 151914 127308 151920
rect 127452 151814 127480 155926
rect 127532 154352 127584 154358
rect 127532 154294 127584 154300
rect 127544 153950 127572 154294
rect 127532 153944 127584 153950
rect 127532 153886 127584 153892
rect 128372 153882 128400 160074
rect 128452 155372 128504 155378
rect 128452 155314 128504 155320
rect 128360 153876 128412 153882
rect 128360 153818 128412 153824
rect 128464 152114 128492 155314
rect 128832 155242 128860 163200
rect 129660 159390 129688 163200
rect 129648 159384 129700 159390
rect 129648 159326 129700 159332
rect 128820 155236 128872 155242
rect 128820 155178 128872 155184
rect 129464 154080 129516 154086
rect 129556 154080 129608 154086
rect 129464 154022 129516 154028
rect 129554 154048 129556 154057
rect 129608 154048 129610 154057
rect 128820 152516 128872 152522
rect 128820 152458 128872 152464
rect 128176 152108 128228 152114
rect 128176 152050 128228 152056
rect 128452 152108 128504 152114
rect 128452 152050 128504 152056
rect 127452 151786 127572 151814
rect 127544 150226 127572 151786
rect 128188 150226 128216 152050
rect 128832 150226 128860 152458
rect 129476 150226 129504 154022
rect 129554 153983 129610 153992
rect 129752 152522 129780 163254
rect 130396 163146 130424 163254
rect 130474 163200 130530 164400
rect 131394 163200 131450 164400
rect 132222 163200 132278 164400
rect 133050 163200 133106 164400
rect 133878 163200 133934 164400
rect 134706 163200 134762 164400
rect 135534 163200 135590 164400
rect 136362 163200 136418 164400
rect 137190 163200 137246 164400
rect 138110 163200 138166 164400
rect 138938 163200 138994 164400
rect 139766 163200 139822 164400
rect 140594 163200 140650 164400
rect 141422 163200 141478 164400
rect 142250 163200 142306 164400
rect 143078 163200 143134 164400
rect 143552 163254 143856 163282
rect 130488 163146 130516 163200
rect 130396 163118 130516 163146
rect 131302 159352 131358 159361
rect 131302 159287 131358 159296
rect 130108 156732 130160 156738
rect 130108 156674 130160 156680
rect 129740 152516 129792 152522
rect 129740 152458 129792 152464
rect 130120 150226 130148 156674
rect 130752 152244 130804 152250
rect 130752 152186 130804 152192
rect 130764 150226 130792 152186
rect 131316 151814 131344 159287
rect 131408 155990 131436 163200
rect 131396 155984 131448 155990
rect 131396 155926 131448 155932
rect 132236 155310 132264 163200
rect 132868 159520 132920 159526
rect 132868 159462 132920 159468
rect 132684 156936 132736 156942
rect 132684 156878 132736 156884
rect 132224 155304 132276 155310
rect 132224 155246 132276 155252
rect 132040 154012 132092 154018
rect 132040 153954 132092 153960
rect 131316 151786 131436 151814
rect 131408 150226 131436 151786
rect 132052 150226 132080 153954
rect 132696 150226 132724 156878
rect 132880 153105 132908 159462
rect 133064 159458 133092 163200
rect 133604 159928 133656 159934
rect 133604 159870 133656 159876
rect 133696 159928 133748 159934
rect 133696 159870 133748 159876
rect 133616 159769 133644 159870
rect 133602 159760 133658 159769
rect 133602 159695 133658 159704
rect 133708 159594 133736 159870
rect 133696 159588 133748 159594
rect 133696 159530 133748 159536
rect 133788 159588 133840 159594
rect 133788 159530 133840 159536
rect 133052 159452 133104 159458
rect 133052 159394 133104 159400
rect 133800 159050 133828 159530
rect 133892 159050 133920 163200
rect 133788 159044 133840 159050
rect 133788 158986 133840 158992
rect 133880 159044 133932 159050
rect 133880 158986 133932 158992
rect 134720 158030 134748 163200
rect 135168 158840 135220 158846
rect 135168 158782 135220 158788
rect 134708 158024 134760 158030
rect 134708 157966 134760 157972
rect 134614 154184 134670 154193
rect 134614 154119 134670 154128
rect 132866 153096 132922 153105
rect 132866 153031 132922 153040
rect 133328 152584 133380 152590
rect 133328 152526 133380 152532
rect 133970 152552 134026 152561
rect 133340 150226 133368 152526
rect 133970 152487 134026 152496
rect 133984 150226 134012 152487
rect 134628 150226 134656 154119
rect 135180 152250 135208 158782
rect 135548 156874 135576 163200
rect 136376 159662 136404 163200
rect 137100 159928 137152 159934
rect 137100 159870 137152 159876
rect 136272 159656 136324 159662
rect 136272 159598 136324 159604
rect 136364 159656 136416 159662
rect 136364 159598 136416 159604
rect 136284 158846 136312 159598
rect 136548 159520 136600 159526
rect 136548 159462 136600 159468
rect 136272 158840 136324 158846
rect 136272 158782 136324 158788
rect 135260 156868 135312 156874
rect 135260 156810 135312 156816
rect 135536 156868 135588 156874
rect 135536 156810 135588 156816
rect 135168 152244 135220 152250
rect 135168 152186 135220 152192
rect 135272 150226 135300 156810
rect 136088 154216 136140 154222
rect 136088 154158 136140 154164
rect 136100 154018 136128 154158
rect 136088 154012 136140 154018
rect 136088 153954 136140 153960
rect 135904 151972 135956 151978
rect 135904 151914 135956 151920
rect 135916 150226 135944 151914
rect 136560 150226 136588 159462
rect 137112 159338 137140 159870
rect 137204 159526 137232 163200
rect 137284 159928 137336 159934
rect 137284 159870 137336 159876
rect 137296 159730 137324 159870
rect 137374 159760 137430 159769
rect 137284 159724 137336 159730
rect 137374 159695 137376 159704
rect 137284 159666 137336 159672
rect 137428 159695 137430 159704
rect 137376 159666 137428 159672
rect 137192 159520 137244 159526
rect 137192 159462 137244 159468
rect 137112 159310 137600 159338
rect 137192 157004 137244 157010
rect 137192 156946 137244 156952
rect 137100 154148 137152 154154
rect 137100 154090 137152 154096
rect 137112 150498 137140 154090
rect 137204 151814 137232 156946
rect 137284 154284 137336 154290
rect 137284 154226 137336 154232
rect 137296 154086 137324 154226
rect 137572 154154 137600 159310
rect 138124 156942 138152 163200
rect 138112 156936 138164 156942
rect 138112 156878 138164 156884
rect 138952 156738 138980 163200
rect 139780 159730 139808 163200
rect 139308 159724 139360 159730
rect 139308 159666 139360 159672
rect 139768 159724 139820 159730
rect 139768 159666 139820 159672
rect 138940 156732 138992 156738
rect 138940 156674 138992 156680
rect 137560 154148 137612 154154
rect 137560 154090 137612 154096
rect 137284 154080 137336 154086
rect 137284 154022 137336 154028
rect 137284 152856 137336 152862
rect 137284 152798 137336 152804
rect 137296 152590 137324 152798
rect 139124 152788 139176 152794
rect 139124 152730 139176 152736
rect 139216 152788 139268 152794
rect 139216 152730 139268 152736
rect 138478 152688 138534 152697
rect 138478 152623 138534 152632
rect 137284 152584 137336 152590
rect 137284 152526 137336 152532
rect 137204 151786 137876 151814
rect 137112 150470 137232 150498
rect 137204 150226 137232 150470
rect 137848 150226 137876 151786
rect 138492 150226 138520 152623
rect 139136 150226 139164 152730
rect 139228 152250 139256 152730
rect 139320 152250 139348 159666
rect 139398 159624 139454 159633
rect 140608 159594 140636 163200
rect 139398 159559 139454 159568
rect 139492 159588 139544 159594
rect 139412 152862 139440 159559
rect 139492 159530 139544 159536
rect 140596 159588 140648 159594
rect 140596 159530 140648 159536
rect 139504 154222 139532 159530
rect 141436 157418 141464 163200
rect 141424 157412 141476 157418
rect 141424 157354 141476 157360
rect 142264 157078 142292 163200
rect 142724 160126 143028 160154
rect 142724 159934 142752 160126
rect 142804 160064 142856 160070
rect 142804 160006 142856 160012
rect 142896 160064 142948 160070
rect 142896 160006 142948 160012
rect 142816 159934 142844 160006
rect 142712 159928 142764 159934
rect 142712 159870 142764 159876
rect 142804 159928 142856 159934
rect 142804 159870 142856 159876
rect 142804 159520 142856 159526
rect 142804 159462 142856 159468
rect 142816 157334 142844 159462
rect 142908 159390 142936 160006
rect 143000 159526 143028 160126
rect 142988 159520 143040 159526
rect 142988 159462 143040 159468
rect 142896 159384 142948 159390
rect 142896 159326 142948 159332
rect 142988 159384 143040 159390
rect 142988 159326 143040 159332
rect 143000 158778 143028 159326
rect 143092 158778 143120 163200
rect 142988 158772 143040 158778
rect 142988 158714 143040 158720
rect 143080 158772 143132 158778
rect 143080 158714 143132 158720
rect 142816 157306 142936 157334
rect 139952 157072 140004 157078
rect 139952 157014 140004 157020
rect 142252 157072 142304 157078
rect 142252 157014 142304 157020
rect 139492 154216 139544 154222
rect 139492 154158 139544 154164
rect 139768 154012 139820 154018
rect 139768 153954 139820 153960
rect 139400 152856 139452 152862
rect 139400 152798 139452 152804
rect 139216 152244 139268 152250
rect 139216 152186 139268 152192
rect 139308 152244 139360 152250
rect 139308 152186 139360 152192
rect 139780 150226 139808 153954
rect 139964 151814 139992 157014
rect 142344 154080 142396 154086
rect 142344 154022 142396 154028
rect 141054 153096 141110 153105
rect 141054 153031 141110 153040
rect 139964 151786 140452 151814
rect 140424 150226 140452 151786
rect 141068 150226 141096 153031
rect 141700 152856 141752 152862
rect 141700 152798 141752 152804
rect 141792 152856 141844 152862
rect 141792 152798 141844 152804
rect 141712 150226 141740 152798
rect 141804 152250 141832 152798
rect 141792 152244 141844 152250
rect 141792 152186 141844 152192
rect 142356 150226 142384 154022
rect 142908 151978 142936 157306
rect 142988 157140 143040 157146
rect 142988 157082 143040 157088
rect 142896 151972 142948 151978
rect 142896 151914 142948 151920
rect 143000 150226 143028 157082
rect 143552 152250 143580 163254
rect 143828 163146 143856 163254
rect 143906 163200 143962 164400
rect 144826 163200 144882 164400
rect 144932 163254 145604 163282
rect 143920 163146 143948 163200
rect 143828 163118 143948 163146
rect 144460 159520 144512 159526
rect 144460 159462 144512 159468
rect 144472 152658 144500 159462
rect 144840 157010 144868 163200
rect 144828 157004 144880 157010
rect 144828 156946 144880 156952
rect 144932 154086 144960 163254
rect 145576 163146 145604 163254
rect 145654 163200 145710 164400
rect 146482 163200 146538 164400
rect 146588 163254 147076 163282
rect 145668 163146 145696 163200
rect 145576 163118 145696 163146
rect 146496 163146 146524 163200
rect 146588 163146 146616 163254
rect 146496 163118 146616 163146
rect 146300 158092 146352 158098
rect 146300 158034 146352 158040
rect 145010 157992 145066 158001
rect 145010 157927 145066 157936
rect 144920 154080 144972 154086
rect 144920 154022 144972 154028
rect 143632 152652 143684 152658
rect 143632 152594 143684 152600
rect 144460 152652 144512 152658
rect 144460 152594 144512 152600
rect 143540 152244 143592 152250
rect 143540 152186 143592 152192
rect 143644 150226 143672 152594
rect 144276 152584 144328 152590
rect 144276 152526 144328 152532
rect 144288 150226 144316 152526
rect 145024 150226 145052 157927
rect 145102 156632 145158 156641
rect 145102 156567 145158 156576
rect 119816 150198 119890 150226
rect 120460 150198 120534 150226
rect 121104 150198 121178 150226
rect 121748 150198 121822 150226
rect 122392 150198 122466 150226
rect 123036 150198 123110 150226
rect 123680 150198 123754 150226
rect 124324 150198 124398 150226
rect 124968 150198 125042 150226
rect 125612 150198 125686 150226
rect 126256 150198 126330 150226
rect 126900 150198 126974 150226
rect 127544 150198 127618 150226
rect 128188 150198 128262 150226
rect 128832 150198 128906 150226
rect 129476 150198 129550 150226
rect 130120 150198 130194 150226
rect 130764 150198 130838 150226
rect 131408 150198 131482 150226
rect 132052 150198 132126 150226
rect 132696 150198 132770 150226
rect 133340 150198 133414 150226
rect 133984 150198 134058 150226
rect 134628 150198 134702 150226
rect 135272 150198 135346 150226
rect 135916 150198 135990 150226
rect 136560 150198 136634 150226
rect 137204 150198 137278 150226
rect 137848 150198 137922 150226
rect 138492 150198 138566 150226
rect 139136 150198 139210 150226
rect 139780 150198 139854 150226
rect 140424 150198 140498 150226
rect 141068 150198 141142 150226
rect 141712 150198 141786 150226
rect 142356 150198 142430 150226
rect 143000 150198 143074 150226
rect 143644 150198 143718 150226
rect 144288 150198 144362 150226
rect 118896 149926 119324 149954
rect 119862 149940 119890 150198
rect 120506 149940 120534 150198
rect 121150 149940 121178 150198
rect 121794 149940 121822 150198
rect 122438 149940 122466 150198
rect 123082 149940 123110 150198
rect 123726 149940 123754 150198
rect 124370 149940 124398 150198
rect 125014 149940 125042 150198
rect 125658 149940 125686 150198
rect 126302 149940 126330 150198
rect 126946 149940 126974 150198
rect 127590 149940 127618 150198
rect 128234 149940 128262 150198
rect 128878 149940 128906 150198
rect 129522 149940 129550 150198
rect 130166 149940 130194 150198
rect 130810 149940 130838 150198
rect 131454 149940 131482 150198
rect 132098 149940 132126 150198
rect 132742 149940 132770 150198
rect 133386 149940 133414 150198
rect 134030 149940 134058 150198
rect 134674 149940 134702 150198
rect 135318 149940 135346 150198
rect 135962 149940 135990 150198
rect 136606 149940 136634 150198
rect 137250 149940 137278 150198
rect 137894 149940 137922 150198
rect 138538 149940 138566 150198
rect 139182 149940 139210 150198
rect 139826 149940 139854 150198
rect 140470 149940 140498 150198
rect 141114 149940 141142 150198
rect 141758 149940 141786 150198
rect 142402 149940 142430 150198
rect 143046 149940 143074 150198
rect 143690 149940 143718 150198
rect 144334 149940 144362 150198
rect 144978 150198 145052 150226
rect 145116 150210 145144 156567
rect 145564 153264 145616 153270
rect 145564 153206 145616 153212
rect 145576 150226 145604 153206
rect 146312 151814 146340 158034
rect 147048 154494 147076 163254
rect 147310 163200 147366 164400
rect 148138 163200 148194 164400
rect 148966 163200 149022 164400
rect 149794 163200 149850 164400
rect 150622 163200 150678 164400
rect 151542 163200 151598 164400
rect 151832 163254 152320 163282
rect 147324 159526 147352 163200
rect 147312 159520 147364 159526
rect 147312 159462 147364 159468
rect 147128 159384 147180 159390
rect 147128 159326 147180 159332
rect 146760 154488 146812 154494
rect 146760 154430 146812 154436
rect 147036 154488 147088 154494
rect 147036 154430 147088 154436
rect 146576 154420 146628 154426
rect 146576 154362 146628 154368
rect 146312 151786 146432 151814
rect 145104 150204 145156 150210
rect 144978 149940 145006 150198
rect 145576 150198 145650 150226
rect 146404 150210 146432 151786
rect 145104 150146 145156 150152
rect 145622 149940 145650 150198
rect 146254 150204 146306 150210
rect 146254 150146 146306 150152
rect 146392 150204 146444 150210
rect 146392 150146 146444 150152
rect 146266 149940 146294 150146
rect 146588 150142 146616 154362
rect 146772 153950 146800 154430
rect 146944 154420 146996 154426
rect 146944 154362 146996 154368
rect 146956 154222 146984 154362
rect 147140 154222 147168 159326
rect 148152 158098 148180 163200
rect 148140 158092 148192 158098
rect 148140 158034 148192 158040
rect 148784 157208 148836 157214
rect 148784 157150 148836 157156
rect 148324 154488 148376 154494
rect 148060 154414 148272 154442
rect 148324 154430 148376 154436
rect 146944 154216 146996 154222
rect 146850 154184 146906 154193
rect 146944 154158 146996 154164
rect 147128 154216 147180 154222
rect 147128 154158 147180 154164
rect 146850 154119 146852 154128
rect 146904 154119 146906 154128
rect 146852 154090 146904 154096
rect 148060 154034 148088 154414
rect 148138 154320 148194 154329
rect 148138 154255 148194 154264
rect 147784 154006 148088 154034
rect 147784 153950 147812 154006
rect 146668 153944 146720 153950
rect 146668 153886 146720 153892
rect 146760 153944 146812 153950
rect 146760 153886 146812 153892
rect 147772 153944 147824 153950
rect 147772 153886 147824 153892
rect 146680 153270 146708 153886
rect 146668 153264 146720 153270
rect 146668 153206 146720 153212
rect 146944 152856 146996 152862
rect 146944 152798 146996 152804
rect 146956 152590 146984 152798
rect 146944 152584 146996 152590
rect 146944 152526 146996 152532
rect 146852 152040 146904 152046
rect 146852 151982 146904 151988
rect 146864 150226 146892 151982
rect 146864 150198 146938 150226
rect 146576 150136 146628 150142
rect 146576 150078 146628 150084
rect 146910 149940 146938 150198
rect 147542 150204 147594 150210
rect 147542 150146 147594 150152
rect 147554 149940 147582 150146
rect 148152 150090 148180 154255
rect 148244 154222 148272 154414
rect 148232 154216 148284 154222
rect 148232 154158 148284 154164
rect 148336 154018 148364 154430
rect 148324 154012 148376 154018
rect 148324 153954 148376 153960
rect 148796 150090 148824 157150
rect 148980 155378 149008 163200
rect 149808 159798 149836 163200
rect 149060 159792 149112 159798
rect 149060 159734 149112 159740
rect 149796 159792 149848 159798
rect 149796 159734 149848 159740
rect 148968 155372 149020 155378
rect 148968 155314 149020 155320
rect 149072 152862 149100 159734
rect 150636 159390 150664 163200
rect 150624 159384 150676 159390
rect 150624 159326 150676 159332
rect 149610 158128 149666 158137
rect 149610 158063 149666 158072
rect 149624 157334 149652 158063
rect 149624 157306 150020 157334
rect 149060 152856 149112 152862
rect 149060 152798 149112 152804
rect 149428 152788 149480 152794
rect 149428 152730 149480 152736
rect 149440 150090 149468 152730
rect 149992 150226 150020 157306
rect 151556 157146 151584 163200
rect 151832 157214 151860 163254
rect 152292 163146 152320 163254
rect 152370 163200 152426 164400
rect 153198 163200 153254 164400
rect 154026 163200 154082 164400
rect 154854 163200 154910 164400
rect 155682 163200 155738 164400
rect 156510 163200 156566 164400
rect 157338 163200 157394 164400
rect 158258 163200 158314 164400
rect 159086 163200 159142 164400
rect 159914 163200 159970 164400
rect 160742 163200 160798 164400
rect 161570 163200 161626 164400
rect 162398 163200 162454 164400
rect 163226 163200 163282 164400
rect 163516 163254 164096 163282
rect 152384 163146 152412 163200
rect 152292 163118 152412 163146
rect 153016 160132 153068 160138
rect 153016 160074 153068 160080
rect 153028 159866 153056 160074
rect 153212 159934 153240 163200
rect 153200 159928 153252 159934
rect 153200 159870 153252 159876
rect 153016 159860 153068 159866
rect 153016 159802 153068 159808
rect 154040 159390 154068 163200
rect 154488 160064 154540 160070
rect 154488 160006 154540 160012
rect 154396 159860 154448 159866
rect 154396 159802 154448 159808
rect 152740 159384 152792 159390
rect 152740 159326 152792 159332
rect 154028 159384 154080 159390
rect 154028 159326 154080 159332
rect 152370 158264 152426 158273
rect 152370 158199 152426 158208
rect 152384 157334 152412 158199
rect 152292 157306 152412 157334
rect 152752 157334 152780 159326
rect 153016 158296 153068 158302
rect 153014 158264 153016 158273
rect 153068 158264 153070 158273
rect 153014 158199 153070 158208
rect 153108 158228 153160 158234
rect 153108 158170 153160 158176
rect 153120 158114 153148 158170
rect 153476 158160 153528 158166
rect 153120 158108 153476 158114
rect 153120 158102 153528 158108
rect 153120 158086 153516 158102
rect 153844 157344 153896 157350
rect 152752 157306 152872 157334
rect 151820 157208 151872 157214
rect 151820 157150 151872 157156
rect 151544 157140 151596 157146
rect 151544 157082 151596 157088
rect 151266 156768 151322 156777
rect 151266 156703 151322 156712
rect 149992 150198 150066 150226
rect 148152 150062 148226 150090
rect 148796 150062 148870 150090
rect 149440 150062 149514 150090
rect 148198 149940 148226 150062
rect 148842 149940 148870 150062
rect 149486 149940 149514 150062
rect 150038 149940 150066 150198
rect 150670 150136 150722 150142
rect 150670 150078 150722 150084
rect 151280 150090 151308 156703
rect 151728 155440 151780 155446
rect 151728 155382 151780 155388
rect 151740 155145 151768 155382
rect 151726 155136 151782 155145
rect 151726 155071 151782 155080
rect 151912 151904 151964 151910
rect 151912 151846 151964 151852
rect 151924 150090 151952 151846
rect 152292 150226 152320 157306
rect 152740 155440 152792 155446
rect 152740 155382 152792 155388
rect 152752 155145 152780 155382
rect 152738 155136 152794 155145
rect 152738 155071 152794 155080
rect 152740 154556 152792 154562
rect 152740 154498 152792 154504
rect 152752 154442 152780 154498
rect 152384 154426 152780 154442
rect 152372 154420 152780 154426
rect 152424 154414 152780 154420
rect 152372 154362 152424 154368
rect 152844 152794 152872 157306
rect 153844 157286 153896 157292
rect 152924 157208 152976 157214
rect 152924 157150 152976 157156
rect 152936 154086 152964 157150
rect 153016 154488 153068 154494
rect 153016 154430 153068 154436
rect 153028 154193 153056 154430
rect 153200 154216 153252 154222
rect 153014 154184 153070 154193
rect 153200 154158 153252 154164
rect 153014 154119 153070 154128
rect 152924 154080 152976 154086
rect 152924 154022 152976 154028
rect 152832 152788 152884 152794
rect 152832 152730 152884 152736
rect 152292 150198 152642 150226
rect 150682 149940 150710 150078
rect 151280 150062 151354 150090
rect 151924 150062 151998 150090
rect 151326 149940 151354 150062
rect 151970 149940 151998 150062
rect 152614 149940 152642 150198
rect 153212 150090 153240 154158
rect 153856 150090 153884 157286
rect 154408 152266 154436 159802
rect 154500 154222 154528 160006
rect 154868 158234 154896 163200
rect 155222 158264 155278 158273
rect 154856 158228 154908 158234
rect 155222 158199 155278 158208
rect 154856 158170 154908 158176
rect 155236 158166 155264 158199
rect 155132 158160 155184 158166
rect 155132 158102 155184 158108
rect 155224 158160 155276 158166
rect 155224 158102 155276 158108
rect 154488 154216 154540 154222
rect 154488 154158 154540 154164
rect 154408 152238 154620 152266
rect 154592 152182 154620 152238
rect 154488 152176 154540 152182
rect 154488 152118 154540 152124
rect 154580 152176 154632 152182
rect 154580 152118 154632 152124
rect 154500 150090 154528 152118
rect 155144 150226 155172 158102
rect 155696 155446 155724 163200
rect 156524 159866 156552 163200
rect 156512 159860 156564 159866
rect 156512 159802 156564 159808
rect 156604 159452 156656 159458
rect 156604 159394 156656 159400
rect 156616 157282 156644 159394
rect 156420 157276 156472 157282
rect 156420 157218 156472 157224
rect 156604 157276 156656 157282
rect 156604 157218 156656 157224
rect 155592 155440 155644 155446
rect 155592 155382 155644 155388
rect 155684 155440 155736 155446
rect 155684 155382 155736 155388
rect 155604 150226 155632 155382
rect 155144 150198 155218 150226
rect 155604 150198 155862 150226
rect 153212 150062 153286 150090
rect 153856 150062 153930 150090
rect 154500 150062 154574 150090
rect 153258 149940 153286 150062
rect 153902 149940 153930 150062
rect 154546 149940 154574 150062
rect 155190 149940 155218 150198
rect 155834 149940 155862 150198
rect 156432 150090 156460 157218
rect 157352 152590 157380 163200
rect 158272 158302 158300 163200
rect 158812 160064 158864 160070
rect 158812 160006 158864 160012
rect 158720 159724 158772 159730
rect 158720 159666 158772 159672
rect 157432 158296 157484 158302
rect 157432 158238 157484 158244
rect 158260 158296 158312 158302
rect 158260 158238 158312 158244
rect 157064 152584 157116 152590
rect 157064 152526 157116 152532
rect 157340 152584 157392 152590
rect 157340 152526 157392 152532
rect 157076 150090 157104 152526
rect 157444 151814 157472 158238
rect 158732 157214 158760 159666
rect 158720 157208 158772 157214
rect 158720 157150 158772 157156
rect 158352 155576 158404 155582
rect 158352 155518 158404 155524
rect 157444 151786 157748 151814
rect 157720 150226 157748 151786
rect 158364 150226 158392 155518
rect 158824 152046 158852 160006
rect 158994 156904 159050 156913
rect 158994 156839 159050 156848
rect 158812 152040 158864 152046
rect 158812 151982 158864 151988
rect 159008 150226 159036 156839
rect 159100 155582 159128 163200
rect 159928 160070 159956 163200
rect 159916 160064 159968 160070
rect 159916 160006 159968 160012
rect 160756 159458 160784 163200
rect 160744 159452 160796 159458
rect 160744 159394 160796 159400
rect 161584 158166 161612 163200
rect 162124 158432 162176 158438
rect 162176 158380 162348 158386
rect 162124 158374 162348 158380
rect 162136 158370 162348 158374
rect 162136 158364 162360 158370
rect 162136 158358 162308 158364
rect 162308 158306 162360 158312
rect 161940 158296 161992 158302
rect 162216 158296 162268 158302
rect 161992 158244 162216 158250
rect 161940 158238 162268 158244
rect 161952 158222 162256 158238
rect 160100 158160 160152 158166
rect 160100 158102 160152 158108
rect 161572 158160 161624 158166
rect 161572 158102 161624 158108
rect 159088 155576 159140 155582
rect 159088 155518 159140 155524
rect 159640 152652 159692 152658
rect 159640 152594 159692 152600
rect 159652 150226 159680 152594
rect 160112 151814 160140 158102
rect 161570 157040 161626 157049
rect 161570 156975 161626 156984
rect 160928 155508 160980 155514
rect 160928 155450 160980 155456
rect 160112 151786 160324 151814
rect 160296 150226 160324 151786
rect 160940 150226 160968 155450
rect 161584 150226 161612 156975
rect 162412 155514 162440 163200
rect 163240 159662 163268 163200
rect 163228 159656 163280 159662
rect 163228 159598 163280 159604
rect 162950 158400 163006 158409
rect 162950 158335 163006 158344
rect 162400 155508 162452 155514
rect 162400 155450 162452 155456
rect 162216 152312 162268 152318
rect 162216 152254 162268 152260
rect 162228 150226 162256 152254
rect 162964 150226 162992 158335
rect 163410 155408 163466 155417
rect 163410 155343 163466 155352
rect 163320 154420 163372 154426
rect 163320 154362 163372 154368
rect 157720 150198 157794 150226
rect 158364 150198 158438 150226
rect 159008 150198 159082 150226
rect 159652 150198 159726 150226
rect 160296 150198 160370 150226
rect 160940 150198 161014 150226
rect 161584 150198 161658 150226
rect 162228 150198 162302 150226
rect 156432 150062 156506 150090
rect 157076 150062 157150 150090
rect 156478 149940 156506 150062
rect 157122 149940 157150 150062
rect 157766 149940 157794 150198
rect 158410 149940 158438 150198
rect 159054 149940 159082 150198
rect 159698 149940 159726 150198
rect 160342 149940 160370 150198
rect 160986 149940 161014 150198
rect 161630 149940 161658 150198
rect 162274 149940 162302 150198
rect 162918 150198 162992 150226
rect 163332 150210 163360 154362
rect 163424 151814 163452 155343
rect 163516 152658 163544 163254
rect 164068 163146 164096 163254
rect 164146 163200 164202 164400
rect 164974 163200 165030 164400
rect 165802 163200 165858 164400
rect 166630 163200 166686 164400
rect 167458 163200 167514 164400
rect 168286 163200 168342 164400
rect 169114 163200 169170 164400
rect 169942 163200 169998 164400
rect 170048 163254 170812 163282
rect 164160 163146 164188 163200
rect 164068 163118 164188 163146
rect 164516 159996 164568 160002
rect 164516 159938 164568 159944
rect 164148 159724 164200 159730
rect 164148 159666 164200 159672
rect 164160 154426 164188 159666
rect 164332 158500 164384 158506
rect 164332 158442 164384 158448
rect 164424 158500 164476 158506
rect 164424 158442 164476 158448
rect 164148 154420 164200 154426
rect 164148 154362 164200 154368
rect 163504 152652 163556 152658
rect 163504 152594 163556 152600
rect 163424 151786 163544 151814
rect 163516 150226 163544 151786
rect 163320 150204 163372 150210
rect 162918 149940 162946 150198
rect 163516 150198 163590 150226
rect 164344 150210 164372 158442
rect 164436 158166 164464 158442
rect 164424 158160 164476 158166
rect 164424 158102 164476 158108
rect 164528 151910 164556 159938
rect 164988 158302 165016 163200
rect 164884 158296 164936 158302
rect 164620 158234 164832 158250
rect 164884 158238 164936 158244
rect 164976 158296 165028 158302
rect 164976 158238 165028 158244
rect 164608 158228 164844 158234
rect 164660 158222 164792 158228
rect 164608 158170 164660 158176
rect 164792 158170 164844 158176
rect 164896 158166 164924 158238
rect 164884 158160 164936 158166
rect 164884 158102 164936 158108
rect 165816 154426 165844 163200
rect 166644 160002 166672 163200
rect 166632 159996 166684 160002
rect 166632 159938 166684 159944
rect 167472 159730 167500 163200
rect 167460 159724 167512 159730
rect 167460 159666 167512 159672
rect 167000 159316 167052 159322
rect 167000 159258 167052 159264
rect 166172 157208 166224 157214
rect 166172 157150 166224 157156
rect 166264 157208 166316 157214
rect 166264 157150 166316 157156
rect 166184 156482 166212 157150
rect 166276 156602 166304 157150
rect 166264 156596 166316 156602
rect 166264 156538 166316 156544
rect 166356 156596 166408 156602
rect 166356 156538 166408 156544
rect 166368 156482 166396 156538
rect 166184 156454 166396 156482
rect 166078 155272 166134 155281
rect 166078 155207 166134 155216
rect 165712 154420 165764 154426
rect 165712 154362 165764 154368
rect 165804 154420 165856 154426
rect 165804 154362 165856 154368
rect 165724 154329 165752 154362
rect 165710 154320 165766 154329
rect 165710 154255 165766 154264
rect 164884 152856 164936 152862
rect 164884 152798 164936 152804
rect 164516 151904 164568 151910
rect 164516 151846 164568 151852
rect 164896 150226 164924 152798
rect 163320 150146 163372 150152
rect 163562 149940 163590 150198
rect 164194 150204 164246 150210
rect 164194 150146 164246 150152
rect 164332 150204 164384 150210
rect 164332 150146 164384 150152
rect 164850 150198 164924 150226
rect 166092 150226 166120 155207
rect 166354 154320 166410 154329
rect 166354 154255 166410 154264
rect 166368 154154 166396 154255
rect 166264 154148 166316 154154
rect 166264 154090 166316 154096
rect 166356 154148 166408 154154
rect 166356 154090 166408 154096
rect 166276 153814 166304 154090
rect 166172 153808 166224 153814
rect 166172 153750 166224 153756
rect 166264 153808 166316 153814
rect 166264 153750 166316 153756
rect 166184 151814 166212 153750
rect 167012 152318 167040 159258
rect 168300 158438 168328 163200
rect 168288 158432 168340 158438
rect 168288 158374 168340 158380
rect 167552 158364 167604 158370
rect 167552 158306 167604 158312
rect 167000 152312 167052 152318
rect 167000 152254 167052 152260
rect 167368 151836 167420 151842
rect 166184 151786 166764 151814
rect 166736 150226 166764 151786
rect 167564 151814 167592 158306
rect 169128 155650 169156 163200
rect 169956 159322 169984 163200
rect 169944 159316 169996 159322
rect 169944 159258 169996 159264
rect 168656 155644 168708 155650
rect 168656 155586 168708 155592
rect 169116 155644 169168 155650
rect 169116 155586 169168 155592
rect 167564 151786 168052 151814
rect 167368 151778 167420 151784
rect 167380 150226 167408 151778
rect 168024 150226 168052 151786
rect 168668 150226 168696 155586
rect 169298 154456 169354 154465
rect 169298 154391 169354 154400
rect 169312 150226 169340 154391
rect 170048 152862 170076 163254
rect 170784 163146 170812 163254
rect 170862 163200 170918 164400
rect 171690 163200 171746 164400
rect 172518 163200 172574 164400
rect 172624 163254 173204 163282
rect 170876 163146 170904 163200
rect 170784 163118 170904 163146
rect 171704 158370 171732 163200
rect 172532 163146 172560 163200
rect 172624 163146 172652 163254
rect 172532 163118 172652 163146
rect 172428 159860 172480 159866
rect 172428 159802 172480 159808
rect 170588 158364 170640 158370
rect 170588 158306 170640 158312
rect 171692 158364 171744 158370
rect 171692 158306 171744 158312
rect 170036 152856 170088 152862
rect 170036 152798 170088 152804
rect 169944 152176 169996 152182
rect 169944 152118 169996 152124
rect 169956 150226 169984 152118
rect 170600 150226 170628 158306
rect 172440 157214 172468 159802
rect 172704 158636 172756 158642
rect 172704 158578 172756 158584
rect 171140 157208 171192 157214
rect 171140 157150 171192 157156
rect 172428 157208 172480 157214
rect 172428 157150 172480 157156
rect 165482 150204 165534 150210
rect 164206 149940 164234 150146
rect 164850 149940 164878 150198
rect 166092 150198 166166 150226
rect 166736 150198 166810 150226
rect 167380 150198 167454 150226
rect 168024 150198 168098 150226
rect 168668 150198 168742 150226
rect 169312 150198 169386 150226
rect 169956 150198 170030 150226
rect 170600 150198 170674 150226
rect 171152 150210 171180 157150
rect 171230 155544 171286 155553
rect 171230 155479 171286 155488
rect 171244 150226 171272 155479
rect 172520 152040 172572 152046
rect 172520 151982 172572 151988
rect 172532 150226 172560 151982
rect 172716 151814 172744 158578
rect 173176 155718 173204 163254
rect 173346 163200 173402 164400
rect 174174 163200 174230 164400
rect 175002 163200 175058 164400
rect 175476 163254 175780 163282
rect 173360 159254 173388 163200
rect 174188 159662 174216 163200
rect 174084 159656 174136 159662
rect 174084 159598 174136 159604
rect 174176 159656 174228 159662
rect 174176 159598 174228 159604
rect 173256 159248 173308 159254
rect 173256 159190 173308 159196
rect 173348 159248 173400 159254
rect 173348 159190 173400 159196
rect 173072 155712 173124 155718
rect 173072 155654 173124 155660
rect 173164 155712 173216 155718
rect 173164 155654 173216 155660
rect 173084 151814 173112 155654
rect 173268 151910 173296 159190
rect 174096 159118 174124 159598
rect 173992 159112 174044 159118
rect 173992 159054 174044 159060
rect 174084 159112 174136 159118
rect 174084 159054 174136 159060
rect 173900 153740 173952 153746
rect 173900 153682 173952 153688
rect 173256 151904 173308 151910
rect 173256 151846 173308 151852
rect 173912 151814 173940 153682
rect 174004 152182 174032 159054
rect 175016 158642 175044 163200
rect 175004 158636 175056 158642
rect 175004 158578 175056 158584
rect 175372 158568 175424 158574
rect 175372 158510 175424 158516
rect 175096 152448 175148 152454
rect 175096 152390 175148 152396
rect 173992 152176 174044 152182
rect 173992 152118 174044 152124
rect 172716 151786 173020 151814
rect 173084 151786 173848 151814
rect 173912 151786 174492 151814
rect 172992 150498 173020 151786
rect 172992 150470 173204 150498
rect 173176 150226 173204 150470
rect 173820 150226 173848 151786
rect 174464 150226 174492 151786
rect 175108 150226 175136 152390
rect 175384 151814 175412 158510
rect 175476 156482 175504 163254
rect 175752 163146 175780 163254
rect 175830 163200 175886 164400
rect 176658 163200 176714 164400
rect 176764 163254 177528 163282
rect 175844 163146 175872 163200
rect 175752 163118 175872 163146
rect 176672 159866 176700 163200
rect 176660 159860 176712 159866
rect 176660 159802 176712 159808
rect 176476 158772 176528 158778
rect 176476 158714 176528 158720
rect 175936 156602 176240 156618
rect 175924 156596 176240 156602
rect 175976 156590 176240 156596
rect 175924 156538 175976 156544
rect 176212 156534 176240 156590
rect 176200 156528 176252 156534
rect 175476 156454 176148 156482
rect 176200 156470 176252 156476
rect 175660 154546 176056 154574
rect 175660 153678 175688 154546
rect 176028 154426 176056 154546
rect 175924 154420 175976 154426
rect 175924 154362 175976 154368
rect 176016 154420 176068 154426
rect 176016 154362 176068 154368
rect 175832 154216 175884 154222
rect 175832 154158 175884 154164
rect 175740 154148 175792 154154
rect 175740 154090 175792 154096
rect 175752 153678 175780 154090
rect 175844 153746 175872 154158
rect 175936 154154 175964 154362
rect 176120 154222 176148 156454
rect 176488 155854 176516 158714
rect 176384 155848 176436 155854
rect 176384 155790 176436 155796
rect 176476 155848 176528 155854
rect 176476 155790 176528 155796
rect 176108 154216 176160 154222
rect 176108 154158 176160 154164
rect 175924 154148 175976 154154
rect 175924 154090 175976 154096
rect 175832 153740 175884 153746
rect 175832 153682 175884 153688
rect 175648 153672 175700 153678
rect 175648 153614 175700 153620
rect 175740 153672 175792 153678
rect 175740 153614 175792 153620
rect 175384 151786 175780 151814
rect 175752 150226 175780 151786
rect 176396 150226 176424 155790
rect 176764 152454 176792 163254
rect 177500 163146 177528 163254
rect 177578 163200 177634 164400
rect 178406 163200 178462 164400
rect 179234 163200 179290 164400
rect 180062 163200 180118 164400
rect 180890 163200 180946 164400
rect 181718 163200 181774 164400
rect 182546 163200 182602 164400
rect 183374 163200 183430 164400
rect 184294 163200 184350 164400
rect 185122 163200 185178 164400
rect 185950 163200 186006 164400
rect 186778 163200 186834 164400
rect 187606 163200 187662 164400
rect 188434 163200 188490 164400
rect 189262 163200 189318 164400
rect 190090 163200 190146 164400
rect 190564 163254 190960 163282
rect 177592 163146 177620 163200
rect 177500 163118 177620 163146
rect 178420 158574 178448 163200
rect 179052 159112 179104 159118
rect 179052 159054 179104 159060
rect 178408 158568 178460 158574
rect 178408 158510 178460 158516
rect 178040 157956 178092 157962
rect 178040 157898 178092 157904
rect 177028 155916 177080 155922
rect 177028 155858 177080 155864
rect 176752 152448 176804 152454
rect 176752 152390 176804 152396
rect 177040 150226 177068 155858
rect 177672 151836 177724 151842
rect 178052 151814 178080 157898
rect 179064 155786 179092 159054
rect 179248 155922 179276 163200
rect 180076 158778 180104 163200
rect 180904 159798 180932 163200
rect 180800 159792 180852 159798
rect 180800 159734 180852 159740
rect 180892 159792 180944 159798
rect 180892 159734 180944 159740
rect 180812 159118 180840 159734
rect 180800 159112 180852 159118
rect 180800 159054 180852 159060
rect 181628 159112 181680 159118
rect 181628 159054 181680 159060
rect 180064 158772 180116 158778
rect 180064 158714 180116 158720
rect 180800 158704 180852 158710
rect 180800 158646 180852 158652
rect 179696 157208 179748 157214
rect 179696 157150 179748 157156
rect 179708 156602 179736 157150
rect 179604 156596 179656 156602
rect 179604 156538 179656 156544
rect 179696 156596 179748 156602
rect 179696 156538 179748 156544
rect 179236 155916 179288 155922
rect 179236 155858 179288 155864
rect 178960 155780 179012 155786
rect 178960 155722 179012 155728
rect 179052 155780 179104 155786
rect 179052 155722 179104 155728
rect 178052 151786 178356 151814
rect 177672 151778 177724 151784
rect 177684 150226 177712 151778
rect 178328 150226 178356 151786
rect 178972 150226 179000 155722
rect 179616 150226 179644 156538
rect 180248 152380 180300 152386
rect 180248 152322 180300 152328
rect 180260 150226 180288 152322
rect 180812 150226 180840 158646
rect 181536 157820 181588 157826
rect 181536 157762 181588 157768
rect 181548 157690 181576 157762
rect 181640 157690 181668 159054
rect 181732 158710 181760 163200
rect 181996 159860 182048 159866
rect 181996 159802 182048 159808
rect 181720 158704 181772 158710
rect 181720 158646 181772 158652
rect 181536 157684 181588 157690
rect 181536 157626 181588 157632
rect 181628 157684 181680 157690
rect 181628 157626 181680 157632
rect 181352 155168 181404 155174
rect 181352 155110 181404 155116
rect 181260 154420 181312 154426
rect 181260 154362 181312 154368
rect 165482 150146 165534 150152
rect 165494 149940 165522 150146
rect 166138 149940 166166 150198
rect 166782 149940 166810 150198
rect 167426 149940 167454 150198
rect 168070 149940 168098 150198
rect 168714 149940 168742 150198
rect 169358 149940 169386 150198
rect 170002 149940 170030 150198
rect 170646 149940 170674 150198
rect 171140 150204 171192 150210
rect 171244 150198 171318 150226
rect 171140 150146 171192 150152
rect 171290 149940 171318 150198
rect 171922 150204 171974 150210
rect 172532 150198 172606 150226
rect 173176 150198 173250 150226
rect 173820 150198 173894 150226
rect 174464 150198 174538 150226
rect 175108 150198 175182 150226
rect 175752 150198 175826 150226
rect 176396 150198 176470 150226
rect 177040 150198 177114 150226
rect 177684 150198 177758 150226
rect 178328 150198 178402 150226
rect 178972 150198 179046 150226
rect 179616 150198 179690 150226
rect 180260 150198 180334 150226
rect 180812 150198 180886 150226
rect 181272 150210 181300 154362
rect 181364 151814 181392 155110
rect 182008 154426 182036 159802
rect 182364 157752 182416 157758
rect 182364 157694 182416 157700
rect 181996 154420 182048 154426
rect 181996 154362 182048 154368
rect 181364 151786 181484 151814
rect 181456 150226 181484 151786
rect 171922 150146 171974 150152
rect 171934 149940 171962 150146
rect 172578 149940 172606 150198
rect 173222 149940 173250 150198
rect 173866 149940 173894 150198
rect 174510 149940 174538 150198
rect 175154 149940 175182 150198
rect 175798 149940 175826 150198
rect 176442 149940 176470 150198
rect 177086 149940 177114 150198
rect 177730 149940 177758 150198
rect 178374 149940 178402 150198
rect 179018 149940 179046 150198
rect 179662 149940 179690 150198
rect 180306 149940 180334 150198
rect 180858 149940 180886 150198
rect 181260 150204 181312 150210
rect 181456 150198 181530 150226
rect 182376 150210 182404 157694
rect 182560 155174 182588 163200
rect 183100 159180 183152 159186
rect 183100 159122 183152 159128
rect 182548 155168 182600 155174
rect 182548 155110 182600 155116
rect 182824 152312 182876 152318
rect 182824 152254 182876 152260
rect 182836 150226 182864 152254
rect 183112 152046 183140 159122
rect 183388 157214 183416 163200
rect 184308 159866 184336 163200
rect 184296 159860 184348 159866
rect 184296 159802 184348 159808
rect 185032 159860 185084 159866
rect 185032 159802 185084 159808
rect 183376 157208 183428 157214
rect 183376 157150 183428 157156
rect 184018 155680 184074 155689
rect 184018 155615 184074 155624
rect 183560 154964 183612 154970
rect 183560 154906 183612 154912
rect 183100 152040 183152 152046
rect 183100 151982 183152 151988
rect 181260 150146 181312 150152
rect 181502 149940 181530 150198
rect 182134 150204 182186 150210
rect 182134 150146 182186 150152
rect 182364 150204 182416 150210
rect 182364 150146 182416 150152
rect 182790 150198 182864 150226
rect 183572 150210 183600 154906
rect 184032 150226 184060 155615
rect 185044 152386 185072 159802
rect 185136 157758 185164 163200
rect 185308 157956 185360 157962
rect 185308 157898 185360 157904
rect 185124 157752 185176 157758
rect 185124 157694 185176 157700
rect 185320 154986 185348 157898
rect 185412 155910 185900 155938
rect 185412 155174 185440 155910
rect 185676 155848 185728 155854
rect 185676 155790 185728 155796
rect 185400 155168 185452 155174
rect 185400 155110 185452 155116
rect 185492 155168 185544 155174
rect 185492 155110 185544 155116
rect 185320 154958 185440 154986
rect 185308 152720 185360 152726
rect 185308 152662 185360 152668
rect 185032 152380 185084 152386
rect 185032 152322 185084 152328
rect 185320 150226 185348 152662
rect 185412 151814 185440 154958
rect 185504 154902 185532 155110
rect 185584 154964 185636 154970
rect 185584 154906 185636 154912
rect 185492 154896 185544 154902
rect 185492 154838 185544 154844
rect 185596 154766 185624 154906
rect 185688 154902 185716 155790
rect 185872 155786 185900 155910
rect 185964 155854 185992 163200
rect 186792 159118 186820 163200
rect 187620 159798 187648 163200
rect 187608 159792 187660 159798
rect 187608 159734 187660 159740
rect 186780 159112 186832 159118
rect 186780 159054 186832 159060
rect 186412 158976 186464 158982
rect 186412 158918 186464 158924
rect 185952 155848 186004 155854
rect 185952 155790 186004 155796
rect 185768 155780 185820 155786
rect 185768 155722 185820 155728
rect 185860 155780 185912 155786
rect 185860 155722 185912 155728
rect 185676 154896 185728 154902
rect 185676 154838 185728 154844
rect 185780 154766 185808 155722
rect 185584 154760 185636 154766
rect 185584 154702 185636 154708
rect 185768 154760 185820 154766
rect 185768 154702 185820 154708
rect 186424 152318 186452 158918
rect 188448 157962 188476 163200
rect 188436 157956 188488 157962
rect 188436 157898 188488 157904
rect 188528 157888 188580 157894
rect 188528 157830 188580 157836
rect 187882 156496 187938 156505
rect 187882 156431 187884 156440
rect 187936 156431 187938 156440
rect 187884 156402 187936 156408
rect 187240 156392 187292 156398
rect 187240 156334 187292 156340
rect 186596 155100 186648 155106
rect 186596 155042 186648 155048
rect 186412 152312 186464 152318
rect 186412 152254 186464 152260
rect 185412 151786 185992 151814
rect 185964 150226 185992 151786
rect 183422 150204 183474 150210
rect 182146 149940 182174 150146
rect 182790 149940 182818 150198
rect 183422 150146 183474 150152
rect 183560 150204 183612 150210
rect 184032 150198 184106 150226
rect 183560 150146 183612 150152
rect 183434 149940 183462 150146
rect 184078 149940 184106 150198
rect 184710 150204 184762 150210
rect 185320 150198 185394 150226
rect 185964 150198 186038 150226
rect 184710 150146 184762 150152
rect 184722 149940 184750 150146
rect 185366 149940 185394 150198
rect 186010 149940 186038 150198
rect 186608 150090 186636 155042
rect 187252 150090 187280 156334
rect 187884 151904 187936 151910
rect 187884 151846 187936 151852
rect 187896 150090 187924 151846
rect 188540 150226 188568 157830
rect 189276 155174 189304 163200
rect 189724 159928 189776 159934
rect 189724 159870 189776 159876
rect 189264 155168 189316 155174
rect 189264 155110 189316 155116
rect 189172 155032 189224 155038
rect 189172 154974 189224 154980
rect 189184 150226 189212 154974
rect 189540 154284 189592 154290
rect 189540 154226 189592 154232
rect 189446 153368 189502 153377
rect 189446 153303 189502 153312
rect 189460 153270 189488 153303
rect 189552 153270 189580 154226
rect 189736 153649 189764 159870
rect 190104 157894 190132 163200
rect 190092 157888 190144 157894
rect 190092 157830 190144 157836
rect 189816 154352 189868 154358
rect 189816 154294 189868 154300
rect 189722 153640 189778 153649
rect 189722 153575 189778 153584
rect 189448 153264 189500 153270
rect 189448 153206 189500 153212
rect 189540 153264 189592 153270
rect 189540 153206 189592 153212
rect 188540 150198 188614 150226
rect 189184 150198 189258 150226
rect 186608 150062 186682 150090
rect 187252 150062 187326 150090
rect 187896 150062 187970 150090
rect 186654 149940 186682 150062
rect 187298 149940 187326 150062
rect 187942 149940 187970 150062
rect 188586 149940 188614 150198
rect 189230 149940 189258 150198
rect 189828 150090 189856 154294
rect 190460 152924 190512 152930
rect 190460 152866 190512 152872
rect 190472 150090 190500 152866
rect 190564 152726 190592 163254
rect 190932 163146 190960 163254
rect 191010 163200 191066 164400
rect 191838 163200 191894 164400
rect 192666 163200 192722 164400
rect 193494 163200 193550 164400
rect 194322 163200 194378 164400
rect 195150 163200 195206 164400
rect 195978 163200 196034 164400
rect 196898 163200 196954 164400
rect 197726 163200 197782 164400
rect 198554 163200 198610 164400
rect 199382 163200 199438 164400
rect 200210 163200 200266 164400
rect 201038 163200 201094 164400
rect 201866 163200 201922 164400
rect 202694 163200 202750 164400
rect 203614 163200 203670 164400
rect 204442 163200 204498 164400
rect 204548 163254 205220 163282
rect 191024 163146 191052 163200
rect 190932 163118 191052 163146
rect 191104 157820 191156 157826
rect 191104 157762 191156 157768
rect 191012 156596 191064 156602
rect 191012 156538 191064 156544
rect 191024 156330 191052 156538
rect 191012 156324 191064 156330
rect 191012 156266 191064 156272
rect 191012 154284 191064 154290
rect 191012 154226 191064 154232
rect 191024 153542 191052 154226
rect 191012 153536 191064 153542
rect 191012 153478 191064 153484
rect 190552 152720 190604 152726
rect 190552 152662 190604 152668
rect 191116 150226 191144 157762
rect 191852 157350 191880 163200
rect 191840 157344 191892 157350
rect 191840 157286 191892 157292
rect 191196 156596 191248 156602
rect 191196 156538 191248 156544
rect 191208 156505 191236 156538
rect 191194 156496 191250 156505
rect 191194 156431 191250 156440
rect 192680 155106 192708 163200
rect 193508 159186 193536 163200
rect 194336 159934 194364 163200
rect 194324 159928 194376 159934
rect 194324 159870 194376 159876
rect 193496 159180 193548 159186
rect 193496 159122 193548 159128
rect 194508 158908 194560 158914
rect 194508 158850 194560 158856
rect 193680 156392 193732 156398
rect 193680 156334 193732 156340
rect 192392 155100 192444 155106
rect 192392 155042 192444 155048
rect 192668 155100 192720 155106
rect 192668 155042 192720 155048
rect 191748 154964 191800 154970
rect 191748 154906 191800 154912
rect 191196 154352 191248 154358
rect 191196 154294 191248 154300
rect 191208 153474 191236 154294
rect 191286 153640 191342 153649
rect 191286 153575 191288 153584
rect 191340 153575 191342 153584
rect 191288 153546 191340 153552
rect 191196 153468 191248 153474
rect 191196 153410 191248 153416
rect 191288 153468 191340 153474
rect 191288 153410 191340 153416
rect 191300 153377 191328 153410
rect 191286 153368 191342 153377
rect 191286 153303 191342 153312
rect 191116 150198 191190 150226
rect 189828 150062 189902 150090
rect 190472 150062 190546 150090
rect 189874 149940 189902 150062
rect 190518 149940 190546 150062
rect 191162 149940 191190 150198
rect 191760 150090 191788 154906
rect 192404 150090 192432 155042
rect 193036 152176 193088 152182
rect 193036 152118 193088 152124
rect 193048 150090 193076 152118
rect 193692 150090 193720 156334
rect 194324 154828 194376 154834
rect 194324 154770 194376 154776
rect 194336 150090 194364 154770
rect 194520 152930 194548 158850
rect 195164 157826 195192 163200
rect 195336 159316 195388 159322
rect 195336 159258 195388 159264
rect 195244 159248 195296 159254
rect 195244 159190 195296 159196
rect 195256 158982 195284 159190
rect 195244 158976 195296 158982
rect 195244 158918 195296 158924
rect 195348 158914 195376 159258
rect 195336 158908 195388 158914
rect 195336 158850 195388 158856
rect 195152 157820 195204 157826
rect 195152 157762 195204 157768
rect 195992 155038 196020 163200
rect 196164 160064 196216 160070
rect 196164 160006 196216 160012
rect 196072 158840 196124 158846
rect 196072 158782 196124 158788
rect 195980 155032 196032 155038
rect 195980 154974 196032 154980
rect 194968 153468 195020 153474
rect 194968 153410 195020 153416
rect 194508 152924 194560 152930
rect 194508 152866 194560 152872
rect 194980 150090 195008 153410
rect 196084 152998 196112 158782
rect 196176 153474 196204 160006
rect 196912 159254 196940 163200
rect 197636 159996 197688 160002
rect 197636 159938 197688 159944
rect 196900 159248 196952 159254
rect 196900 159190 196952 159196
rect 196254 158536 196310 158545
rect 196254 158471 196310 158480
rect 196164 153468 196216 153474
rect 196164 153410 196216 153416
rect 195612 152992 195664 152998
rect 195612 152934 195664 152940
rect 196072 152992 196124 152998
rect 196072 152934 196124 152940
rect 195624 150090 195652 152934
rect 196268 150226 196296 158471
rect 196900 153536 196952 153542
rect 196900 153478 196952 153484
rect 196268 150198 196342 150226
rect 191760 150062 191834 150090
rect 192404 150062 192478 150090
rect 193048 150062 193122 150090
rect 193692 150062 193766 150090
rect 194336 150062 194410 150090
rect 194980 150062 195054 150090
rect 195624 150062 195698 150090
rect 191806 149940 191834 150062
rect 192450 149940 192478 150062
rect 193094 149940 193122 150062
rect 193738 149940 193766 150062
rect 194382 149940 194410 150062
rect 195026 149940 195054 150062
rect 195670 149940 195698 150062
rect 196314 149940 196342 150198
rect 196912 150090 196940 153478
rect 197648 153270 197676 159938
rect 197740 159322 197768 163200
rect 197728 159316 197780 159322
rect 197728 159258 197780 159264
rect 198568 156534 198596 163200
rect 198740 158908 198792 158914
rect 198740 158850 198792 158856
rect 198556 156528 198608 156534
rect 198556 156470 198608 156476
rect 198752 153542 198780 158850
rect 198830 157176 198886 157185
rect 198830 157111 198886 157120
rect 198740 153536 198792 153542
rect 198740 153478 198792 153484
rect 197544 153264 197596 153270
rect 197544 153206 197596 153212
rect 197636 153264 197688 153270
rect 197636 153206 197688 153212
rect 197556 150090 197584 153206
rect 198188 152040 198240 152046
rect 198188 151982 198240 151988
rect 198200 150090 198228 151982
rect 198844 150090 198872 157111
rect 199396 154970 199424 163200
rect 200224 158846 200252 163200
rect 201052 160002 201080 163200
rect 201040 159996 201092 160002
rect 201040 159938 201092 159944
rect 200212 158840 200264 158846
rect 200212 158782 200264 158788
rect 200304 157684 200356 157690
rect 200304 157626 200356 157632
rect 200316 157554 200344 157626
rect 200580 157616 200632 157622
rect 200764 157616 200816 157622
rect 200632 157564 200764 157570
rect 200580 157558 200816 157564
rect 200212 157548 200264 157554
rect 200212 157490 200264 157496
rect 200304 157548 200356 157554
rect 200592 157542 200804 157558
rect 200304 157490 200356 157496
rect 199384 154964 199436 154970
rect 199384 154906 199436 154912
rect 199476 154284 199528 154290
rect 199476 154226 199528 154232
rect 199488 150090 199516 154226
rect 200118 153776 200174 153785
rect 200118 153711 200174 153720
rect 200132 150090 200160 153711
rect 200224 150210 200252 157490
rect 201880 156602 201908 163200
rect 202708 157334 202736 163200
rect 203628 158982 203656 163200
rect 203616 158976 203668 158982
rect 203616 158918 203668 158924
rect 204076 158908 204128 158914
rect 204076 158850 204128 158856
rect 202880 158772 202932 158778
rect 202880 158714 202932 158720
rect 202892 157690 202920 158714
rect 202880 157684 202932 157690
rect 202880 157626 202932 157632
rect 204088 157622 204116 158850
rect 204456 158778 204484 163200
rect 204444 158772 204496 158778
rect 204444 158714 204496 158720
rect 203984 157616 204036 157622
rect 203984 157558 204036 157564
rect 204076 157616 204128 157622
rect 204076 157558 204128 157564
rect 202708 157306 202828 157334
rect 200672 156596 200724 156602
rect 200672 156538 200724 156544
rect 201868 156596 201920 156602
rect 201868 156538 201920 156544
rect 200684 156194 200712 156538
rect 200856 156528 200908 156534
rect 200856 156470 200908 156476
rect 202696 156528 202748 156534
rect 202696 156470 202748 156476
rect 200672 156188 200724 156194
rect 200672 156130 200724 156136
rect 200764 156188 200816 156194
rect 200764 156130 200816 156136
rect 200776 156058 200804 156130
rect 200868 156058 200896 156470
rect 200764 156052 200816 156058
rect 200764 155994 200816 156000
rect 200856 156052 200908 156058
rect 200856 155994 200908 156000
rect 202052 154352 202104 154358
rect 202052 154294 202104 154300
rect 200764 153196 200816 153202
rect 200764 153138 200816 153144
rect 200212 150204 200264 150210
rect 200212 150146 200264 150152
rect 200776 150090 200804 153138
rect 201454 150204 201506 150210
rect 201454 150146 201506 150152
rect 196912 150062 196986 150090
rect 197556 150062 197630 150090
rect 198200 150062 198274 150090
rect 198844 150062 198918 150090
rect 199488 150062 199562 150090
rect 200132 150062 200206 150090
rect 200776 150062 200850 150090
rect 196958 149940 196986 150062
rect 197602 149940 197630 150062
rect 198246 149940 198274 150062
rect 198890 149940 198918 150062
rect 199534 149940 199562 150062
rect 200178 149940 200206 150062
rect 200822 149940 200850 150062
rect 201466 149940 201494 150146
rect 202064 150090 202092 154294
rect 202708 150090 202736 156470
rect 202800 154902 202828 157306
rect 202788 154896 202840 154902
rect 202788 154838 202840 154844
rect 203340 153060 203392 153066
rect 203340 153002 203392 153008
rect 203352 150090 203380 153002
rect 203996 150226 204024 157558
rect 204548 154290 204576 163254
rect 205192 163146 205220 163254
rect 205270 163200 205326 164400
rect 206098 163200 206154 164400
rect 206926 163200 206982 164400
rect 207754 163200 207810 164400
rect 208582 163200 208638 164400
rect 209410 163200 209466 164400
rect 210330 163200 210386 164400
rect 211158 163200 211214 164400
rect 211264 163254 211936 163282
rect 205284 163146 205312 163200
rect 205192 163118 205312 163146
rect 206112 156534 206140 163200
rect 206940 158914 206968 163200
rect 207768 160070 207796 163200
rect 207756 160064 207808 160070
rect 207756 160006 207808 160012
rect 206928 158908 206980 158914
rect 206928 158850 206980 158856
rect 206100 156528 206152 156534
rect 206100 156470 206152 156476
rect 207204 156460 207256 156466
rect 207204 156402 207256 156408
rect 206560 156256 206612 156262
rect 206560 156198 206612 156204
rect 204536 154284 204588 154290
rect 204536 154226 204588 154232
rect 204628 153400 204680 153406
rect 204628 153342 204680 153348
rect 203996 150198 204070 150226
rect 202064 150062 202138 150090
rect 202708 150062 202782 150090
rect 203352 150062 203426 150090
rect 202110 149940 202138 150062
rect 202754 149940 202782 150062
rect 203398 149940 203426 150062
rect 204042 149940 204070 150198
rect 204640 150090 204668 153342
rect 205272 153332 205324 153338
rect 205272 153274 205324 153280
rect 205284 150090 205312 153274
rect 205916 152312 205968 152318
rect 205916 152254 205968 152260
rect 205928 150226 205956 152254
rect 206572 150226 206600 156198
rect 207216 150226 207244 156402
rect 207848 154488 207900 154494
rect 207848 154430 207900 154436
rect 207860 150226 207888 154430
rect 208596 154358 208624 163200
rect 209136 157480 209188 157486
rect 209136 157422 209188 157428
rect 208584 154352 208636 154358
rect 208584 154294 208636 154300
rect 208492 153128 208544 153134
rect 208492 153070 208544 153076
rect 208504 150226 208532 153070
rect 209148 150226 209176 157422
rect 209424 156466 209452 163200
rect 210344 159050 210372 163200
rect 210240 159044 210292 159050
rect 210240 158986 210292 158992
rect 210332 159044 210384 159050
rect 210332 158986 210384 158992
rect 209412 156460 209464 156466
rect 209412 156402 209464 156408
rect 209780 154692 209832 154698
rect 209780 154634 209832 154640
rect 209792 150226 209820 154634
rect 210252 153066 210280 158986
rect 210516 154556 210568 154562
rect 210516 154498 210568 154504
rect 210240 153060 210292 153066
rect 210240 153002 210292 153008
rect 210528 150226 210556 154498
rect 211172 152930 211200 163200
rect 211264 154494 211292 163254
rect 211908 163146 211936 163254
rect 211986 163200 212042 164400
rect 212814 163200 212870 164400
rect 213642 163200 213698 164400
rect 214470 163200 214526 164400
rect 215298 163200 215354 164400
rect 216126 163200 216182 164400
rect 216692 163254 216996 163282
rect 212000 163146 212028 163200
rect 211908 163118 212028 163146
rect 211804 159248 211856 159254
rect 211804 159190 211856 159196
rect 211344 156664 211396 156670
rect 211344 156606 211396 156612
rect 211252 154488 211304 154494
rect 211252 154430 211304 154436
rect 211068 152924 211120 152930
rect 211068 152866 211120 152872
rect 211160 152924 211212 152930
rect 211160 152866 211212 152872
rect 205928 150198 206002 150226
rect 206572 150198 206646 150226
rect 207216 150198 207290 150226
rect 207860 150198 207934 150226
rect 208504 150198 208578 150226
rect 209148 150198 209222 150226
rect 209792 150198 209866 150226
rect 204640 150062 204714 150090
rect 205284 150062 205358 150090
rect 204686 149940 204714 150062
rect 205330 149940 205358 150062
rect 205974 149940 206002 150198
rect 206618 149940 206646 150198
rect 207262 149940 207290 150198
rect 207906 149940 207934 150198
rect 208550 149940 208578 150198
rect 209194 149940 209222 150198
rect 209838 149940 209866 150198
rect 210482 150198 210556 150226
rect 211080 150226 211108 152866
rect 211356 151814 211384 156606
rect 211816 156262 211844 159190
rect 211804 156256 211856 156262
rect 211804 156198 211856 156204
rect 212828 154698 212856 163200
rect 213656 159254 213684 163200
rect 214484 159322 214512 163200
rect 214380 159316 214432 159322
rect 214380 159258 214432 159264
rect 214472 159316 214524 159322
rect 214472 159258 214524 159264
rect 213644 159248 213696 159254
rect 213644 159190 213696 159196
rect 214392 159050 214420 159258
rect 214564 159112 214616 159118
rect 214564 159054 214616 159060
rect 214012 159044 214064 159050
rect 214012 158986 214064 158992
rect 214380 159044 214432 159050
rect 214380 158986 214432 158992
rect 213920 156188 213972 156194
rect 213920 156130 213972 156136
rect 212816 154692 212868 154698
rect 212816 154634 212868 154640
rect 212264 154624 212316 154630
rect 212264 154566 212316 154572
rect 211356 151786 211660 151814
rect 211632 150226 211660 151786
rect 212276 150226 212304 154566
rect 212908 153808 212960 153814
rect 212908 153750 212960 153756
rect 212920 150226 212948 153750
rect 213552 152108 213604 152114
rect 213552 152050 213604 152056
rect 213564 150226 213592 152050
rect 211080 150198 211154 150226
rect 211632 150198 211706 150226
rect 212276 150198 212350 150226
rect 212920 150198 212994 150226
rect 213564 150198 213638 150226
rect 213932 150210 213960 156130
rect 214024 153134 214052 158986
rect 214576 156126 214604 159054
rect 214196 156120 214248 156126
rect 214196 156062 214248 156068
rect 214564 156120 214616 156126
rect 214564 156062 214616 156068
rect 214012 153128 214064 153134
rect 214012 153070 214064 153076
rect 214208 150226 214236 156062
rect 215312 154562 215340 163200
rect 215392 159044 215444 159050
rect 215392 158986 215444 158992
rect 215300 154556 215352 154562
rect 215300 154498 215352 154504
rect 215404 151842 215432 158986
rect 216140 156670 216168 163200
rect 216128 156664 216180 156670
rect 216128 156606 216180 156612
rect 215484 153876 215536 153882
rect 215484 153818 215536 153824
rect 215392 151836 215444 151842
rect 215392 151778 215444 151784
rect 215496 150226 215524 153818
rect 216692 152998 216720 163254
rect 216968 163146 216996 163254
rect 217046 163200 217102 164400
rect 217152 163254 217824 163282
rect 217060 163146 217088 163200
rect 216968 163118 217088 163146
rect 216864 156800 216916 156806
rect 216864 156742 216916 156748
rect 216128 152992 216180 152998
rect 216128 152934 216180 152940
rect 216680 152992 216732 152998
rect 216680 152934 216732 152940
rect 216140 150226 216168 152934
rect 216876 150226 216904 156742
rect 217152 152425 217180 163254
rect 217796 163146 217824 163254
rect 217874 163200 217930 164400
rect 218072 163254 218652 163282
rect 217888 163146 217916 163200
rect 217796 163118 217916 163146
rect 217416 155236 217468 155242
rect 217416 155178 217468 155184
rect 217138 152416 217194 152425
rect 217138 152351 217194 152360
rect 210482 149940 210510 150198
rect 211126 149940 211154 150198
rect 211678 149940 211706 150198
rect 212322 149940 212350 150198
rect 212966 149940 212994 150198
rect 213610 149940 213638 150198
rect 213920 150204 213972 150210
rect 214208 150198 214282 150226
rect 213920 150146 213972 150152
rect 214254 149940 214282 150198
rect 214886 150204 214938 150210
rect 215496 150198 215570 150226
rect 216140 150198 216214 150226
rect 214886 150146 214938 150152
rect 214898 149940 214926 150146
rect 215542 149940 215570 150198
rect 216186 149940 216214 150198
rect 216830 150198 216904 150226
rect 217428 150226 217456 155178
rect 218072 153882 218100 163254
rect 218624 163146 218652 163254
rect 218702 163200 218758 164400
rect 219530 163200 219586 164400
rect 220358 163200 220414 164400
rect 221186 163200 221242 164400
rect 221292 163254 221964 163282
rect 218716 163146 218744 163200
rect 218624 163118 218744 163146
rect 218152 159588 218204 159594
rect 218152 159530 218204 159536
rect 218060 153876 218112 153882
rect 218060 153818 218112 153824
rect 218060 153740 218112 153746
rect 218060 153682 218112 153688
rect 218072 150226 218100 153682
rect 218164 153202 218192 159530
rect 219544 156806 219572 163200
rect 220372 159118 220400 163200
rect 221200 159594 221228 163200
rect 221188 159588 221240 159594
rect 221188 159530 221240 159536
rect 220360 159112 220412 159118
rect 220360 159054 220412 159060
rect 219900 158772 219952 158778
rect 219900 158714 219952 158720
rect 219532 156800 219584 156806
rect 219532 156742 219584 156748
rect 218244 155984 218296 155990
rect 218244 155926 218296 155932
rect 218152 153196 218204 153202
rect 218152 153138 218204 153144
rect 217428 150198 217502 150226
rect 218072 150198 218146 150226
rect 218256 150210 218284 155926
rect 219532 155304 219584 155310
rect 219532 155246 219584 155252
rect 218704 152516 218756 152522
rect 218704 152458 218756 152464
rect 218716 150226 218744 152458
rect 219544 151814 219572 155246
rect 219912 151910 219940 158714
rect 219992 157276 220044 157282
rect 219992 157218 220044 157224
rect 219900 151904 219952 151910
rect 219900 151846 219952 151852
rect 220004 151814 220032 157218
rect 221292 153785 221320 163254
rect 221936 163146 221964 163254
rect 222014 163200 222070 164400
rect 222842 163200 222898 164400
rect 223762 163200 223818 164400
rect 224590 163200 224646 164400
rect 224972 163254 225368 163282
rect 222028 163146 222056 163200
rect 221936 163118 222056 163146
rect 221924 158024 221976 158030
rect 221924 157966 221976 157972
rect 221278 153776 221334 153785
rect 221278 153711 221334 153720
rect 221280 153060 221332 153066
rect 221280 153002 221332 153008
rect 219544 151786 219940 151814
rect 220004 151786 220676 151814
rect 219912 150498 219940 151786
rect 219912 150470 220032 150498
rect 220004 150226 220032 150470
rect 220648 150226 220676 151786
rect 221292 150226 221320 153002
rect 221936 150226 221964 157966
rect 222856 156874 222884 163200
rect 223580 159180 223632 159186
rect 223580 159122 223632 159128
rect 222568 156868 222620 156874
rect 222568 156810 222620 156816
rect 222844 156868 222896 156874
rect 222844 156810 222896 156816
rect 222580 150226 222608 156810
rect 223592 156126 223620 159122
rect 223580 156120 223632 156126
rect 223580 156062 223632 156068
rect 223212 153672 223264 153678
rect 223212 153614 223264 153620
rect 223224 150226 223252 153614
rect 223776 152522 223804 163200
rect 224224 159044 224276 159050
rect 224224 158986 224276 158992
rect 224236 158846 224264 158986
rect 224604 158846 224632 163200
rect 224224 158840 224276 158846
rect 224224 158782 224276 158788
rect 224592 158840 224644 158846
rect 224592 158782 224644 158788
rect 224500 156936 224552 156942
rect 224500 156878 224552 156884
rect 223764 152516 223816 152522
rect 223764 152458 223816 152464
rect 223856 151972 223908 151978
rect 223856 151914 223908 151920
rect 223868 150226 223896 151914
rect 224512 150226 224540 156878
rect 224972 153814 225000 163254
rect 225340 163146 225368 163254
rect 225418 163200 225474 164400
rect 226246 163200 226302 164400
rect 227074 163200 227130 164400
rect 227902 163200 227958 164400
rect 228008 163254 228680 163282
rect 225432 163146 225460 163200
rect 225340 163118 225460 163146
rect 225144 156732 225196 156738
rect 225144 156674 225196 156680
rect 224960 153808 225012 153814
rect 224960 153750 225012 153756
rect 216830 149940 216858 150198
rect 217474 149940 217502 150198
rect 218118 149940 218146 150198
rect 218244 150204 218296 150210
rect 218716 150198 218790 150226
rect 218244 150146 218296 150152
rect 218762 149940 218790 150198
rect 219394 150204 219446 150210
rect 220004 150198 220078 150226
rect 220648 150198 220722 150226
rect 221292 150198 221366 150226
rect 221936 150198 222010 150226
rect 222580 150198 222654 150226
rect 223224 150198 223298 150226
rect 223868 150198 223942 150226
rect 224512 150198 224586 150226
rect 219394 150146 219446 150152
rect 219406 149940 219434 150146
rect 220050 149940 220078 150198
rect 220694 149940 220722 150198
rect 221338 149940 221366 150198
rect 221982 149940 222010 150198
rect 222626 149940 222654 150198
rect 223270 149940 223298 150198
rect 223914 149940 223942 150198
rect 224558 149940 224586 150198
rect 225156 150090 225184 156674
rect 226260 156398 226288 163200
rect 226340 159520 226392 159526
rect 226340 159462 226392 159468
rect 225788 156392 225840 156398
rect 225788 156334 225840 156340
rect 226248 156392 226300 156398
rect 226248 156334 226300 156340
rect 225800 150090 225828 156334
rect 226352 153202 226380 159462
rect 227088 158778 227116 163200
rect 227916 159526 227944 163200
rect 227904 159520 227956 159526
rect 227904 159462 227956 159468
rect 227720 159044 227772 159050
rect 227720 158986 227772 158992
rect 227076 158772 227128 158778
rect 227076 158714 227128 158720
rect 226892 157412 226944 157418
rect 226892 157354 226944 157360
rect 226248 153196 226300 153202
rect 226248 153138 226300 153144
rect 226340 153196 226392 153202
rect 226340 153138 226392 153144
rect 226260 153082 226288 153138
rect 226260 153054 226472 153082
rect 226444 150226 226472 153054
rect 226904 150226 226932 157354
rect 227732 154630 227760 158986
rect 227812 157072 227864 157078
rect 227812 157014 227864 157020
rect 227720 154624 227772 154630
rect 227720 154566 227772 154572
rect 226444 150198 226518 150226
rect 226904 150198 227162 150226
rect 225156 150062 225230 150090
rect 225800 150062 225874 150090
rect 225202 149940 225230 150062
rect 225846 149940 225874 150062
rect 226490 149940 226518 150198
rect 227134 149940 227162 150198
rect 227824 150090 227852 157014
rect 228008 153746 228036 163254
rect 228652 163146 228680 163254
rect 228730 163200 228786 164400
rect 229650 163200 229706 164400
rect 230478 163200 230534 164400
rect 230584 163254 231256 163282
rect 228744 163146 228772 163200
rect 228652 163118 228772 163146
rect 229376 159112 229428 159118
rect 229376 159054 229428 159060
rect 228364 154828 228416 154834
rect 228364 154770 228416 154776
rect 227996 153740 228048 153746
rect 227996 153682 228048 153688
rect 227778 150062 227852 150090
rect 228376 150090 228404 154770
rect 229008 152244 229060 152250
rect 229008 152186 229060 152192
rect 229020 150090 229048 152186
rect 229388 152182 229416 159054
rect 229560 157004 229612 157010
rect 229560 156946 229612 156952
rect 229376 152176 229428 152182
rect 229376 152118 229428 152124
rect 229572 150226 229600 156946
rect 229664 156942 229692 163200
rect 230492 159118 230520 163200
rect 230480 159112 230532 159118
rect 230480 159054 230532 159060
rect 229652 156936 229704 156942
rect 229652 156878 229704 156884
rect 229652 154760 229704 154766
rect 229836 154760 229888 154766
rect 229704 154708 229836 154714
rect 229652 154702 229888 154708
rect 229664 154686 229876 154702
rect 230296 153944 230348 153950
rect 230296 153886 230348 153892
rect 229572 150198 229738 150226
rect 228376 150062 228450 150090
rect 229020 150062 229094 150090
rect 227778 149940 227806 150062
rect 228422 149940 228450 150062
rect 229066 149940 229094 150062
rect 229710 149940 229738 150198
rect 230308 150090 230336 153886
rect 230584 153066 230612 163254
rect 231228 163146 231256 163254
rect 231306 163200 231362 164400
rect 231872 163254 232084 163282
rect 231320 163146 231348 163200
rect 231228 163118 231348 163146
rect 230756 158840 230808 158846
rect 230756 158782 230808 158788
rect 230572 153060 230624 153066
rect 230572 153002 230624 153008
rect 230768 152318 230796 158782
rect 231872 154018 231900 163254
rect 232056 163146 232084 163254
rect 232134 163200 232190 164400
rect 232962 163200 233018 164400
rect 233790 163200 233846 164400
rect 234618 163200 234674 164400
rect 234724 163254 235396 163282
rect 232148 163146 232176 163200
rect 232056 163118 232176 163146
rect 231952 158092 232004 158098
rect 231952 158034 232004 158040
rect 231964 157334 231992 158034
rect 231964 157306 232268 157334
rect 230940 154012 230992 154018
rect 230940 153954 230992 153960
rect 231860 154012 231912 154018
rect 231860 153954 231912 153960
rect 230756 152312 230808 152318
rect 230756 152254 230808 152260
rect 230952 150090 230980 153954
rect 231584 153196 231636 153202
rect 231584 153138 231636 153144
rect 231596 150090 231624 153138
rect 232240 150226 232268 157306
rect 232976 157010 233004 163200
rect 233804 159050 233832 163200
rect 234632 159186 234660 163200
rect 234620 159180 234672 159186
rect 234620 159122 234672 159128
rect 233792 159044 233844 159050
rect 233792 158986 233844 158992
rect 233148 158976 233200 158982
rect 233148 158918 233200 158924
rect 233160 157486 233188 158918
rect 233884 158908 233936 158914
rect 233884 158850 233936 158856
rect 233516 157548 233568 157554
rect 233516 157490 233568 157496
rect 233148 157480 233200 157486
rect 233148 157422 233200 157428
rect 232964 157004 233016 157010
rect 232964 156946 233016 156952
rect 232872 155372 232924 155378
rect 232872 155314 232924 155320
rect 232240 150198 232314 150226
rect 230308 150062 230382 150090
rect 230952 150062 231026 150090
rect 231596 150062 231670 150090
rect 230354 149940 230382 150062
rect 230998 149940 231026 150062
rect 231642 149940 231670 150062
rect 232286 149940 232314 150198
rect 232884 150090 232912 155314
rect 233528 150226 233556 157490
rect 233896 155242 233924 158850
rect 233884 155236 233936 155242
rect 233884 155178 233936 155184
rect 234724 153950 234752 163254
rect 235368 163146 235396 163254
rect 235446 163200 235502 164400
rect 236366 163200 236422 164400
rect 237194 163200 237250 164400
rect 237392 163254 237972 163282
rect 235460 163146 235488 163200
rect 235368 163118 235488 163146
rect 236380 158030 236408 163200
rect 236736 159384 236788 159390
rect 236736 159326 236788 159332
rect 236368 158024 236420 158030
rect 236368 157966 236420 157972
rect 234804 157140 234856 157146
rect 234804 157082 234856 157088
rect 234712 153944 234764 153950
rect 234712 153886 234764 153892
rect 234160 152788 234212 152794
rect 234160 152730 234212 152736
rect 233528 150198 233602 150226
rect 232884 150062 232958 150090
rect 232930 149940 232958 150062
rect 233574 149940 233602 150198
rect 234172 150090 234200 152730
rect 234816 150226 234844 157082
rect 235448 154080 235500 154086
rect 235448 154022 235500 154028
rect 235460 150226 235488 154022
rect 236092 153604 236144 153610
rect 236092 153546 236144 153552
rect 236104 150226 236132 153546
rect 236748 150226 236776 159326
rect 237208 153202 237236 163200
rect 237196 153196 237248 153202
rect 237196 153138 237248 153144
rect 237392 152794 237420 163254
rect 237944 163146 237972 163254
rect 238022 163200 238078 164400
rect 238850 163200 238906 164400
rect 239678 163200 239734 164400
rect 240506 163200 240562 164400
rect 241334 163200 241390 164400
rect 241532 163254 242112 163282
rect 238036 163146 238064 163200
rect 237944 163118 238064 163146
rect 238864 161474 238892 163200
rect 238864 161446 238984 161474
rect 237472 158228 237524 158234
rect 237472 158170 237524 158176
rect 237380 152788 237432 152794
rect 237380 152730 237432 152736
rect 237484 150226 237512 158170
rect 238852 158160 238904 158166
rect 238852 158102 238904 158108
rect 238668 156324 238720 156330
rect 238668 156266 238720 156272
rect 237564 155440 237616 155446
rect 237564 155382 237616 155388
rect 237576 151814 237604 155382
rect 237576 151786 238064 151814
rect 234816 150198 234890 150226
rect 235460 150198 235534 150226
rect 236104 150198 236178 150226
rect 236748 150198 236822 150226
rect 234172 150062 234246 150090
rect 234218 149940 234246 150062
rect 234862 149940 234890 150198
rect 235506 149940 235534 150198
rect 236150 149940 236178 150198
rect 236794 149940 236822 150198
rect 237438 150198 237512 150226
rect 238036 150226 238064 151786
rect 238680 150226 238708 156266
rect 238036 150198 238110 150226
rect 238680 150198 238754 150226
rect 238864 150210 238892 158102
rect 238956 153610 238984 161446
rect 239692 158098 239720 163200
rect 240324 159452 240376 159458
rect 240324 159394 240376 159400
rect 239680 158092 239732 158098
rect 239680 158034 239732 158040
rect 238944 153604 238996 153610
rect 238944 153546 238996 153552
rect 240336 152590 240364 159394
rect 240520 158982 240548 163200
rect 241348 159390 241376 163200
rect 241336 159384 241388 159390
rect 241336 159326 241388 159332
rect 240508 158976 240560 158982
rect 240508 158918 240560 158924
rect 241428 158772 241480 158778
rect 241428 158714 241480 158720
rect 240600 155576 240652 155582
rect 240600 155518 240652 155524
rect 239312 152584 239364 152590
rect 239312 152526 239364 152532
rect 240324 152584 240376 152590
rect 240324 152526 240376 152532
rect 239324 150226 239352 152526
rect 240612 150226 240640 155518
rect 241440 154698 241468 158714
rect 241428 154692 241480 154698
rect 241428 154634 241480 154640
rect 241532 153678 241560 163254
rect 242084 163146 242112 163254
rect 242162 163200 242218 164400
rect 243082 163200 243138 164400
rect 243910 163200 243966 164400
rect 244738 163200 244794 164400
rect 245566 163200 245622 164400
rect 246394 163200 246450 164400
rect 247222 163200 247278 164400
rect 248050 163200 248106 164400
rect 248432 163254 248828 163282
rect 242176 163146 242204 163200
rect 242084 163118 242204 163146
rect 243096 161474 243124 163200
rect 243096 161446 243216 161474
rect 242992 159724 243044 159730
rect 242992 159666 243044 159672
rect 242440 158500 242492 158506
rect 242440 158442 242492 158448
rect 241520 153672 241572 153678
rect 241520 153614 241572 153620
rect 241244 153468 241296 153474
rect 241244 153410 241296 153416
rect 241256 150226 241284 153410
rect 241888 152584 241940 152590
rect 241888 152526 241940 152532
rect 241900 150226 241928 152526
rect 242452 150226 242480 158442
rect 242900 154760 242952 154766
rect 242900 154702 242952 154708
rect 237438 149940 237466 150198
rect 238082 149940 238110 150198
rect 238726 149940 238754 150198
rect 238852 150204 238904 150210
rect 239324 150198 239398 150226
rect 238852 150146 238904 150152
rect 239370 149940 239398 150198
rect 240002 150204 240054 150210
rect 240612 150198 240686 150226
rect 241256 150198 241330 150226
rect 241900 150198 241974 150226
rect 242452 150198 242526 150226
rect 242912 150210 242940 154702
rect 243004 152590 243032 159666
rect 243084 155508 243136 155514
rect 243084 155450 243136 155456
rect 242992 152584 243044 152590
rect 242992 152526 243044 152532
rect 243096 150226 243124 155450
rect 243188 155310 243216 161446
rect 243924 158846 243952 163200
rect 243912 158840 243964 158846
rect 243912 158782 243964 158788
rect 244752 158778 244780 163200
rect 244740 158772 244792 158778
rect 244740 158714 244792 158720
rect 245016 158296 245068 158302
rect 245016 158238 245068 158244
rect 243176 155304 243228 155310
rect 243176 155246 243228 155252
rect 243544 155236 243596 155242
rect 243544 155178 243596 155184
rect 243556 154766 243584 155178
rect 243544 154760 243596 154766
rect 243544 154702 243596 154708
rect 244372 152652 244424 152658
rect 244372 152594 244424 152600
rect 244384 150226 244412 152594
rect 245028 150226 245056 158238
rect 245580 154086 245608 163200
rect 246120 158840 246172 158846
rect 246120 158782 246172 158788
rect 245752 158772 245804 158778
rect 245752 158714 245804 158720
rect 245660 154148 245712 154154
rect 245660 154090 245712 154096
rect 245568 154080 245620 154086
rect 245568 154022 245620 154028
rect 245672 150226 245700 154090
rect 245764 152658 245792 158714
rect 245752 152652 245804 152658
rect 245752 152594 245804 152600
rect 246132 152250 246160 158782
rect 246408 158166 246436 163200
rect 247236 159458 247264 163200
rect 248064 159730 248092 163200
rect 248052 159724 248104 159730
rect 248052 159666 248104 159672
rect 247224 159452 247276 159458
rect 247224 159394 247276 159400
rect 247592 158432 247644 158438
rect 247592 158374 247644 158380
rect 246396 158160 246448 158166
rect 246396 158102 246448 158108
rect 247132 155644 247184 155650
rect 247132 155586 247184 155592
rect 246304 153264 246356 153270
rect 246304 153206 246356 153212
rect 246120 152244 246172 152250
rect 246120 152186 246172 152192
rect 246316 150226 246344 153206
rect 246948 152584 247000 152590
rect 246948 152526 247000 152532
rect 246960 150226 246988 152526
rect 240002 150146 240054 150152
rect 240014 149940 240042 150146
rect 240658 149940 240686 150198
rect 241302 149940 241330 150198
rect 241946 149940 241974 150198
rect 242498 149940 242526 150198
rect 242900 150204 242952 150210
rect 243096 150198 243170 150226
rect 242900 150146 242952 150152
rect 243142 149940 243170 150198
rect 243774 150204 243826 150210
rect 244384 150198 244458 150226
rect 245028 150198 245102 150226
rect 245672 150198 245746 150226
rect 246316 150198 246390 150226
rect 246960 150198 247034 150226
rect 247144 150210 247172 155586
rect 247604 150226 247632 158374
rect 248432 154154 248460 163254
rect 248800 163146 248828 163254
rect 248878 163200 248934 164400
rect 249798 163200 249854 164400
rect 249996 163254 250576 163282
rect 248892 163146 248920 163200
rect 248800 163118 248920 163146
rect 249812 158234 249840 163200
rect 249892 158364 249944 158370
rect 249892 158306 249944 158312
rect 249800 158228 249852 158234
rect 249800 158170 249852 158176
rect 248420 154148 248472 154154
rect 248420 154090 248472 154096
rect 248880 153536 248932 153542
rect 248880 153478 248932 153484
rect 248892 150226 248920 153478
rect 249524 152856 249576 152862
rect 249524 152798 249576 152804
rect 249536 150226 249564 152798
rect 249904 151814 249932 158306
rect 249996 152590 250024 163254
rect 250548 163146 250576 163254
rect 250626 163200 250682 164400
rect 251454 163200 251510 164400
rect 251560 163254 252232 163282
rect 250640 163146 250668 163200
rect 250548 163118 250668 163146
rect 251180 159656 251232 159662
rect 251180 159598 251232 159604
rect 250812 155712 250864 155718
rect 250812 155654 250864 155660
rect 249984 152584 250036 152590
rect 249984 152526 250036 152532
rect 249904 151786 250208 151814
rect 250180 150226 250208 151786
rect 250824 150226 250852 155654
rect 243774 150146 243826 150152
rect 243786 149940 243814 150146
rect 244430 149940 244458 150198
rect 245074 149940 245102 150198
rect 245718 149940 245746 150198
rect 246362 149940 246390 150198
rect 247006 149940 247034 150198
rect 247132 150204 247184 150210
rect 247604 150198 247678 150226
rect 247132 150146 247184 150152
rect 247650 149940 247678 150198
rect 248282 150204 248334 150210
rect 248892 150198 248966 150226
rect 249536 150198 249610 150226
rect 250180 150198 250254 150226
rect 250824 150198 250898 150226
rect 251192 150210 251220 159598
rect 251468 158778 251496 163200
rect 251456 158772 251508 158778
rect 251456 158714 251508 158720
rect 251456 157616 251508 157622
rect 251456 157558 251508 157564
rect 251468 150226 251496 157558
rect 251560 153542 251588 163254
rect 252204 163146 252232 163254
rect 252282 163200 252338 164400
rect 253110 163200 253166 164400
rect 253938 163200 253994 164400
rect 254766 163200 254822 164400
rect 255332 163254 255544 163282
rect 252296 163146 252324 163200
rect 252204 163118 252324 163146
rect 252928 158772 252980 158778
rect 252928 158714 252980 158720
rect 252744 158636 252796 158642
rect 252744 158578 252796 158584
rect 251548 153536 251600 153542
rect 251548 153478 251600 153484
rect 252756 150226 252784 158578
rect 252940 152114 252968 158714
rect 253124 155310 253152 163200
rect 253952 158914 253980 163200
rect 254780 159662 254808 163200
rect 254768 159656 254820 159662
rect 254768 159598 254820 159604
rect 253940 158908 253992 158914
rect 253940 158850 253992 158856
rect 253112 155304 253164 155310
rect 253112 155246 253164 155252
rect 254032 154420 254084 154426
rect 254032 154362 254084 154368
rect 253388 154216 253440 154222
rect 253388 154158 253440 154164
rect 252928 152108 252980 152114
rect 252928 152050 252980 152056
rect 253400 150226 253428 154158
rect 254044 150226 254072 154362
rect 255332 154222 255360 163254
rect 255516 163146 255544 163254
rect 255594 163200 255650 164400
rect 256514 163200 256570 164400
rect 256712 163254 257292 163282
rect 255608 163146 255636 163200
rect 255516 163118 255636 163146
rect 255504 159860 255556 159866
rect 255504 159802 255556 159808
rect 255412 158568 255464 158574
rect 255412 158510 255464 158516
rect 255320 154216 255372 154222
rect 255320 154158 255372 154164
rect 254676 152448 254728 152454
rect 254676 152390 254728 152396
rect 254688 150226 254716 152390
rect 255424 150226 255452 158510
rect 255516 152862 255544 159802
rect 255872 157684 255924 157690
rect 255872 157626 255924 157632
rect 255688 155916 255740 155922
rect 255688 155858 255740 155864
rect 255504 152856 255556 152862
rect 255504 152798 255556 152804
rect 255700 151814 255728 155858
rect 255884 151814 255912 157626
rect 256528 155378 256556 163200
rect 256516 155372 256568 155378
rect 256516 155314 256568 155320
rect 256712 152454 256740 163254
rect 257264 163146 257292 163254
rect 257342 163200 257398 164400
rect 258170 163200 258226 164400
rect 258276 163254 258948 163282
rect 257356 163146 257384 163200
rect 257264 163118 257384 163146
rect 258184 161474 258212 163200
rect 258092 161446 258212 161474
rect 256792 158704 256844 158710
rect 256792 158646 256844 158652
rect 256700 152448 256752 152454
rect 256700 152390 256752 152396
rect 255700 151786 255820 151814
rect 255884 151786 256648 151814
rect 248282 150146 248334 150152
rect 248294 149940 248322 150146
rect 248938 149940 248966 150198
rect 249582 149940 249610 150198
rect 250226 149940 250254 150198
rect 250870 149940 250898 150198
rect 251180 150204 251232 150210
rect 251468 150198 251542 150226
rect 251180 150146 251232 150152
rect 251514 149940 251542 150198
rect 252146 150204 252198 150210
rect 252756 150198 252830 150226
rect 253400 150198 253474 150226
rect 254044 150198 254118 150226
rect 254688 150198 254762 150226
rect 252146 150146 252198 150152
rect 252158 149940 252186 150146
rect 252802 149940 252830 150198
rect 253446 149940 253474 150198
rect 254090 149940 254118 150198
rect 254734 149940 254762 150198
rect 255378 150198 255452 150226
rect 255792 150226 255820 151786
rect 256620 150226 256648 151786
rect 255792 150198 256050 150226
rect 256620 150198 256694 150226
rect 256804 150210 256832 158646
rect 258092 152862 258120 161446
rect 258172 157208 258224 157214
rect 258172 157150 258224 157156
rect 257252 152856 257304 152862
rect 257252 152798 257304 152804
rect 258080 152856 258132 152862
rect 258080 152798 258132 152804
rect 257264 150226 257292 152798
rect 255378 149940 255406 150198
rect 256022 149940 256050 150198
rect 256666 149940 256694 150198
rect 256792 150204 256844 150210
rect 257264 150198 257338 150226
rect 258184 150210 258212 157150
rect 258276 154426 258304 163254
rect 258920 163146 258948 163254
rect 258998 163200 259054 164400
rect 259826 163200 259882 164400
rect 260654 163200 260710 164400
rect 261482 163200 261538 164400
rect 262402 163200 262458 164400
rect 263230 163200 263286 164400
rect 263612 163254 264008 163282
rect 259012 163146 259040 163200
rect 258920 163118 259040 163146
rect 258540 155780 258592 155786
rect 258540 155722 258592 155728
rect 258264 154420 258316 154426
rect 258264 154362 258316 154368
rect 258552 150226 258580 155722
rect 259840 155446 259868 163200
rect 260668 159866 260696 163200
rect 260656 159860 260708 159866
rect 260656 159802 260708 159808
rect 261496 158846 261524 163200
rect 262220 159792 262272 159798
rect 262220 159734 262272 159740
rect 261484 158840 261536 158846
rect 261484 158782 261536 158788
rect 260472 157752 260524 157758
rect 260472 157694 260524 157700
rect 259828 155440 259880 155446
rect 259828 155382 259880 155388
rect 259828 152380 259880 152386
rect 259828 152322 259880 152328
rect 259840 150226 259868 152322
rect 260484 150226 260512 157694
rect 260840 156188 260892 156194
rect 260840 156130 260892 156136
rect 256792 150146 256844 150152
rect 257310 149940 257338 150198
rect 257942 150204 257994 150210
rect 257942 150146 257994 150152
rect 258172 150204 258224 150210
rect 258552 150198 258626 150226
rect 258172 150146 258224 150152
rect 257954 149940 257982 150146
rect 258598 149940 258626 150198
rect 259230 150204 259282 150210
rect 259840 150198 259914 150226
rect 260484 150198 260558 150226
rect 260852 150210 260880 156130
rect 261116 155848 261168 155854
rect 261116 155790 261168 155796
rect 261128 150226 261156 155790
rect 262232 151814 262260 159734
rect 262416 153406 262444 163200
rect 263048 157956 263100 157962
rect 263048 157898 263100 157904
rect 262404 153400 262456 153406
rect 262404 153342 262456 153348
rect 262232 151786 262444 151814
rect 262416 150226 262444 151786
rect 263060 150226 263088 157898
rect 263244 155514 263272 163200
rect 263232 155508 263284 155514
rect 263232 155450 263284 155456
rect 263612 152386 263640 163254
rect 263980 163146 264008 163254
rect 264058 163200 264114 164400
rect 264164 163254 264836 163282
rect 264072 163146 264100 163200
rect 263980 163118 264100 163146
rect 263784 155168 263836 155174
rect 263784 155110 263836 155116
rect 263600 152380 263652 152386
rect 263600 152322 263652 152328
rect 263796 150226 263824 155110
rect 264164 152046 264192 163254
rect 264808 163146 264836 163254
rect 264886 163200 264942 164400
rect 264992 163254 265664 163282
rect 264900 163146 264928 163200
rect 264808 163118 264928 163146
rect 264336 157888 264388 157894
rect 264336 157830 264388 157836
rect 264152 152040 264204 152046
rect 264152 151982 264204 151988
rect 259230 150146 259282 150152
rect 259242 149940 259270 150146
rect 259886 149940 259914 150198
rect 260530 149940 260558 150198
rect 260840 150204 260892 150210
rect 261128 150198 261202 150226
rect 260840 150146 260892 150152
rect 261174 149940 261202 150198
rect 261806 150204 261858 150210
rect 262416 150198 262490 150226
rect 263060 150198 263134 150226
rect 261806 150146 261858 150152
rect 261818 149940 261846 150146
rect 262462 149940 262490 150198
rect 263106 149940 263134 150198
rect 263750 150198 263824 150226
rect 264348 150226 264376 157830
rect 264992 153474 265020 163254
rect 265636 163146 265664 163254
rect 265714 163200 265770 164400
rect 266542 163200 266598 164400
rect 267370 163200 267426 164400
rect 268198 163200 268254 164400
rect 269118 163200 269174 164400
rect 269946 163200 270002 164400
rect 270774 163200 270830 164400
rect 270880 163254 271552 163282
rect 265728 163146 265756 163200
rect 265636 163118 265756 163146
rect 265164 157344 265216 157350
rect 265164 157286 265216 157292
rect 264980 153468 265032 153474
rect 264980 153410 265032 153416
rect 264980 152720 265032 152726
rect 264980 152662 265032 152668
rect 264992 150226 265020 152662
rect 265176 151814 265204 157286
rect 266452 156120 266504 156126
rect 266452 156062 266504 156068
rect 266268 155100 266320 155106
rect 266268 155042 266320 155048
rect 265176 151786 265664 151814
rect 265636 150226 265664 151786
rect 266280 150226 266308 155042
rect 266464 151814 266492 156062
rect 266556 155582 266584 163200
rect 267384 159798 267412 163200
rect 267556 159928 267608 159934
rect 267556 159870 267608 159876
rect 267372 159792 267424 159798
rect 267372 159734 267424 159740
rect 266544 155576 266596 155582
rect 266544 155518 266596 155524
rect 266464 151786 266952 151814
rect 266924 150226 266952 151786
rect 267568 150226 267596 159870
rect 268212 158778 268240 163200
rect 268200 158772 268252 158778
rect 268200 158714 268252 158720
rect 267740 157820 267792 157826
rect 267740 157762 267792 157768
rect 267752 151814 267780 157762
rect 268844 155032 268896 155038
rect 268844 154974 268896 154980
rect 267752 151786 268240 151814
rect 268212 150226 268240 151786
rect 268856 150226 268884 154974
rect 269132 153338 269160 163200
rect 269488 156256 269540 156262
rect 269488 156198 269540 156204
rect 269120 153332 269172 153338
rect 269120 153274 269172 153280
rect 269500 150226 269528 156198
rect 269960 155650 269988 163200
rect 270788 159934 270816 163200
rect 270776 159928 270828 159934
rect 270776 159870 270828 159876
rect 270592 156052 270644 156058
rect 270592 155994 270644 156000
rect 269948 155644 270000 155650
rect 269948 155586 270000 155592
rect 270132 151836 270184 151842
rect 270604 151814 270632 155994
rect 270880 152726 270908 163254
rect 271524 163146 271552 163254
rect 271602 163200 271658 164400
rect 271984 163254 272380 163282
rect 271616 163146 271644 163200
rect 271524 163118 271644 163146
rect 271880 159996 271932 160002
rect 271880 159938 271932 159944
rect 271420 154964 271472 154970
rect 271420 154906 271472 154912
rect 270868 152720 270920 152726
rect 270868 152662 270920 152668
rect 270604 151786 270816 151814
rect 270132 151778 270184 151784
rect 270144 150226 270172 151778
rect 270788 150226 270816 151786
rect 271432 150226 271460 154906
rect 264348 150198 264422 150226
rect 264992 150198 265066 150226
rect 265636 150198 265710 150226
rect 266280 150198 266354 150226
rect 266924 150198 266998 150226
rect 267568 150198 267642 150226
rect 268212 150198 268286 150226
rect 268856 150198 268930 150226
rect 269500 150198 269574 150226
rect 270144 150198 270218 150226
rect 270788 150198 270862 150226
rect 271432 150198 271506 150226
rect 271892 150210 271920 159938
rect 271984 153270 272012 163254
rect 272352 163146 272380 163254
rect 272430 163200 272486 164400
rect 273258 163200 273314 164400
rect 274086 163200 274142 164400
rect 274914 163200 274970 164400
rect 275112 163254 275784 163282
rect 272444 163146 272472 163200
rect 272352 163118 272472 163146
rect 273272 157214 273300 163200
rect 274100 159934 274128 163200
rect 274928 160002 274956 163200
rect 274916 159996 274968 160002
rect 274916 159938 274968 159944
rect 273352 159928 273404 159934
rect 273352 159870 273404 159876
rect 274088 159928 274140 159934
rect 274088 159870 274140 159876
rect 273260 157208 273312 157214
rect 273260 157150 273312 157156
rect 273260 156596 273312 156602
rect 273260 156538 273312 156544
rect 272064 154624 272116 154630
rect 272064 154566 272116 154572
rect 271972 153264 272024 153270
rect 271972 153206 272024 153212
rect 272076 150226 272104 154566
rect 273272 150226 273300 156538
rect 273364 151842 273392 159870
rect 273812 157480 273864 157486
rect 273812 157422 273864 157428
rect 273444 154896 273496 154902
rect 273444 154838 273496 154844
rect 273352 151836 273404 151842
rect 273456 151814 273484 154838
rect 273824 151814 273852 157422
rect 275112 154290 275140 163254
rect 275756 163146 275784 163254
rect 275834 163200 275890 164400
rect 276662 163200 276718 164400
rect 277490 163200 277546 164400
rect 278056 163254 278268 163282
rect 275848 163146 275876 163200
rect 275756 163118 275876 163146
rect 276112 160064 276164 160070
rect 276112 160006 276164 160012
rect 276020 156528 276072 156534
rect 276020 156470 276072 156476
rect 274640 154284 274692 154290
rect 274640 154226 274692 154232
rect 275100 154284 275152 154290
rect 275100 154226 275152 154232
rect 274546 153368 274602 153377
rect 274652 153338 274680 154226
rect 275926 153368 275982 153377
rect 274546 153303 274548 153312
rect 274600 153303 274602 153312
rect 274640 153332 274692 153338
rect 274548 153274 274600 153280
rect 274640 153274 274692 153280
rect 275836 153332 275888 153338
rect 275926 153303 275928 153312
rect 275836 153274 275888 153280
rect 275980 153303 275982 153312
rect 275928 153274 275980 153280
rect 275192 151904 275244 151910
rect 275192 151846 275244 151852
rect 273456 151786 273760 151814
rect 273824 151786 274588 151814
rect 273352 151778 273404 151784
rect 273732 150362 273760 151786
rect 273732 150334 273944 150362
rect 273916 150226 273944 150334
rect 274560 150226 274588 151786
rect 275204 150226 275232 151846
rect 275848 150226 275876 153274
rect 276032 151814 276060 156470
rect 276124 151910 276152 160006
rect 276676 157078 276704 163200
rect 277504 160070 277532 163200
rect 277492 160064 277544 160070
rect 277492 160006 277544 160012
rect 276664 157072 276716 157078
rect 276664 157014 276716 157020
rect 276480 154760 276532 154766
rect 276480 154702 276532 154708
rect 276112 151904 276164 151910
rect 276112 151846 276164 151852
rect 276492 151814 276520 154702
rect 278056 151978 278084 163254
rect 278240 163146 278268 163254
rect 278318 163200 278374 164400
rect 278792 163254 279096 163282
rect 278332 163146 278360 163200
rect 278240 163118 278360 163146
rect 278792 154358 278820 163254
rect 279068 163146 279096 163254
rect 279146 163200 279202 164400
rect 279974 163200 280030 164400
rect 280802 163200 280858 164400
rect 281630 163200 281686 164400
rect 281736 163254 282500 163282
rect 279160 163146 279188 163200
rect 279068 163118 279188 163146
rect 279792 159248 279844 159254
rect 279792 159190 279844 159196
rect 279056 156460 279108 156466
rect 279056 156402 279108 156408
rect 278412 154352 278464 154358
rect 278412 154294 278464 154300
rect 278780 154352 278832 154358
rect 278780 154294 278832 154300
rect 278044 151972 278096 151978
rect 278044 151914 278096 151920
rect 277768 151904 277820 151910
rect 277768 151846 277820 151852
rect 276032 151786 276428 151814
rect 276492 151786 277164 151814
rect 276400 150226 276428 151786
rect 277136 150226 277164 151786
rect 277780 150226 277808 151846
rect 278424 150226 278452 154294
rect 279068 150226 279096 156402
rect 279804 153134 279832 159190
rect 279988 157146 280016 163200
rect 280816 160070 280844 163200
rect 280160 160064 280212 160070
rect 280160 160006 280212 160012
rect 280804 160064 280856 160070
rect 280804 160006 280856 160012
rect 279976 157140 280028 157146
rect 279976 157082 280028 157088
rect 279332 153128 279384 153134
rect 279332 153070 279384 153076
rect 279792 153128 279844 153134
rect 279792 153070 279844 153076
rect 279344 151814 279372 153070
rect 280172 151910 280200 160006
rect 281644 159254 281672 163200
rect 281632 159248 281684 159254
rect 281632 159190 281684 159196
rect 281632 154828 281684 154834
rect 281632 154770 281684 154776
rect 280988 154488 281040 154494
rect 280988 154430 281040 154436
rect 280344 152924 280396 152930
rect 280344 152866 280396 152872
rect 280160 151904 280212 151910
rect 280160 151846 280212 151852
rect 279344 151786 279740 151814
rect 279712 150226 279740 151786
rect 280356 150226 280384 152866
rect 281000 150226 281028 154430
rect 281644 150226 281672 154770
rect 281736 154494 281764 163254
rect 282472 163146 282500 163254
rect 282550 163200 282606 164400
rect 283378 163200 283434 164400
rect 284206 163200 284262 164400
rect 284312 163254 284984 163282
rect 282564 163146 282592 163200
rect 282472 163118 282592 163146
rect 282828 159316 282880 159322
rect 282828 159258 282880 159264
rect 281724 154488 281776 154494
rect 281724 154430 281776 154436
rect 282276 153128 282328 153134
rect 282276 153070 282328 153076
rect 282288 150226 282316 153070
rect 282840 151814 282868 159258
rect 283392 157282 283420 163200
rect 284220 161474 284248 163200
rect 284128 161446 284248 161474
rect 283380 157276 283432 157282
rect 283380 157218 283432 157224
rect 283196 154556 283248 154562
rect 283196 154498 283248 154504
rect 283208 151814 283236 154498
rect 284128 152930 284156 161446
rect 284208 156664 284260 156670
rect 284208 156606 284260 156612
rect 284116 152924 284168 152930
rect 284116 152866 284168 152872
rect 282840 151786 282960 151814
rect 283208 151786 283604 151814
rect 282932 150226 282960 151786
rect 283576 150226 283604 151786
rect 284220 150226 284248 156606
rect 284312 153134 284340 163254
rect 284956 163146 284984 163254
rect 285034 163200 285090 164400
rect 285862 163200 285918 164400
rect 286690 163200 286746 164400
rect 287518 163200 287574 164400
rect 288346 163200 288402 164400
rect 289266 163200 289322 164400
rect 290094 163200 290150 164400
rect 290200 163254 290872 163282
rect 285048 163146 285076 163200
rect 284956 163118 285076 163146
rect 285876 154562 285904 163200
rect 286704 156670 286732 163200
rect 287532 159594 287560 163200
rect 287520 159588 287572 159594
rect 287520 159530 287572 159536
rect 287336 159520 287388 159526
rect 287336 159462 287388 159468
rect 288072 159520 288124 159526
rect 288072 159462 288124 159468
rect 287348 159322 287376 159462
rect 287336 159316 287388 159322
rect 287336 159258 287388 159264
rect 286784 156800 286836 156806
rect 286784 156742 286836 156748
rect 286692 156664 286744 156670
rect 286692 156606 286744 156612
rect 285864 154556 285916 154562
rect 285864 154498 285916 154504
rect 286140 153876 286192 153882
rect 286140 153818 286192 153824
rect 284300 153128 284352 153134
rect 284300 153070 284352 153076
rect 284852 152992 284904 152998
rect 284852 152934 284904 152940
rect 284864 150226 284892 152934
rect 285494 152416 285550 152425
rect 285494 152351 285550 152360
rect 285508 150226 285536 152351
rect 286152 150226 286180 153818
rect 286796 150226 286824 156742
rect 287428 152176 287480 152182
rect 287428 152118 287480 152124
rect 287440 150226 287468 152118
rect 288084 150226 288112 159462
rect 288360 159361 288388 163200
rect 288346 159352 288402 159361
rect 288346 159287 288402 159296
rect 289280 155718 289308 163200
rect 289360 156868 289412 156874
rect 289360 156810 289412 156816
rect 289268 155712 289320 155718
rect 289268 155654 289320 155660
rect 288714 153776 288770 153785
rect 288714 153711 288770 153720
rect 288728 150226 288756 153711
rect 289372 150226 289400 156810
rect 290108 156806 290136 163200
rect 290096 156800 290148 156806
rect 290096 156742 290148 156748
rect 290200 152998 290228 163254
rect 290844 163146 290872 163254
rect 290922 163200 290978 164400
rect 291750 163200 291806 164400
rect 292578 163200 292634 164400
rect 293406 163200 293462 164400
rect 294234 163200 294290 164400
rect 295154 163200 295210 164400
rect 295982 163200 296038 164400
rect 296810 163200 296866 164400
rect 297638 163200 297694 164400
rect 298466 163200 298522 164400
rect 299294 163200 299350 164400
rect 300122 163200 300178 164400
rect 300950 163200 301006 164400
rect 301870 163200 301926 164400
rect 302698 163200 302754 164400
rect 303526 163200 303582 164400
rect 303632 163254 304304 163282
rect 290936 163146 290964 163200
rect 290844 163118 290964 163146
rect 291660 159520 291712 159526
rect 291660 159462 291712 159468
rect 291672 159050 291700 159462
rect 291764 159050 291792 163200
rect 291660 159044 291712 159050
rect 291660 158986 291712 158992
rect 291752 159044 291804 159050
rect 291752 158986 291804 158992
rect 291936 156392 291988 156398
rect 291936 156334 291988 156340
rect 291292 153808 291344 153814
rect 291292 153750 291344 153756
rect 290188 152992 290240 152998
rect 290188 152934 290240 152940
rect 290004 152516 290056 152522
rect 290004 152458 290056 152464
rect 290016 150226 290044 152458
rect 290648 152312 290700 152318
rect 290648 152254 290700 152260
rect 290660 150226 290688 152254
rect 291304 150226 291332 153750
rect 291948 150226 291976 156334
rect 292592 155922 292620 163200
rect 293224 159316 293276 159322
rect 293224 159258 293276 159264
rect 292580 155916 292632 155922
rect 292580 155858 292632 155864
rect 292580 154692 292632 154698
rect 292580 154634 292632 154640
rect 292592 150226 292620 154634
rect 293236 150226 293264 159258
rect 293420 156738 293448 163200
rect 294248 159322 294276 163200
rect 295168 159526 295196 163200
rect 295064 159520 295116 159526
rect 295064 159462 295116 159468
rect 295156 159520 295208 159526
rect 295156 159462 295208 159468
rect 295076 159338 295104 159462
rect 294236 159316 294288 159322
rect 295076 159310 295380 159338
rect 294236 159258 294288 159264
rect 294512 159112 294564 159118
rect 294512 159054 294564 159060
rect 293960 159044 294012 159050
rect 293960 158986 294012 158992
rect 293408 156732 293460 156738
rect 293408 156674 293460 156680
rect 293868 153740 293920 153746
rect 293868 153682 293920 153688
rect 293880 150226 293908 153682
rect 293972 152318 294000 158986
rect 294052 156936 294104 156942
rect 294052 156878 294104 156884
rect 293960 152312 294012 152318
rect 293960 152254 294012 152260
rect 294064 151814 294092 156878
rect 294524 151814 294552 159054
rect 295352 152182 295380 159310
rect 295996 155786 296024 163200
rect 296824 156942 296852 163200
rect 297088 157004 297140 157010
rect 297088 156946 297140 156952
rect 296812 156936 296864 156942
rect 296812 156878 296864 156884
rect 295984 155780 296036 155786
rect 295984 155722 296036 155728
rect 296444 154012 296496 154018
rect 296444 153954 296496 153960
rect 295800 153060 295852 153066
rect 295800 153002 295852 153008
rect 295340 152176 295392 152182
rect 295340 152118 295392 152124
rect 294064 151786 294460 151814
rect 294524 151786 295196 151814
rect 294432 150226 294460 151786
rect 295168 150226 295196 151786
rect 295812 150226 295840 153002
rect 296456 150226 296484 153954
rect 297100 150226 297128 156946
rect 297652 152522 297680 163200
rect 298376 159180 298428 159186
rect 298376 159122 298428 159128
rect 297640 152516 297692 152522
rect 297640 152458 297692 152464
rect 297732 152176 297784 152182
rect 297732 152118 297784 152124
rect 297744 150226 297772 152118
rect 298388 150226 298416 159122
rect 298480 159050 298508 163200
rect 298468 159044 298520 159050
rect 298468 158986 298520 158992
rect 299308 155854 299336 163200
rect 299480 159044 299532 159050
rect 299480 158986 299532 158992
rect 299296 155848 299348 155854
rect 299296 155790 299348 155796
rect 299020 153944 299072 153950
rect 299020 153886 299072 153892
rect 299032 150226 299060 153886
rect 299492 152182 299520 158986
rect 299664 158024 299716 158030
rect 299664 157966 299716 157972
rect 299480 152176 299532 152182
rect 299480 152118 299532 152124
rect 299676 150226 299704 157966
rect 300136 156874 300164 163200
rect 300964 159118 300992 163200
rect 301884 159186 301912 163200
rect 301872 159180 301924 159186
rect 301872 159122 301924 159128
rect 300952 159112 301004 159118
rect 300952 159054 301004 159060
rect 300860 158976 300912 158982
rect 300860 158918 300912 158924
rect 300124 156868 300176 156874
rect 300124 156810 300176 156816
rect 300872 153202 300900 158918
rect 302332 158092 302384 158098
rect 302332 158034 302384 158040
rect 301596 153604 301648 153610
rect 301596 153546 301648 153552
rect 300308 153196 300360 153202
rect 300308 153138 300360 153144
rect 300860 153196 300912 153202
rect 300860 153138 300912 153144
rect 300320 150226 300348 153138
rect 300952 152788 301004 152794
rect 300952 152730 301004 152736
rect 300964 150226 300992 152730
rect 301608 150226 301636 153546
rect 302344 150226 302372 158034
rect 302712 155174 302740 163200
rect 303436 159384 303488 159390
rect 303436 159326 303488 159332
rect 302700 155168 302752 155174
rect 302700 155110 302752 155116
rect 302884 153196 302936 153202
rect 302884 153138 302936 153144
rect 263750 149940 263778 150198
rect 264394 149940 264422 150198
rect 265038 149940 265066 150198
rect 265682 149940 265710 150198
rect 266326 149940 266354 150198
rect 266970 149940 266998 150198
rect 267614 149940 267642 150198
rect 268258 149940 268286 150198
rect 268902 149940 268930 150198
rect 269546 149940 269574 150198
rect 270190 149940 270218 150198
rect 270834 149940 270862 150198
rect 271478 149940 271506 150198
rect 271880 150204 271932 150210
rect 272076 150198 272150 150226
rect 271880 150146 271932 150152
rect 272122 149940 272150 150198
rect 272754 150204 272806 150210
rect 273272 150198 273346 150226
rect 273916 150198 273990 150226
rect 274560 150198 274634 150226
rect 275204 150198 275278 150226
rect 275848 150198 275922 150226
rect 276400 150198 276566 150226
rect 277136 150198 277210 150226
rect 277780 150198 277854 150226
rect 278424 150198 278498 150226
rect 279068 150198 279142 150226
rect 279712 150198 279786 150226
rect 280356 150198 280430 150226
rect 281000 150198 281074 150226
rect 281644 150198 281718 150226
rect 282288 150198 282362 150226
rect 282932 150198 283006 150226
rect 283576 150198 283650 150226
rect 284220 150198 284294 150226
rect 284864 150198 284938 150226
rect 285508 150198 285582 150226
rect 286152 150198 286226 150226
rect 286796 150198 286870 150226
rect 287440 150198 287514 150226
rect 288084 150198 288158 150226
rect 288728 150198 288802 150226
rect 289372 150198 289446 150226
rect 290016 150198 290090 150226
rect 290660 150198 290734 150226
rect 291304 150198 291378 150226
rect 291948 150198 292022 150226
rect 292592 150198 292666 150226
rect 293236 150198 293310 150226
rect 293880 150198 293954 150226
rect 294432 150198 294598 150226
rect 295168 150198 295242 150226
rect 295812 150198 295886 150226
rect 296456 150198 296530 150226
rect 297100 150198 297174 150226
rect 297744 150198 297818 150226
rect 298388 150198 298462 150226
rect 299032 150198 299106 150226
rect 299676 150198 299750 150226
rect 300320 150198 300394 150226
rect 300964 150198 301038 150226
rect 301608 150198 301682 150226
rect 272754 150146 272806 150152
rect 272766 149940 272794 150146
rect 273318 149940 273346 150198
rect 273962 149940 273990 150198
rect 274606 149940 274634 150198
rect 275250 149940 275278 150198
rect 275894 149940 275922 150198
rect 276538 149940 276566 150198
rect 277182 149940 277210 150198
rect 277826 149940 277854 150198
rect 278470 149940 278498 150198
rect 279114 149940 279142 150198
rect 279758 149940 279786 150198
rect 280402 149940 280430 150198
rect 281046 149940 281074 150198
rect 281690 149940 281718 150198
rect 282334 149940 282362 150198
rect 282978 149940 283006 150198
rect 283622 149940 283650 150198
rect 284266 149940 284294 150198
rect 284910 149940 284938 150198
rect 285554 149940 285582 150198
rect 286198 149940 286226 150198
rect 286842 149940 286870 150198
rect 287486 149940 287514 150198
rect 288130 149940 288158 150198
rect 288774 149940 288802 150198
rect 289418 149940 289446 150198
rect 290062 149940 290090 150198
rect 290706 149940 290734 150198
rect 291350 149940 291378 150198
rect 291994 149940 292022 150198
rect 292638 149940 292666 150198
rect 293282 149940 293310 150198
rect 293926 149940 293954 150198
rect 294570 149940 294598 150198
rect 295214 149940 295242 150198
rect 295858 149940 295886 150198
rect 296502 149940 296530 150198
rect 297146 149940 297174 150198
rect 297790 149940 297818 150198
rect 298434 149940 298462 150198
rect 299078 149940 299106 150198
rect 299722 149940 299750 150198
rect 300366 149940 300394 150198
rect 301010 149940 301038 150198
rect 301654 149940 301682 150198
rect 302298 150198 302372 150226
rect 302896 150226 302924 153138
rect 303448 151814 303476 159326
rect 303540 152794 303568 163200
rect 303632 153202 303660 163254
rect 304276 163146 304304 163254
rect 304354 163200 304410 164400
rect 305182 163200 305238 164400
rect 306010 163200 306066 164400
rect 306838 163200 306894 164400
rect 307666 163200 307722 164400
rect 308586 163200 308642 164400
rect 309152 163254 309364 163282
rect 304368 163146 304396 163200
rect 304276 163118 304396 163146
rect 304724 155236 304776 155242
rect 304724 155178 304776 155184
rect 304080 153672 304132 153678
rect 304080 153614 304132 153620
rect 303620 153196 303672 153202
rect 303620 153138 303672 153144
rect 303528 152788 303580 152794
rect 303528 152730 303580 152736
rect 303448 151786 303568 151814
rect 303540 150226 303568 151786
rect 304092 150226 304120 153614
rect 304736 150226 304764 155178
rect 305196 153066 305224 163200
rect 306024 155242 306052 163200
rect 306852 159050 306880 163200
rect 307680 159390 307708 163200
rect 308496 159724 308548 159730
rect 308496 159666 308548 159672
rect 307760 159452 307812 159458
rect 307760 159394 307812 159400
rect 307668 159384 307720 159390
rect 307668 159326 307720 159332
rect 306840 159044 306892 159050
rect 306840 158986 306892 158992
rect 307300 158160 307352 158166
rect 307300 158102 307352 158108
rect 306012 155236 306064 155242
rect 306012 155178 306064 155184
rect 306656 154080 306708 154086
rect 306656 154022 306708 154028
rect 305184 153060 305236 153066
rect 305184 153002 305236 153008
rect 306012 152652 306064 152658
rect 306012 152594 306064 152600
rect 305368 152244 305420 152250
rect 305368 152186 305420 152192
rect 305380 150226 305408 152186
rect 306024 150226 306052 152594
rect 306668 150226 306696 154022
rect 307312 150226 307340 158102
rect 307772 151814 307800 159394
rect 308508 151814 308536 159666
rect 308600 159458 308628 163200
rect 308588 159452 308640 159458
rect 308588 159394 308640 159400
rect 309152 153882 309180 163254
rect 309336 163146 309364 163254
rect 309414 163200 309470 164400
rect 310242 163200 310298 164400
rect 310624 163254 311020 163282
rect 309428 163146 309456 163200
rect 309336 163118 309456 163146
rect 310256 158982 310284 163200
rect 310244 158976 310296 158982
rect 310244 158918 310296 158924
rect 309876 158228 309928 158234
rect 309876 158170 309928 158176
rect 309232 154148 309284 154154
rect 309232 154090 309284 154096
rect 309140 153876 309192 153882
rect 309140 153818 309192 153824
rect 307772 151786 307984 151814
rect 308508 151786 308628 151814
rect 307956 150226 307984 151786
rect 308600 150226 308628 151786
rect 309244 150226 309272 154090
rect 309888 150226 309916 158170
rect 310624 152658 310652 163254
rect 310992 163146 311020 163254
rect 311070 163200 311126 164400
rect 311898 163200 311954 164400
rect 312726 163200 312782 164400
rect 313554 163200 313610 164400
rect 314382 163200 314438 164400
rect 315302 163200 315358 164400
rect 316130 163200 316186 164400
rect 316958 163200 317014 164400
rect 317786 163200 317842 164400
rect 318614 163200 318670 164400
rect 318812 163254 319392 163282
rect 311084 163146 311112 163200
rect 310992 163118 311112 163146
rect 310704 158976 310756 158982
rect 310704 158918 310756 158924
rect 310612 152652 310664 152658
rect 310612 152594 310664 152600
rect 310520 152584 310572 152590
rect 310520 152526 310572 152532
rect 310532 150226 310560 152526
rect 310716 152425 310744 158918
rect 311808 153536 311860 153542
rect 311808 153478 311860 153484
rect 310702 152416 310758 152425
rect 310702 152351 310758 152360
rect 311164 152108 311216 152114
rect 311164 152050 311216 152056
rect 311176 150226 311204 152050
rect 311820 150226 311848 153478
rect 311912 152590 311940 163200
rect 311992 158908 312044 158914
rect 311992 158850 312044 158856
rect 311900 152584 311952 152590
rect 311900 152526 311952 152532
rect 302896 150198 302970 150226
rect 303540 150198 303614 150226
rect 304092 150198 304166 150226
rect 304736 150198 304810 150226
rect 305380 150198 305454 150226
rect 306024 150198 306098 150226
rect 306668 150198 306742 150226
rect 307312 150198 307386 150226
rect 307956 150198 308030 150226
rect 308600 150198 308674 150226
rect 309244 150198 309318 150226
rect 309888 150198 309962 150226
rect 310532 150198 310606 150226
rect 311176 150198 311250 150226
rect 311820 150198 311894 150226
rect 312004 150210 312032 158850
rect 312452 155304 312504 155310
rect 312452 155246 312504 155252
rect 312464 150226 312492 155246
rect 312740 155106 312768 163200
rect 313568 158982 313596 163200
rect 314396 159662 314424 163200
rect 315316 159730 315344 163200
rect 315304 159724 315356 159730
rect 315304 159666 315356 159672
rect 313740 159656 313792 159662
rect 313740 159598 313792 159604
rect 314384 159656 314436 159662
rect 314384 159598 314436 159604
rect 313556 158976 313608 158982
rect 313556 158918 313608 158924
rect 312728 155100 312780 155106
rect 312728 155042 312780 155048
rect 313752 150226 313780 159598
rect 315028 155372 315080 155378
rect 315028 155314 315080 155320
rect 314384 154216 314436 154222
rect 314384 154158 314436 154164
rect 314396 150226 314424 154158
rect 315040 150226 315068 155314
rect 316144 154086 316172 163200
rect 316972 161474 317000 163200
rect 316972 161446 317092 161474
rect 316960 154420 317012 154426
rect 316960 154362 317012 154368
rect 316132 154080 316184 154086
rect 316132 154022 316184 154028
rect 316316 152856 316368 152862
rect 316316 152798 316368 152804
rect 315672 152448 315724 152454
rect 315672 152390 315724 152396
rect 315684 150226 315712 152390
rect 316328 150226 316356 152798
rect 316972 150226 317000 154362
rect 317064 152454 317092 161446
rect 317144 159860 317196 159866
rect 317144 159802 317196 159808
rect 317156 152862 317184 159802
rect 317800 159798 317828 163200
rect 317788 159792 317840 159798
rect 317788 159734 317840 159740
rect 318628 158914 318656 163200
rect 318616 158908 318668 158914
rect 318616 158850 318668 158856
rect 318708 158840 318760 158846
rect 318708 158782 318760 158788
rect 317604 155440 317656 155446
rect 317604 155382 317656 155388
rect 317144 152856 317196 152862
rect 317144 152798 317196 152804
rect 317052 152448 317104 152454
rect 317052 152390 317104 152396
rect 317616 150226 317644 155382
rect 318248 152856 318300 152862
rect 318248 152798 318300 152804
rect 318260 150226 318288 152798
rect 318720 151814 318748 158782
rect 318812 153950 318840 163254
rect 319364 163146 319392 163254
rect 319442 163200 319498 164400
rect 320270 163200 320326 164400
rect 321098 163200 321154 164400
rect 322018 163200 322074 164400
rect 322846 163200 322902 164400
rect 322952 163254 323624 163282
rect 319456 163146 319484 163200
rect 319364 163118 319484 163146
rect 318892 159792 318944 159798
rect 318892 159734 318944 159740
rect 318800 153944 318852 153950
rect 318800 153886 318852 153892
rect 318904 152114 318932 159734
rect 319168 158908 319220 158914
rect 319168 158850 319220 158856
rect 319180 152250 319208 158850
rect 320284 158778 320312 163200
rect 321112 159866 321140 163200
rect 321100 159860 321152 159866
rect 321100 159802 321152 159808
rect 321560 159792 321612 159798
rect 321560 159734 321612 159740
rect 320272 158772 320324 158778
rect 320272 158714 320324 158720
rect 320180 155508 320232 155514
rect 320180 155450 320232 155456
rect 319536 153400 319588 153406
rect 319536 153342 319588 153348
rect 319168 152244 319220 152250
rect 319168 152186 319220 152192
rect 318892 152108 318944 152114
rect 318892 152050 318944 152056
rect 318720 151786 318932 151814
rect 318904 150226 318932 151786
rect 319548 150226 319576 153342
rect 320192 150226 320220 155450
rect 321572 152386 321600 159734
rect 322032 158778 322060 163200
rect 322020 158772 322072 158778
rect 322020 158714 322072 158720
rect 321836 155576 321888 155582
rect 321836 155518 321888 155524
rect 321744 153468 321796 153474
rect 321744 153410 321796 153416
rect 320824 152380 320876 152386
rect 320824 152322 320876 152328
rect 321560 152380 321612 152386
rect 321560 152322 321612 152328
rect 320836 150226 320864 152322
rect 321468 152040 321520 152046
rect 321468 151982 321520 151988
rect 321480 150226 321508 151982
rect 321756 150498 321784 153410
rect 321848 151814 321876 155518
rect 322860 154018 322888 163200
rect 322848 154012 322900 154018
rect 322848 153954 322900 153960
rect 322952 152862 322980 163254
rect 323596 163146 323624 163254
rect 323674 163200 323730 164400
rect 324502 163200 324558 164400
rect 324608 163254 325280 163282
rect 323688 163146 323716 163200
rect 323596 163118 323716 163146
rect 324516 160002 324544 163200
rect 324412 159996 324464 160002
rect 324412 159938 324464 159944
rect 324504 159996 324556 160002
rect 324504 159938 324556 159944
rect 324424 158914 324452 159938
rect 324044 158908 324096 158914
rect 324044 158850 324096 158856
rect 324412 158908 324464 158914
rect 324412 158850 324464 158856
rect 322940 152856 322992 152862
rect 322940 152798 322992 152804
rect 323400 152380 323452 152386
rect 323400 152322 323452 152328
rect 321848 151786 322796 151814
rect 321756 150470 322152 150498
rect 322124 150226 322152 150470
rect 322768 150226 322796 151786
rect 323412 150226 323440 152322
rect 324056 150226 324084 158850
rect 324608 152386 324636 163254
rect 325252 163146 325280 163254
rect 325330 163200 325386 164400
rect 325712 163254 326108 163282
rect 325344 163146 325372 163200
rect 325252 163118 325372 163146
rect 325332 155644 325384 155650
rect 325332 155586 325384 155592
rect 324688 153332 324740 153338
rect 324688 153274 324740 153280
rect 324596 152380 324648 152386
rect 324596 152322 324648 152328
rect 324700 150226 324728 153274
rect 325344 150226 325372 155586
rect 325712 154154 325740 163254
rect 326080 163146 326108 163254
rect 326158 163200 326214 164400
rect 326986 163200 327042 164400
rect 327906 163200 327962 164400
rect 328734 163200 328790 164400
rect 329562 163200 329618 164400
rect 329852 163254 330340 163282
rect 326172 163146 326200 163200
rect 326080 163118 326200 163146
rect 327000 159798 327028 163200
rect 326988 159792 327040 159798
rect 326988 159734 327040 159740
rect 327920 158778 327948 163200
rect 328368 159996 328420 160002
rect 328368 159938 328420 159944
rect 328460 159996 328512 160002
rect 328460 159938 328512 159944
rect 327908 158772 327960 158778
rect 327908 158714 327960 158720
rect 327632 157208 327684 157214
rect 327632 157150 327684 157156
rect 325700 154148 325752 154154
rect 325700 154090 325752 154096
rect 327264 153264 327316 153270
rect 327264 153206 327316 153212
rect 326620 152720 326672 152726
rect 326620 152662 326672 152668
rect 325976 151836 326028 151842
rect 325976 151778 326028 151784
rect 325988 150226 326016 151778
rect 326632 150226 326660 152662
rect 327276 150226 327304 153206
rect 327644 151814 327672 157150
rect 328380 151842 328408 159938
rect 328472 159254 328500 159938
rect 328748 159934 328776 163200
rect 328552 159928 328604 159934
rect 328552 159870 328604 159876
rect 328736 159928 328788 159934
rect 328736 159870 328788 159876
rect 328460 159248 328512 159254
rect 328460 159190 328512 159196
rect 328460 158908 328512 158914
rect 328460 158850 328512 158856
rect 328368 151836 328420 151842
rect 327644 151786 327948 151814
rect 327920 150226 327948 151786
rect 328368 151778 328420 151784
rect 302298 149940 302326 150198
rect 302942 149940 302970 150198
rect 303586 149940 303614 150198
rect 304138 149940 304166 150198
rect 304782 149940 304810 150198
rect 305426 149940 305454 150198
rect 306070 149940 306098 150198
rect 306714 149940 306742 150198
rect 307358 149940 307386 150198
rect 308002 149940 308030 150198
rect 308646 149940 308674 150198
rect 309290 149940 309318 150198
rect 309934 149940 309962 150198
rect 310578 149940 310606 150198
rect 311222 149940 311250 150198
rect 311866 149940 311894 150198
rect 311992 150204 312044 150210
rect 312464 150198 312538 150226
rect 311992 150146 312044 150152
rect 312510 149940 312538 150198
rect 313142 150204 313194 150210
rect 313752 150198 313826 150226
rect 314396 150198 314470 150226
rect 315040 150198 315114 150226
rect 315684 150198 315758 150226
rect 316328 150198 316402 150226
rect 316972 150198 317046 150226
rect 317616 150198 317690 150226
rect 318260 150198 318334 150226
rect 318904 150198 318978 150226
rect 319548 150198 319622 150226
rect 320192 150198 320266 150226
rect 320836 150198 320910 150226
rect 321480 150198 321554 150226
rect 322124 150198 322198 150226
rect 322768 150198 322842 150226
rect 323412 150198 323486 150226
rect 324056 150198 324130 150226
rect 324700 150198 324774 150226
rect 325344 150198 325418 150226
rect 325988 150198 326062 150226
rect 326632 150198 326706 150226
rect 327276 150198 327350 150226
rect 327920 150198 327994 150226
rect 328472 150210 328500 158850
rect 328564 150226 328592 159870
rect 328644 158908 328696 158914
rect 328644 158850 328696 158856
rect 328656 158710 328684 158850
rect 328644 158704 328696 158710
rect 328644 158646 328696 158652
rect 329576 155378 329604 163200
rect 329564 155372 329616 155378
rect 329564 155314 329616 155320
rect 329852 152726 329880 163254
rect 330312 163146 330340 163254
rect 330390 163200 330446 164400
rect 331218 163200 331274 164400
rect 331324 163254 331536 163282
rect 330404 163146 330432 163200
rect 330312 163118 330432 163146
rect 331232 163146 331260 163200
rect 331324 163146 331352 163254
rect 331232 163118 331352 163146
rect 331508 160070 331536 163254
rect 332046 163200 332102 164400
rect 332874 163200 332930 164400
rect 333702 163200 333758 164400
rect 334622 163200 334678 164400
rect 335450 163200 335506 164400
rect 335648 163254 336228 163282
rect 331496 160064 331548 160070
rect 331496 160006 331548 160012
rect 331312 159996 331364 160002
rect 331312 159938 331364 159944
rect 330484 157072 330536 157078
rect 330484 157014 330536 157020
rect 329932 154284 329984 154290
rect 329932 154226 329984 154232
rect 329840 152720 329892 152726
rect 329840 152662 329892 152668
rect 329944 150226 329972 154226
rect 313142 150146 313194 150152
rect 313154 149940 313182 150146
rect 313798 149940 313826 150198
rect 314442 149940 314470 150198
rect 315086 149940 315114 150198
rect 315730 149940 315758 150198
rect 316374 149940 316402 150198
rect 317018 149940 317046 150198
rect 317662 149940 317690 150198
rect 318306 149940 318334 150198
rect 318950 149940 318978 150198
rect 319594 149940 319622 150198
rect 320238 149940 320266 150198
rect 320882 149940 320910 150198
rect 321526 149940 321554 150198
rect 322170 149940 322198 150198
rect 322814 149940 322842 150198
rect 323458 149940 323486 150198
rect 324102 149940 324130 150198
rect 324746 149940 324774 150198
rect 325390 149940 325418 150198
rect 326034 149940 326062 150198
rect 326678 149940 326706 150198
rect 327322 149940 327350 150198
rect 327966 149940 327994 150198
rect 328460 150204 328512 150210
rect 328564 150198 328638 150226
rect 328460 150146 328512 150152
rect 328610 149940 328638 150198
rect 329242 150204 329294 150210
rect 329242 150146 329294 150152
rect 329898 150198 329972 150226
rect 330496 150226 330524 157014
rect 331324 152046 331352 159938
rect 332060 159254 332088 163200
rect 332600 159996 332652 160002
rect 332600 159938 332652 159944
rect 332048 159248 332100 159254
rect 332048 159190 332100 159196
rect 332416 154352 332468 154358
rect 332416 154294 332468 154300
rect 331312 152040 331364 152046
rect 331312 151982 331364 151988
rect 331772 151972 331824 151978
rect 331772 151914 331824 151920
rect 331128 151904 331180 151910
rect 331128 151846 331180 151852
rect 331140 150226 331168 151846
rect 331784 150226 331812 151914
rect 332428 150226 332456 154294
rect 330496 150198 330570 150226
rect 331140 150198 331214 150226
rect 331784 150198 331858 150226
rect 332428 150198 332502 150226
rect 332612 150210 332640 159938
rect 332888 155446 332916 163200
rect 333716 160002 333744 163200
rect 334636 160070 334664 163200
rect 334072 160064 334124 160070
rect 334072 160006 334124 160012
rect 334624 160064 334676 160070
rect 334624 160006 334676 160012
rect 333704 159996 333756 160002
rect 333704 159938 333756 159944
rect 333060 157140 333112 157146
rect 333060 157082 333112 157088
rect 332876 155440 332928 155446
rect 332876 155382 332928 155388
rect 333072 150226 333100 157082
rect 334084 151842 334112 160006
rect 335464 159254 335492 163200
rect 334532 159248 334584 159254
rect 334532 159190 334584 159196
rect 335452 159248 335504 159254
rect 335452 159190 335504 159196
rect 334348 152040 334400 152046
rect 334348 151982 334400 151988
rect 334072 151836 334124 151842
rect 334072 151778 334124 151784
rect 334360 150226 334388 151982
rect 334544 151910 334572 159190
rect 335544 157276 335596 157282
rect 335544 157218 335596 157224
rect 334900 154488 334952 154494
rect 334900 154430 334952 154436
rect 334532 151904 334584 151910
rect 334532 151846 334584 151852
rect 334912 150226 334940 154430
rect 335556 150226 335584 157218
rect 335648 154222 335676 163254
rect 336200 163146 336228 163254
rect 336278 163200 336334 164400
rect 337106 163200 337162 164400
rect 337934 163200 337990 164400
rect 338132 163254 338712 163282
rect 336292 163146 336320 163200
rect 336200 163118 336320 163146
rect 337016 159588 337068 159594
rect 337016 159530 337068 159536
rect 335636 154216 335688 154222
rect 335636 154158 335688 154164
rect 337028 153134 337056 159530
rect 337120 155514 337148 163200
rect 337948 159526 337976 163200
rect 337936 159520 337988 159526
rect 337936 159462 337988 159468
rect 337108 155508 337160 155514
rect 337108 155450 337160 155456
rect 337476 154556 337528 154562
rect 337476 154498 337528 154504
rect 336832 153128 336884 153134
rect 336832 153070 336884 153076
rect 337016 153128 337068 153134
rect 337016 153070 337068 153076
rect 336188 152924 336240 152930
rect 336188 152866 336240 152872
rect 336200 150226 336228 152866
rect 336844 150226 336872 153070
rect 337488 150226 337516 154498
rect 338132 152930 338160 163254
rect 338684 163146 338712 163254
rect 338762 163200 338818 164400
rect 339590 163200 339646 164400
rect 340418 163200 340474 164400
rect 340892 163254 341288 163282
rect 338776 163146 338804 163200
rect 338684 163118 338804 163146
rect 339500 159520 339552 159526
rect 339500 159462 339552 159468
rect 339406 159352 339462 159361
rect 339406 159287 339462 159296
rect 338212 156664 338264 156670
rect 338212 156606 338264 156612
rect 338120 152924 338172 152930
rect 338120 152866 338172 152872
rect 338224 150226 338252 156606
rect 338764 153128 338816 153134
rect 338764 153070 338816 153076
rect 329254 149940 329282 150146
rect 329898 149940 329926 150198
rect 330542 149940 330570 150198
rect 331186 149940 331214 150198
rect 331830 149940 331858 150198
rect 332474 149940 332502 150198
rect 332600 150204 332652 150210
rect 333072 150198 333146 150226
rect 332600 150146 332652 150152
rect 333118 149940 333146 150198
rect 333750 150204 333802 150210
rect 334360 150198 334434 150226
rect 334912 150198 334986 150226
rect 335556 150198 335630 150226
rect 336200 150198 336274 150226
rect 336844 150198 336918 150226
rect 337488 150198 337562 150226
rect 333750 150146 333802 150152
rect 333762 149940 333790 150146
rect 334406 149940 334434 150198
rect 334958 149940 334986 150198
rect 335602 149940 335630 150198
rect 336246 149940 336274 150198
rect 336890 149940 336918 150198
rect 337534 149940 337562 150198
rect 338178 150198 338252 150226
rect 338776 150226 338804 153070
rect 339420 150226 339448 159287
rect 339512 151910 339540 159462
rect 339604 154290 339632 163200
rect 339684 156800 339736 156806
rect 339684 156742 339736 156748
rect 339592 154284 339644 154290
rect 339592 154226 339644 154232
rect 339500 151904 339552 151910
rect 339500 151846 339552 151852
rect 338776 150198 338850 150226
rect 339420 150198 339494 150226
rect 339696 150210 339724 156742
rect 340052 155712 340104 155718
rect 340052 155654 340104 155660
rect 340064 150226 340092 155654
rect 340432 155582 340460 163200
rect 340420 155576 340472 155582
rect 340420 155518 340472 155524
rect 340892 153134 340920 163254
rect 341260 163146 341288 163254
rect 341338 163200 341394 164400
rect 342166 163200 342222 164400
rect 342272 163254 342944 163282
rect 341352 163146 341380 163200
rect 341260 163118 341380 163146
rect 342180 159594 342208 163200
rect 342168 159588 342220 159594
rect 342168 159530 342220 159536
rect 342272 154358 342300 163254
rect 342916 163146 342944 163254
rect 342994 163200 343050 164400
rect 343822 163200 343878 164400
rect 344650 163200 344706 164400
rect 345032 163254 345428 163282
rect 343008 163146 343036 163200
rect 342916 163118 343036 163146
rect 343836 159322 343864 163200
rect 344664 159526 344692 163200
rect 344560 159520 344612 159526
rect 344560 159462 344612 159468
rect 344652 159520 344704 159526
rect 344652 159462 344704 159468
rect 343640 159316 343692 159322
rect 343640 159258 343692 159264
rect 343824 159316 343876 159322
rect 343824 159258 343876 159264
rect 343272 156732 343324 156738
rect 343272 156674 343324 156680
rect 342352 155916 342404 155922
rect 342352 155858 342404 155864
rect 342260 154352 342312 154358
rect 342260 154294 342312 154300
rect 340880 153128 340932 153134
rect 340880 153070 340932 153076
rect 341340 152992 341392 152998
rect 341340 152934 341392 152940
rect 341352 150226 341380 152934
rect 341984 152312 342036 152318
rect 341984 152254 342036 152260
rect 341996 150226 342024 152254
rect 342364 151814 342392 155858
rect 342364 151786 342668 151814
rect 342640 150226 342668 151786
rect 343284 150226 343312 156674
rect 343652 151814 343680 159258
rect 343652 151786 343956 151814
rect 343928 150226 343956 151786
rect 344572 150226 344600 159462
rect 345032 152318 345060 163254
rect 345400 163146 345428 163254
rect 345478 163200 345534 164400
rect 345584 163254 346256 163282
rect 345492 163146 345520 163200
rect 345400 163118 345520 163146
rect 345204 155780 345256 155786
rect 345204 155722 345256 155728
rect 345020 152312 345072 152318
rect 345020 152254 345072 152260
rect 345216 150226 345244 155722
rect 345584 154426 345612 163254
rect 346228 163146 346256 163254
rect 346306 163200 346362 164400
rect 346412 163254 347084 163282
rect 346320 163146 346348 163200
rect 346228 163118 346348 163146
rect 345848 156936 345900 156942
rect 345848 156878 345900 156884
rect 345572 154420 345624 154426
rect 345572 154362 345624 154368
rect 345860 150226 345888 156878
rect 346412 152998 346440 163254
rect 347056 163146 347084 163254
rect 347134 163200 347190 164400
rect 347792 163254 348004 163282
rect 347148 163146 347176 163200
rect 347056 163118 347176 163146
rect 346400 152992 346452 152998
rect 346400 152934 346452 152940
rect 347792 152522 347820 163254
rect 347976 163146 348004 163254
rect 348054 163200 348110 164400
rect 348882 163200 348938 164400
rect 349264 163254 349660 163282
rect 348068 163146 348096 163200
rect 347976 163118 348096 163146
rect 348896 159390 348924 163200
rect 348792 159384 348844 159390
rect 348790 159352 348792 159361
rect 348884 159384 348936 159390
rect 348844 159352 348846 159361
rect 348884 159326 348936 159332
rect 348790 159287 348846 159296
rect 349068 159112 349120 159118
rect 349068 159054 349120 159060
rect 348056 156868 348108 156874
rect 348056 156810 348108 156816
rect 347872 155848 347924 155854
rect 347872 155790 347924 155796
rect 346492 152516 346544 152522
rect 346492 152458 346544 152464
rect 347780 152516 347832 152522
rect 347780 152458 347832 152464
rect 346504 150226 346532 152458
rect 347136 152176 347188 152182
rect 347136 152118 347188 152124
rect 347148 150226 347176 152118
rect 347884 150226 347912 155790
rect 348068 151814 348096 156810
rect 348068 151786 348464 151814
rect 338178 149940 338206 150198
rect 338822 149940 338850 150198
rect 339466 149940 339494 150198
rect 339684 150204 339736 150210
rect 340064 150198 340138 150226
rect 339684 150146 339736 150152
rect 340110 149940 340138 150198
rect 340742 150204 340794 150210
rect 341352 150198 341426 150226
rect 341996 150198 342070 150226
rect 342640 150198 342714 150226
rect 343284 150198 343358 150226
rect 343928 150198 344002 150226
rect 344572 150198 344646 150226
rect 345216 150198 345290 150226
rect 345860 150198 345934 150226
rect 346504 150198 346578 150226
rect 347148 150198 347222 150226
rect 340742 150146 340794 150152
rect 340754 149940 340782 150146
rect 341398 149940 341426 150198
rect 342042 149940 342070 150198
rect 342686 149940 342714 150198
rect 343330 149940 343358 150198
rect 343974 149940 344002 150198
rect 344618 149940 344646 150198
rect 345262 149940 345290 150198
rect 345906 149940 345934 150198
rect 346550 149940 346578 150198
rect 347194 149940 347222 150198
rect 347838 150198 347912 150226
rect 348436 150226 348464 151786
rect 349080 150226 349108 159054
rect 349264 154494 349292 163254
rect 349632 163146 349660 163254
rect 349710 163200 349766 164400
rect 350538 163200 350594 164400
rect 351366 163200 351422 164400
rect 351932 163254 352144 163282
rect 349724 163146 349752 163200
rect 349632 163118 349752 163146
rect 349804 159452 349856 159458
rect 349804 159394 349856 159400
rect 349896 159452 349948 159458
rect 349896 159394 349948 159400
rect 349712 159180 349764 159186
rect 349712 159122 349764 159128
rect 349344 155168 349396 155174
rect 349344 155110 349396 155116
rect 349252 154488 349304 154494
rect 349252 154430 349304 154436
rect 348436 150198 348510 150226
rect 349080 150198 349154 150226
rect 349356 150210 349384 155110
rect 349724 150226 349752 159122
rect 349816 158930 349844 159394
rect 349908 159361 349936 159394
rect 349894 159352 349950 159361
rect 349894 159287 349950 159296
rect 349988 159316 350040 159322
rect 349988 159258 350040 159264
rect 350000 159118 350028 159258
rect 349988 159112 350040 159118
rect 349988 159054 350040 159060
rect 350080 159044 350132 159050
rect 350080 158986 350132 158992
rect 350092 158930 350120 158986
rect 349816 158902 350120 158930
rect 350552 152182 350580 163200
rect 351380 159730 351408 163200
rect 351276 159724 351328 159730
rect 351276 159666 351328 159672
rect 351368 159724 351420 159730
rect 351368 159666 351420 159672
rect 351288 159390 351316 159666
rect 351276 159384 351328 159390
rect 351276 159326 351328 159332
rect 351644 153196 351696 153202
rect 351644 153138 351696 153144
rect 351000 152788 351052 152794
rect 351000 152730 351052 152736
rect 350540 152176 350592 152182
rect 350540 152118 350592 152124
rect 351012 150226 351040 152730
rect 351656 150226 351684 153138
rect 351932 152794 351960 163254
rect 352116 163146 352144 163254
rect 352194 163200 352250 164400
rect 352300 163254 352972 163282
rect 352208 163146 352236 163200
rect 352116 163118 352236 163146
rect 352300 154562 352328 163254
rect 352944 163146 352972 163254
rect 353022 163200 353078 164400
rect 353850 163200 353906 164400
rect 354770 163200 354826 164400
rect 355598 163200 355654 164400
rect 356072 163254 356376 163282
rect 353036 163146 353064 163200
rect 352944 163118 353064 163146
rect 353864 159186 353892 163200
rect 354220 159452 354272 159458
rect 354220 159394 354272 159400
rect 353300 159180 353352 159186
rect 353300 159122 353352 159128
rect 353852 159180 353904 159186
rect 353852 159122 353904 159128
rect 352932 155236 352984 155242
rect 352932 155178 352984 155184
rect 352288 154556 352340 154562
rect 352288 154498 352340 154504
rect 352288 153060 352340 153066
rect 352288 153002 352340 153008
rect 351920 152788 351972 152794
rect 351920 152730 351972 152736
rect 352300 150226 352328 153002
rect 352944 150226 352972 155178
rect 353312 151814 353340 159122
rect 353312 151786 353616 151814
rect 353588 150226 353616 151786
rect 354232 150226 354260 159394
rect 354784 153202 354812 163200
rect 355612 159390 355640 163200
rect 355600 159384 355652 159390
rect 355600 159326 355652 159332
rect 354864 159044 354916 159050
rect 354864 158986 354916 158992
rect 354772 153196 354824 153202
rect 354772 153138 354824 153144
rect 354876 150226 354904 158986
rect 356072 153882 356100 163254
rect 356348 163146 356376 163254
rect 356426 163200 356482 164400
rect 357254 163200 357310 164400
rect 358082 163200 358138 164400
rect 358910 163200 358966 164400
rect 359016 163254 359688 163282
rect 356440 163146 356468 163200
rect 356348 163118 356468 163146
rect 357268 158846 357296 163200
rect 357808 159724 357860 159730
rect 357808 159666 357860 159672
rect 357532 159656 357584 159662
rect 357532 159598 357584 159604
rect 357624 159656 357676 159662
rect 357624 159598 357676 159604
rect 357256 158840 357308 158846
rect 357256 158782 357308 158788
rect 355508 153876 355560 153882
rect 355508 153818 355560 153824
rect 356060 153876 356112 153882
rect 356060 153818 356112 153824
rect 355520 150226 355548 153818
rect 357544 152658 357572 159598
rect 357636 159458 357664 159598
rect 357624 159452 357676 159458
rect 357624 159394 357676 159400
rect 357820 159186 357848 159666
rect 358096 159458 358124 163200
rect 358820 159656 358872 159662
rect 358820 159598 358872 159604
rect 358084 159452 358136 159458
rect 358084 159394 358136 159400
rect 357716 159180 357768 159186
rect 357716 159122 357768 159128
rect 357808 159180 357860 159186
rect 357808 159122 357860 159128
rect 357728 159050 357756 159122
rect 357624 159044 357676 159050
rect 357624 158986 357676 158992
rect 357716 159044 357768 159050
rect 357716 158986 357768 158992
rect 356796 152652 356848 152658
rect 356796 152594 356848 152600
rect 357532 152652 357584 152658
rect 357532 152594 357584 152600
rect 356150 152416 356206 152425
rect 356150 152351 356206 152360
rect 356164 150226 356192 152351
rect 356808 150226 356836 152594
rect 357440 152584 357492 152590
rect 357440 152526 357492 152532
rect 357452 150226 357480 152526
rect 347838 149940 347866 150198
rect 348482 149940 348510 150198
rect 349126 149940 349154 150198
rect 349344 150204 349396 150210
rect 349724 150198 349798 150226
rect 349344 150146 349396 150152
rect 349770 149940 349798 150198
rect 350402 150204 350454 150210
rect 351012 150198 351086 150226
rect 351656 150198 351730 150226
rect 352300 150198 352374 150226
rect 352944 150198 353018 150226
rect 353588 150198 353662 150226
rect 354232 150198 354306 150226
rect 354876 150198 354950 150226
rect 355520 150198 355594 150226
rect 356164 150198 356238 150226
rect 356808 150198 356882 150226
rect 357452 150198 357526 150226
rect 357636 150210 357664 158986
rect 357900 155100 357952 155106
rect 357900 155042 357952 155048
rect 357912 151814 357940 155042
rect 358832 151814 358860 159598
rect 358924 153066 358952 163200
rect 359016 153814 359044 163254
rect 359660 163146 359688 163254
rect 359738 163200 359794 164400
rect 360212 163254 360608 163282
rect 359752 163146 359780 163200
rect 359660 163118 359780 163146
rect 359004 153808 359056 153814
rect 359004 153750 359056 153756
rect 358912 153060 358964 153066
rect 358912 153002 358964 153008
rect 359372 152652 359424 152658
rect 359372 152594 359424 152600
rect 357912 151786 358124 151814
rect 358832 151786 358952 151814
rect 358096 150226 358124 151786
rect 350402 150146 350454 150152
rect 350414 149940 350442 150146
rect 351058 149940 351086 150198
rect 351702 149940 351730 150198
rect 352346 149940 352374 150198
rect 352990 149940 353018 150198
rect 353634 149940 353662 150198
rect 354278 149940 354306 150198
rect 354922 149940 354950 150198
rect 355566 149940 355594 150198
rect 356210 149940 356238 150198
rect 356854 149940 356882 150198
rect 357498 149940 357526 150198
rect 357624 150204 357676 150210
rect 358096 150198 358170 150226
rect 358924 150210 358952 151786
rect 359384 150226 359412 152594
rect 359464 152584 359516 152590
rect 359464 152526 359516 152532
rect 359476 152046 359504 152526
rect 360212 152046 360240 163254
rect 360580 163146 360608 163254
rect 360658 163200 360714 164400
rect 360856 163254 361436 163282
rect 360672 163146 360700 163200
rect 360580 163118 360700 163146
rect 360660 154080 360712 154086
rect 360660 154022 360712 154028
rect 359464 152040 359516 152046
rect 359464 151982 359516 151988
rect 360200 152040 360252 152046
rect 360200 151982 360252 151988
rect 357624 150146 357676 150152
rect 358142 149940 358170 150198
rect 358774 150204 358826 150210
rect 358774 150146 358826 150152
rect 358912 150204 358964 150210
rect 359384 150198 359458 150226
rect 358912 150146 358964 150152
rect 358786 149940 358814 150146
rect 359430 149940 359458 150198
rect 360062 150204 360114 150210
rect 360062 150146 360114 150152
rect 360074 149940 360102 150146
rect 360672 150090 360700 154022
rect 360856 153270 360884 163254
rect 361408 163146 361436 163254
rect 361486 163200 361542 164400
rect 362314 163200 362370 164400
rect 363142 163200 363198 164400
rect 363970 163200 364026 164400
rect 364798 163200 364854 164400
rect 364904 163254 365576 163282
rect 361500 163146 361528 163200
rect 361408 163118 361528 163146
rect 362328 159662 362356 163200
rect 362316 159656 362368 159662
rect 362316 159598 362368 159604
rect 363052 158908 363104 158914
rect 363052 158850 363104 158856
rect 360844 153264 360896 153270
rect 360844 153206 360896 153212
rect 361764 152720 361816 152726
rect 361764 152662 361816 152668
rect 361776 152454 361804 152662
rect 361304 152448 361356 152454
rect 361304 152390 361356 152396
rect 361764 152448 361816 152454
rect 361764 152390 361816 152396
rect 361316 150090 361344 152390
rect 362592 152244 362644 152250
rect 362592 152186 362644 152192
rect 361948 152108 362000 152114
rect 361948 152050 362000 152056
rect 361960 150090 361988 152050
rect 362604 150090 362632 152186
rect 363064 150210 363092 158850
rect 363156 154086 363184 163200
rect 363236 159860 363288 159866
rect 363236 159802 363288 159808
rect 363144 154080 363196 154086
rect 363144 154022 363196 154028
rect 363144 153944 363196 153950
rect 363144 153886 363196 153892
rect 363156 150226 363184 153886
rect 363248 152658 363276 159802
rect 363984 158914 364012 163200
rect 364812 159866 364840 163200
rect 364800 159860 364852 159866
rect 364800 159802 364852 159808
rect 363972 158908 364024 158914
rect 363972 158850 364024 158856
rect 364904 157334 364932 163254
rect 365548 163146 365576 163254
rect 365626 163200 365682 164400
rect 365732 163254 366404 163282
rect 365640 163146 365668 163200
rect 365548 163118 365668 163146
rect 365168 158976 365220 158982
rect 365168 158918 365220 158924
rect 364812 157306 364932 157334
rect 363236 152652 363288 152658
rect 363236 152594 363288 152600
rect 364524 152652 364576 152658
rect 364524 152594 364576 152600
rect 363052 150204 363104 150210
rect 363156 150198 363322 150226
rect 363052 150146 363104 150152
rect 360672 150062 360746 150090
rect 361316 150062 361390 150090
rect 361960 150062 362034 150090
rect 362604 150062 362678 150090
rect 360718 149940 360746 150062
rect 361362 149940 361390 150062
rect 362006 149940 362034 150062
rect 362650 149940 362678 150062
rect 363294 149940 363322 150198
rect 363926 150204 363978 150210
rect 363926 150146 363978 150152
rect 363938 149940 363966 150146
rect 364536 150090 364564 152594
rect 364812 152114 364840 157306
rect 364984 153196 365036 153202
rect 364984 153138 365036 153144
rect 364996 153066 365024 153138
rect 364892 153060 364944 153066
rect 364892 153002 364944 153008
rect 364984 153060 365036 153066
rect 364984 153002 365036 153008
rect 364904 152946 364932 153002
rect 364904 152918 365116 152946
rect 365088 152658 365116 152918
rect 365076 152652 365128 152658
rect 365076 152594 365128 152600
rect 364800 152108 364852 152114
rect 364800 152050 364852 152056
rect 365180 150226 365208 158918
rect 365732 153746 365760 163254
rect 366376 163146 366404 163254
rect 366454 163200 366510 164400
rect 367374 163200 367430 164400
rect 367572 163254 368152 163282
rect 366468 163146 366496 163200
rect 366376 163118 366496 163146
rect 367388 158778 367416 163200
rect 367376 158772 367428 158778
rect 367376 158714 367428 158720
rect 365812 154012 365864 154018
rect 365812 153954 365864 153960
rect 365720 153740 365772 153746
rect 365720 153682 365772 153688
rect 365180 150198 365254 150226
rect 364536 150062 364610 150090
rect 364582 149940 364610 150062
rect 365226 149940 365254 150198
rect 365824 150090 365852 153954
rect 367572 152862 367600 163254
rect 368124 163146 368152 163254
rect 368202 163200 368258 164400
rect 369030 163200 369086 164400
rect 369858 163200 369914 164400
rect 370686 163200 370742 164400
rect 371514 163200 371570 164400
rect 371804 163254 372292 163282
rect 368216 163146 368244 163200
rect 368124 163118 368244 163146
rect 368940 159792 368992 159798
rect 368940 159734 368992 159740
rect 368480 158704 368532 158710
rect 368480 158646 368532 158652
rect 368296 154148 368348 154154
rect 368296 154090 368348 154096
rect 366364 152856 366416 152862
rect 366364 152798 366416 152804
rect 367560 152856 367612 152862
rect 367560 152798 367612 152804
rect 365778 150062 365852 150090
rect 366376 150090 366404 152798
rect 367008 152720 367060 152726
rect 367008 152662 367060 152668
rect 367020 150090 367048 152662
rect 367100 152584 367152 152590
rect 367100 152526 367152 152532
rect 367112 152046 367140 152526
rect 367652 152380 367704 152386
rect 367652 152322 367704 152328
rect 367744 152380 367796 152386
rect 367744 152322 367796 152328
rect 367100 152040 367152 152046
rect 367100 151982 367152 151988
rect 367664 150090 367692 152322
rect 367756 152114 367784 152322
rect 367744 152108 367796 152114
rect 367744 152050 367796 152056
rect 368308 150090 368336 154090
rect 368492 150210 368520 158646
rect 368952 150226 368980 159734
rect 369044 159730 369072 163200
rect 369032 159724 369084 159730
rect 369032 159666 369084 159672
rect 369872 155242 369900 163200
rect 370044 159928 370096 159934
rect 370044 159870 370096 159876
rect 369860 155236 369912 155242
rect 369860 155178 369912 155184
rect 370056 151814 370084 159870
rect 370700 152250 370728 163200
rect 371528 158982 371556 163200
rect 371516 158976 371568 158982
rect 371516 158918 371568 158924
rect 370872 155372 370924 155378
rect 370872 155314 370924 155320
rect 370688 152244 370740 152250
rect 370688 152186 370740 152192
rect 370056 151786 370268 151814
rect 370240 150226 370268 151786
rect 370884 150226 370912 155314
rect 371516 152448 371568 152454
rect 371516 152390 371568 152396
rect 371528 150226 371556 152390
rect 371804 152386 371832 163254
rect 372264 163146 372292 163254
rect 372342 163200 372398 164400
rect 373170 163200 373226 164400
rect 374090 163200 374146 164400
rect 374918 163200 374974 164400
rect 375746 163200 375802 164400
rect 376574 163200 376630 164400
rect 376772 163254 377352 163282
rect 372356 163146 372384 163200
rect 372264 163118 372384 163146
rect 373184 155310 373212 163200
rect 374000 159996 374052 160002
rect 374000 159938 374052 159944
rect 373448 155440 373500 155446
rect 373448 155382 373500 155388
rect 373172 155304 373224 155310
rect 373172 155246 373224 155252
rect 371792 152380 371844 152386
rect 371792 152322 371844 152328
rect 372804 151972 372856 151978
rect 372804 151914 372856 151920
rect 372160 151836 372212 151842
rect 372160 151778 372212 151784
rect 372172 150226 372200 151778
rect 372816 150226 372844 151914
rect 373460 150226 373488 155382
rect 374012 151814 374040 159938
rect 374104 159934 374132 163200
rect 374736 160064 374788 160070
rect 374736 160006 374788 160012
rect 374092 159928 374144 159934
rect 374092 159870 374144 159876
rect 374012 151786 374132 151814
rect 374104 150226 374132 151786
rect 374748 150226 374776 160006
rect 374932 160002 374960 163200
rect 374920 159996 374972 160002
rect 374920 159938 374972 159944
rect 375760 159798 375788 163200
rect 375748 159792 375800 159798
rect 375748 159734 375800 159740
rect 375380 159248 375432 159254
rect 375380 159190 375432 159196
rect 375392 150226 375420 159190
rect 376588 155378 376616 163200
rect 376668 155508 376720 155514
rect 376668 155450 376720 155456
rect 376576 155372 376628 155378
rect 376576 155314 376628 155320
rect 376024 154216 376076 154222
rect 376024 154158 376076 154164
rect 376036 150226 376064 154158
rect 376680 150226 376708 155450
rect 376772 151978 376800 163254
rect 377324 163146 377352 163254
rect 377402 163200 377458 164400
rect 378230 163200 378286 164400
rect 379058 163200 379114 164400
rect 379624 163254 379836 163282
rect 377416 163146 377444 163200
rect 377324 163118 377444 163146
rect 377772 159112 377824 159118
rect 377772 159054 377824 159060
rect 377784 152114 377812 159054
rect 377956 152924 378008 152930
rect 377956 152866 378008 152872
rect 377772 152108 377824 152114
rect 377772 152050 377824 152056
rect 376760 151972 376812 151978
rect 376760 151914 376812 151920
rect 377312 151904 377364 151910
rect 377312 151846 377364 151852
rect 377324 150226 377352 151846
rect 377968 150226 377996 152866
rect 378244 151910 378272 163200
rect 378600 154284 378652 154290
rect 378600 154226 378652 154232
rect 378232 151904 378284 151910
rect 378232 151846 378284 151852
rect 378612 150226 378640 154226
rect 379072 152726 379100 163200
rect 379244 155576 379296 155582
rect 379244 155518 379296 155524
rect 379060 152720 379112 152726
rect 379060 152662 379112 152668
rect 379256 150226 379284 155518
rect 379624 154018 379652 163254
rect 379808 163146 379836 163254
rect 379886 163200 379942 164400
rect 380806 163200 380862 164400
rect 381634 163200 381690 164400
rect 382462 163200 382518 164400
rect 383290 163200 383346 164400
rect 383764 163254 384068 163282
rect 379900 163146 379928 163200
rect 379808 163118 379928 163146
rect 380820 159934 380848 163200
rect 381648 160070 381676 163200
rect 381636 160064 381688 160070
rect 381636 160006 381688 160012
rect 380716 159928 380768 159934
rect 380716 159870 380768 159876
rect 380808 159928 380860 159934
rect 380808 159870 380860 159876
rect 380728 159594 380756 159870
rect 380532 159588 380584 159594
rect 380532 159530 380584 159536
rect 380716 159588 380768 159594
rect 380716 159530 380768 159536
rect 379612 154012 379664 154018
rect 379612 153954 379664 153960
rect 379888 153128 379940 153134
rect 379888 153070 379940 153076
rect 379900 150226 379928 153070
rect 380544 150226 380572 159530
rect 380900 159112 380952 159118
rect 380900 159054 380952 159060
rect 380912 152930 380940 159054
rect 382476 159050 382504 163200
rect 382556 159520 382608 159526
rect 382556 159462 382608 159468
rect 382464 159044 382516 159050
rect 382464 158986 382516 158992
rect 380992 158840 381044 158846
rect 380992 158782 381044 158788
rect 380900 152924 380952 152930
rect 380900 152866 380952 152872
rect 381004 151842 381032 158782
rect 381176 154352 381228 154358
rect 381176 154294 381228 154300
rect 380992 151836 381044 151842
rect 380992 151778 381044 151784
rect 381188 150226 381216 154294
rect 381820 152108 381872 152114
rect 381820 152050 381872 152056
rect 381832 150226 381860 152050
rect 382568 150226 382596 159462
rect 383304 153950 383332 163200
rect 383292 153944 383344 153950
rect 383292 153886 383344 153892
rect 383764 152998 383792 163254
rect 384040 163146 384068 163254
rect 384118 163200 384174 164400
rect 384946 163200 385002 164400
rect 385774 163200 385830 164400
rect 386602 163200 386658 164400
rect 387522 163200 387578 164400
rect 388350 163200 388406 164400
rect 389178 163200 389234 164400
rect 389744 163254 389956 163282
rect 384132 163146 384160 163200
rect 384040 163118 384160 163146
rect 383844 154420 383896 154426
rect 383844 154362 383896 154368
rect 383752 152992 383804 152998
rect 383752 152934 383804 152940
rect 383200 152924 383252 152930
rect 383200 152866 383252 152872
rect 383212 152318 383240 152866
rect 383108 152312 383160 152318
rect 383108 152254 383160 152260
rect 383200 152312 383252 152318
rect 383200 152254 383252 152260
rect 368480 150204 368532 150210
rect 368952 150198 369026 150226
rect 368480 150146 368532 150152
rect 366376 150062 366450 150090
rect 367020 150062 367094 150090
rect 367664 150062 367738 150090
rect 368308 150062 368382 150090
rect 365778 149940 365806 150062
rect 366422 149940 366450 150062
rect 367066 149940 367094 150062
rect 367710 149940 367738 150062
rect 368354 149940 368382 150062
rect 368998 149940 369026 150198
rect 369630 150204 369682 150210
rect 370240 150198 370314 150226
rect 370884 150198 370958 150226
rect 371528 150198 371602 150226
rect 372172 150198 372246 150226
rect 372816 150198 372890 150226
rect 373460 150198 373534 150226
rect 374104 150198 374178 150226
rect 374748 150198 374822 150226
rect 375392 150198 375466 150226
rect 376036 150198 376110 150226
rect 376680 150198 376754 150226
rect 377324 150198 377398 150226
rect 377968 150198 378042 150226
rect 378612 150198 378686 150226
rect 379256 150198 379330 150226
rect 379900 150198 379974 150226
rect 380544 150198 380618 150226
rect 381188 150198 381262 150226
rect 381832 150198 381906 150226
rect 369630 150146 369682 150152
rect 369642 149940 369670 150146
rect 370286 149940 370314 150198
rect 370930 149940 370958 150198
rect 371574 149940 371602 150198
rect 372218 149940 372246 150198
rect 372862 149940 372890 150198
rect 373506 149940 373534 150198
rect 374150 149940 374178 150198
rect 374794 149940 374822 150198
rect 375438 149940 375466 150198
rect 376082 149940 376110 150198
rect 376726 149940 376754 150198
rect 377370 149940 377398 150198
rect 378014 149940 378042 150198
rect 378658 149940 378686 150198
rect 379302 149940 379330 150198
rect 379946 149940 379974 150198
rect 380590 149940 380618 150198
rect 381234 149940 381262 150198
rect 381878 149940 381906 150198
rect 382522 150198 382596 150226
rect 383120 150226 383148 152254
rect 383856 150226 383884 154362
rect 384960 153134 384988 163200
rect 385788 159594 385816 163200
rect 385776 159588 385828 159594
rect 385776 159530 385828 159536
rect 385592 159316 385644 159322
rect 385592 159258 385644 159264
rect 384948 153128 385000 153134
rect 384948 153070 385000 153076
rect 384396 152924 384448 152930
rect 384396 152866 384448 152872
rect 383120 150198 383194 150226
rect 382522 149940 382550 150198
rect 383166 149940 383194 150198
rect 383810 150198 383884 150226
rect 384408 150226 384436 152866
rect 385040 152516 385092 152522
rect 385040 152458 385092 152464
rect 385052 150226 385080 152458
rect 385604 151814 385632 159258
rect 385868 158908 385920 158914
rect 385868 158850 385920 158856
rect 385880 151910 385908 158850
rect 386052 158772 386104 158778
rect 386052 158714 386104 158720
rect 386064 151978 386092 158714
rect 386328 154488 386380 154494
rect 386328 154430 386380 154436
rect 386052 151972 386104 151978
rect 386052 151914 386104 151920
rect 385868 151904 385920 151910
rect 385868 151846 385920 151852
rect 385604 151786 385724 151814
rect 385696 150226 385724 151786
rect 386340 150226 386368 154430
rect 386616 154222 386644 163200
rect 387536 158778 387564 163200
rect 388364 159322 388392 163200
rect 389192 159934 389220 163200
rect 388628 159928 388680 159934
rect 388628 159870 388680 159876
rect 389180 159928 389232 159934
rect 389180 159870 389232 159876
rect 388352 159316 388404 159322
rect 388352 159258 388404 159264
rect 387616 159180 387668 159186
rect 387616 159122 387668 159128
rect 387524 158772 387576 158778
rect 387524 158714 387576 158720
rect 386604 154216 386656 154222
rect 386604 154158 386656 154164
rect 386972 152176 387024 152182
rect 386972 152118 387024 152124
rect 386984 150226 387012 152118
rect 387628 150226 387656 159122
rect 388444 152924 388496 152930
rect 388444 152866 388496 152872
rect 388260 152788 388312 152794
rect 388260 152730 388312 152736
rect 388272 150226 388300 152730
rect 388456 152726 388484 152866
rect 388444 152720 388496 152726
rect 388444 152662 388496 152668
rect 388536 152720 388588 152726
rect 388536 152662 388588 152668
rect 388548 152182 388576 152662
rect 388640 152182 388668 159870
rect 388720 159520 388772 159526
rect 388720 159462 388772 159468
rect 388536 152176 388588 152182
rect 388536 152118 388588 152124
rect 388628 152176 388680 152182
rect 388628 152118 388680 152124
rect 388732 152046 388760 159462
rect 388904 154556 388956 154562
rect 388904 154498 388956 154504
rect 388720 152040 388772 152046
rect 388720 151982 388772 151988
rect 388916 150226 388944 154498
rect 389744 154154 389772 163254
rect 389928 163146 389956 163254
rect 390006 163200 390062 164400
rect 390834 163200 390890 164400
rect 391662 163200 391718 164400
rect 392490 163200 392546 164400
rect 393410 163200 393466 164400
rect 394238 163200 394294 164400
rect 395066 163200 395122 164400
rect 395894 163200 395950 164400
rect 396092 163254 396672 163282
rect 390020 163146 390048 163200
rect 389928 163118 390048 163146
rect 390744 159384 390796 159390
rect 390744 159326 390796 159332
rect 390560 158772 390612 158778
rect 390560 158714 390612 158720
rect 389732 154148 389784 154154
rect 389732 154090 389784 154096
rect 390192 153060 390244 153066
rect 390192 153002 390244 153008
rect 389548 152312 389600 152318
rect 389548 152254 389600 152260
rect 389560 150226 389588 152254
rect 390204 150226 390232 153002
rect 390572 152318 390600 158714
rect 390560 152312 390612 152318
rect 390560 152254 390612 152260
rect 390756 151814 390784 159326
rect 390848 159118 390876 163200
rect 391676 159254 391704 163200
rect 392400 159452 392452 159458
rect 392400 159394 392452 159400
rect 391664 159248 391716 159254
rect 391664 159190 391716 159196
rect 390836 159112 390888 159118
rect 390836 159054 390888 159060
rect 391940 159112 391992 159118
rect 391940 159054 391992 159060
rect 391480 153876 391532 153882
rect 391480 153818 391532 153824
rect 390756 151786 390876 151814
rect 390848 150226 390876 151786
rect 391492 150226 391520 153818
rect 391952 153066 391980 159054
rect 391940 153060 391992 153066
rect 391940 153002 391992 153008
rect 392124 151836 392176 151842
rect 392412 151814 392440 159394
rect 392504 159186 392532 163200
rect 392492 159180 392544 159186
rect 392492 159122 392544 159128
rect 393424 154290 393452 163200
rect 393412 154284 393464 154290
rect 393412 154226 393464 154232
rect 394056 153808 394108 153814
rect 394056 153750 394108 153756
rect 393412 152652 393464 152658
rect 393412 152594 393464 152600
rect 392412 151786 392808 151814
rect 392124 151778 392176 151784
rect 392136 150226 392164 151778
rect 392780 150226 392808 151786
rect 393424 150226 393452 152594
rect 394068 150226 394096 153750
rect 394252 152522 394280 163200
rect 395080 159458 395108 163200
rect 395528 159860 395580 159866
rect 395528 159802 395580 159808
rect 395252 159656 395304 159662
rect 395252 159598 395304 159604
rect 395068 159452 395120 159458
rect 395068 159394 395120 159400
rect 395160 153196 395212 153202
rect 395160 153138 395212 153144
rect 394700 152584 394752 152590
rect 394700 152526 394752 152532
rect 394240 152516 394292 152522
rect 394240 152458 394292 152464
rect 394712 150226 394740 152526
rect 384408 150198 384482 150226
rect 385052 150198 385126 150226
rect 385696 150198 385770 150226
rect 386340 150198 386414 150226
rect 386984 150198 387058 150226
rect 387628 150198 387702 150226
rect 388272 150198 388346 150226
rect 388916 150198 388990 150226
rect 389560 150198 389634 150226
rect 390204 150198 390278 150226
rect 390848 150198 390922 150226
rect 391492 150198 391566 150226
rect 392136 150198 392210 150226
rect 392780 150198 392854 150226
rect 393424 150198 393498 150226
rect 394068 150198 394142 150226
rect 394712 150198 394786 150226
rect 383810 149940 383838 150198
rect 384454 149940 384482 150198
rect 385098 149940 385126 150198
rect 385742 149940 385770 150198
rect 386386 149940 386414 150198
rect 387030 149940 387058 150198
rect 387674 149940 387702 150198
rect 388318 149940 388346 150198
rect 388962 149940 388990 150198
rect 389606 149940 389634 150198
rect 390250 149940 390278 150198
rect 390894 149940 390922 150198
rect 391538 149940 391566 150198
rect 392182 149940 392210 150198
rect 392826 149940 392854 150198
rect 393470 149940 393498 150198
rect 394114 149940 394142 150198
rect 394758 149940 394786 150198
rect 395172 150192 395200 153138
rect 395264 151814 395292 159598
rect 395540 153202 395568 159802
rect 395528 153196 395580 153202
rect 395528 153138 395580 153144
rect 395908 152862 395936 163200
rect 396092 153882 396120 163254
rect 396644 163146 396672 163254
rect 396722 163200 396778 164400
rect 397550 163200 397606 164400
rect 398378 163200 398434 164400
rect 399206 163200 399262 164400
rect 400126 163200 400182 164400
rect 400324 163254 400904 163282
rect 396736 163146 396764 163200
rect 396644 163118 396764 163146
rect 397368 158976 397420 158982
rect 397368 158918 397420 158924
rect 396540 154080 396592 154086
rect 396540 154022 396592 154028
rect 396080 153876 396132 153882
rect 396080 153818 396132 153824
rect 395896 152856 395948 152862
rect 395896 152798 395948 152804
rect 395264 151786 396028 151814
rect 396000 150226 396028 151786
rect 396552 150226 396580 154022
rect 397184 151904 397236 151910
rect 397184 151846 397236 151852
rect 397196 150226 397224 151846
rect 397380 151842 397408 158918
rect 397564 152590 397592 163200
rect 397920 159996 397972 160002
rect 397920 159938 397972 159944
rect 397828 153196 397880 153202
rect 397828 153138 397880 153144
rect 397552 152584 397604 152590
rect 397552 152526 397604 152532
rect 397368 151836 397420 151842
rect 397368 151778 397420 151784
rect 397840 150226 397868 153138
rect 397932 151910 397960 159938
rect 398392 158846 398420 163200
rect 398840 160064 398892 160070
rect 398840 160006 398892 160012
rect 398380 158840 398432 158846
rect 398380 158782 398432 158788
rect 398852 152454 398880 160006
rect 399220 160002 399248 163200
rect 399208 159996 399260 160002
rect 399208 159938 399260 159944
rect 400140 154086 400168 163200
rect 400324 154358 400352 163254
rect 400876 163146 400904 163254
rect 400954 163200 401010 164400
rect 401782 163200 401838 164400
rect 401888 163254 402560 163282
rect 400968 163146 400996 163200
rect 400876 163118 400996 163146
rect 401796 160070 401824 163200
rect 401784 160064 401836 160070
rect 401784 160006 401836 160012
rect 401048 159724 401100 159730
rect 401048 159666 401100 159672
rect 400312 154352 400364 154358
rect 400312 154294 400364 154300
rect 400128 154080 400180 154086
rect 400128 154022 400180 154028
rect 399116 153740 399168 153746
rect 399116 153682 399168 153688
rect 398472 152448 398524 152454
rect 398472 152390 398524 152396
rect 398840 152448 398892 152454
rect 398840 152390 398892 152396
rect 397920 151904 397972 151910
rect 397920 151846 397972 151852
rect 398484 150226 398512 152390
rect 399128 150226 399156 153682
rect 400404 152788 400456 152794
rect 400404 152730 400456 152736
rect 399760 151972 399812 151978
rect 399760 151914 399812 151920
rect 399772 150226 399800 151914
rect 400416 150226 400444 152730
rect 401060 150226 401088 159666
rect 401600 159316 401652 159322
rect 401600 159258 401652 159264
rect 401612 153202 401640 159258
rect 401692 155236 401744 155242
rect 401692 155178 401744 155184
rect 401600 153196 401652 153202
rect 401600 153138 401652 153144
rect 401704 150226 401732 155178
rect 401888 152658 401916 163254
rect 402532 163146 402560 163254
rect 402610 163200 402666 164400
rect 403438 163200 403494 164400
rect 404266 163200 404322 164400
rect 405094 163200 405150 164400
rect 405922 163200 405978 164400
rect 406842 163200 406898 164400
rect 407670 163200 407726 164400
rect 408498 163200 408554 164400
rect 409064 163254 409276 163282
rect 402624 163146 402652 163200
rect 402532 163118 402652 163146
rect 403452 159730 403480 163200
rect 403440 159724 403492 159730
rect 403440 159666 403492 159672
rect 404280 159390 404308 163200
rect 404268 159384 404320 159390
rect 404268 159326 404320 159332
rect 403900 159248 403952 159254
rect 403900 159190 403952 159196
rect 403164 155304 403216 155310
rect 403164 155246 403216 155252
rect 401876 152652 401928 152658
rect 401876 152594 401928 152600
rect 402336 152244 402388 152250
rect 402336 152186 402388 152192
rect 402348 150226 402376 152186
rect 402980 151836 403032 151842
rect 402980 151778 403032 151784
rect 402992 150226 403020 151778
rect 396000 150198 396074 150226
rect 396552 150198 396626 150226
rect 397196 150198 397270 150226
rect 397840 150198 397914 150226
rect 398484 150198 398558 150226
rect 399128 150198 399202 150226
rect 399772 150198 399846 150226
rect 400416 150198 400490 150226
rect 401060 150198 401134 150226
rect 401704 150198 401778 150226
rect 402348 150198 402422 150226
rect 402992 150198 403066 150226
rect 403176 150210 403204 155246
rect 403912 152386 403940 159190
rect 404636 158840 404688 158846
rect 404636 158782 404688 158788
rect 403624 152380 403676 152386
rect 403624 152322 403676 152328
rect 403900 152380 403952 152386
rect 403900 152322 403952 152328
rect 403636 150226 403664 152322
rect 404648 151978 404676 158782
rect 405108 158778 405136 163200
rect 405832 159792 405884 159798
rect 405832 159734 405884 159740
rect 405648 159452 405700 159458
rect 405648 159394 405700 159400
rect 405096 158772 405148 158778
rect 405096 158714 405148 158720
rect 404912 152040 404964 152046
rect 404912 151982 404964 151988
rect 404636 151972 404688 151978
rect 404636 151914 404688 151920
rect 404924 150226 404952 151982
rect 405660 151910 405688 159394
rect 405556 151904 405608 151910
rect 405556 151846 405608 151852
rect 405648 151904 405700 151910
rect 405648 151846 405700 151852
rect 405568 150226 405596 151846
rect 405844 151814 405872 159734
rect 405936 152862 405964 163200
rect 406856 159798 406884 163200
rect 407580 160064 407632 160070
rect 407580 160006 407632 160012
rect 406844 159792 406896 159798
rect 406844 159734 406896 159740
rect 406844 155372 406896 155378
rect 406844 155314 406896 155320
rect 405924 152856 405976 152862
rect 405924 152798 405976 152804
rect 405844 151786 406240 151814
rect 406212 150226 406240 151786
rect 406856 150226 406884 155314
rect 407488 152720 407540 152726
rect 407488 152662 407540 152668
rect 407500 150226 407528 152662
rect 407592 152046 407620 160006
rect 407684 159662 407712 163200
rect 407672 159656 407724 159662
rect 407672 159598 407724 159604
rect 408512 158846 408540 163200
rect 408500 158840 408552 158846
rect 408500 158782 408552 158788
rect 408868 158772 408920 158778
rect 408868 158714 408920 158720
rect 408776 152924 408828 152930
rect 408776 152866 408828 152872
rect 408132 152108 408184 152114
rect 408132 152050 408184 152056
rect 407580 152040 407632 152046
rect 407580 151982 407632 151988
rect 408144 150226 408172 152050
rect 408788 150226 408816 152866
rect 408880 152250 408908 158714
rect 409064 152726 409092 163254
rect 409248 163146 409276 163254
rect 409326 163200 409382 164400
rect 410154 163200 410210 164400
rect 410720 163254 410932 163282
rect 409340 163146 409368 163200
rect 409248 163118 409368 163146
rect 410168 159866 410196 163200
rect 410156 159860 410208 159866
rect 410156 159802 410208 159808
rect 409420 154012 409472 154018
rect 409420 153954 409472 153960
rect 409052 152720 409104 152726
rect 409052 152662 409104 152668
rect 408868 152244 408920 152250
rect 408868 152186 408920 152192
rect 409432 150226 409460 153954
rect 410720 152930 410748 163254
rect 410904 163146 410932 163254
rect 410982 163200 411038 164400
rect 411810 163200 411866 164400
rect 412638 163200 412694 164400
rect 413558 163200 413614 164400
rect 414124 163254 414336 163282
rect 410996 163146 411024 163200
rect 410904 163118 411024 163146
rect 411352 159044 411404 159050
rect 411352 158986 411404 158992
rect 411260 158840 411312 158846
rect 411260 158782 411312 158788
rect 410708 152924 410760 152930
rect 410708 152866 410760 152872
rect 410708 152448 410760 152454
rect 410708 152390 410760 152396
rect 410064 152176 410116 152182
rect 410064 152118 410116 152124
rect 410076 150226 410104 152118
rect 410720 150226 410748 152390
rect 411272 152182 411300 158782
rect 411260 152176 411312 152182
rect 411260 152118 411312 152124
rect 411364 150226 411392 158986
rect 411824 158914 411852 163200
rect 411812 158908 411864 158914
rect 411812 158850 411864 158856
rect 412652 158778 412680 163200
rect 413192 159588 413244 159594
rect 413192 159530 413244 159536
rect 412640 158772 412692 158778
rect 412640 158714 412692 158720
rect 411996 153944 412048 153950
rect 411996 153886 412048 153892
rect 412008 150226 412036 153886
rect 413100 153128 413152 153134
rect 413100 153070 413152 153076
rect 412640 152992 412692 152998
rect 412640 152934 412692 152940
rect 412652 150226 412680 152934
rect 413112 150498 413140 153070
rect 413204 151814 413232 159530
rect 413572 159526 413600 163200
rect 413560 159520 413612 159526
rect 413560 159462 413612 159468
rect 413744 158908 413796 158914
rect 413744 158850 413796 158856
rect 413756 152454 413784 158850
rect 414124 153134 414152 163254
rect 414308 163146 414336 163254
rect 414386 163200 414442 164400
rect 415214 163200 415270 164400
rect 416042 163200 416098 164400
rect 416870 163200 416926 164400
rect 416976 163254 417648 163282
rect 414400 163146 414428 163200
rect 414308 163118 414428 163146
rect 414572 154216 414624 154222
rect 414572 154158 414624 154164
rect 414112 153128 414164 153134
rect 414112 153070 414164 153076
rect 413744 152448 413796 152454
rect 413744 152390 413796 152396
rect 413204 151786 413968 151814
rect 413112 150470 413324 150498
rect 413296 150226 413324 150470
rect 413940 150226 413968 151786
rect 414584 150226 414612 154158
rect 415228 152998 415256 163200
rect 416056 159934 416084 163200
rect 415952 159928 416004 159934
rect 415952 159870 416004 159876
rect 416044 159928 416096 159934
rect 416044 159870 416096 159876
rect 415676 159180 415728 159186
rect 415676 159122 415728 159128
rect 415216 152992 415268 152998
rect 415216 152934 415268 152940
rect 415688 152318 415716 159122
rect 415860 153196 415912 153202
rect 415860 153138 415912 153144
rect 415216 152312 415268 152318
rect 415216 152254 415268 152260
rect 415676 152312 415728 152318
rect 415676 152254 415728 152260
rect 415228 150226 415256 152254
rect 415872 150226 415900 153138
rect 415964 151814 415992 159870
rect 416884 159594 416912 163200
rect 416872 159588 416924 159594
rect 416872 159530 416924 159536
rect 416976 153202 417004 163254
rect 417620 163146 417648 163254
rect 417698 163200 417754 164400
rect 418172 163254 418476 163282
rect 417712 163146 417740 163200
rect 417620 163118 417740 163146
rect 417148 154148 417200 154154
rect 417148 154090 417200 154096
rect 416964 153196 417016 153202
rect 416964 153138 417016 153144
rect 415964 151786 416544 151814
rect 416516 150226 416544 151786
rect 417160 150226 417188 154090
rect 418172 153066 418200 163254
rect 418448 163146 418476 163254
rect 418526 163200 418582 164400
rect 419354 163200 419410 164400
rect 420274 163200 420330 164400
rect 421102 163200 421158 164400
rect 421930 163200 421986 164400
rect 422758 163200 422814 164400
rect 423586 163200 423642 164400
rect 424414 163200 424470 164400
rect 425242 163200 425298 164400
rect 426162 163200 426218 164400
rect 426990 163200 427046 164400
rect 427818 163200 427874 164400
rect 428646 163200 428702 164400
rect 429212 163254 429424 163282
rect 418540 163146 418568 163200
rect 418448 163118 418568 163146
rect 418252 159996 418304 160002
rect 418252 159938 418304 159944
rect 417792 153060 417844 153066
rect 417792 153002 417844 153008
rect 418160 153060 418212 153066
rect 418160 153002 418212 153008
rect 417804 150226 417832 153002
rect 418264 152114 418292 159938
rect 419368 158982 419396 163200
rect 420288 159458 420316 163200
rect 420276 159452 420328 159458
rect 420276 159394 420328 159400
rect 419356 158976 419408 158982
rect 419356 158918 419408 158924
rect 419540 158772 419592 158778
rect 419540 158714 419592 158720
rect 418436 152380 418488 152386
rect 418436 152322 418488 152328
rect 418252 152108 418304 152114
rect 418252 152050 418304 152056
rect 418448 150226 418476 152322
rect 419080 152312 419132 152318
rect 419080 152254 419132 152260
rect 419092 150226 419120 152254
rect 419552 151842 419580 158714
rect 419724 154284 419776 154290
rect 419724 154226 419776 154232
rect 419540 151836 419592 151842
rect 419540 151778 419592 151784
rect 419736 150226 419764 154226
rect 421116 153950 421144 163200
rect 421104 153944 421156 153950
rect 421104 153886 421156 153892
rect 421656 152788 421708 152794
rect 421656 152730 421708 152736
rect 420368 152516 420420 152522
rect 420368 152458 420420 152464
rect 420380 150226 420408 152458
rect 421012 151904 421064 151910
rect 421012 151846 421064 151852
rect 421024 150226 421052 151846
rect 421668 150226 421696 152730
rect 421944 152386 421972 163200
rect 422772 159118 422800 163200
rect 423600 159934 423628 163200
rect 424428 160002 424456 163200
rect 424416 159996 424468 160002
rect 424416 159938 424468 159944
rect 423404 159928 423456 159934
rect 423404 159870 423456 159876
rect 423588 159928 423640 159934
rect 423588 159870 423640 159876
rect 422760 159112 422812 159118
rect 422760 159054 422812 159060
rect 422300 153876 422352 153882
rect 422300 153818 422352 153824
rect 421932 152380 421984 152386
rect 421932 152322 421984 152328
rect 422312 150226 422340 153818
rect 422852 152584 422904 152590
rect 422852 152526 422904 152532
rect 422864 151814 422892 152526
rect 423416 152522 423444 159870
rect 424968 159112 425020 159118
rect 424968 159054 425020 159060
rect 423496 158976 423548 158982
rect 423496 158918 423548 158924
rect 423404 152516 423456 152522
rect 423404 152458 423456 152464
rect 423508 151910 423536 158918
rect 424876 154080 424928 154086
rect 424876 154022 424928 154028
rect 424232 152108 424284 152114
rect 424232 152050 424284 152056
rect 423588 151972 423640 151978
rect 423588 151914 423640 151920
rect 423496 151904 423548 151910
rect 423496 151846 423548 151852
rect 422864 151786 422984 151814
rect 422956 150226 422984 151786
rect 423600 150226 423628 151914
rect 424244 150226 424272 152050
rect 424888 150226 424916 154022
rect 424980 151978 425008 159054
rect 425256 153814 425284 163200
rect 425520 154352 425572 154358
rect 425520 154294 425572 154300
rect 425244 153808 425296 153814
rect 425244 153750 425296 153756
rect 424968 151972 425020 151978
rect 424968 151914 425020 151920
rect 425532 150226 425560 154294
rect 426176 153474 426204 163200
rect 427004 160070 427032 163200
rect 426992 160064 427044 160070
rect 426992 160006 427044 160012
rect 427360 159724 427412 159730
rect 427360 159666 427412 159672
rect 426164 153468 426216 153474
rect 426164 153410 426216 153416
rect 426808 152652 426860 152658
rect 426808 152594 426860 152600
rect 426164 152040 426216 152046
rect 426164 151982 426216 151988
rect 426176 150226 426204 151982
rect 426820 150226 426848 152594
rect 427084 152516 427136 152522
rect 427084 152458 427136 152464
rect 427096 151910 427124 152458
rect 427084 151904 427136 151910
rect 427084 151846 427136 151852
rect 427372 150226 427400 159666
rect 427832 159322 427860 163200
rect 428004 159384 428056 159390
rect 428004 159326 428056 159332
rect 427820 159316 427872 159322
rect 427820 159258 427872 159264
rect 428016 150226 428044 159326
rect 428660 152794 428688 163200
rect 428648 152788 428700 152794
rect 428648 152730 428700 152736
rect 429212 152658 429240 163254
rect 429396 163146 429424 163254
rect 429474 163200 429530 164400
rect 429580 163254 430252 163282
rect 429488 163146 429516 163200
rect 429396 163118 429516 163146
rect 429476 153468 429528 153474
rect 429476 153410 429528 153416
rect 429292 152856 429344 152862
rect 429292 152798 429344 152804
rect 429200 152652 429252 152658
rect 429200 152594 429252 152600
rect 428648 152244 428700 152250
rect 428648 152186 428700 152192
rect 395172 150164 395430 150192
rect 395402 149940 395430 150164
rect 396046 149940 396074 150198
rect 396598 149940 396626 150198
rect 397242 149940 397270 150198
rect 397886 149940 397914 150198
rect 398530 149940 398558 150198
rect 399174 149940 399202 150198
rect 399818 149940 399846 150198
rect 400462 149940 400490 150198
rect 401106 149940 401134 150198
rect 401750 149940 401778 150198
rect 402394 149940 402422 150198
rect 403038 149940 403066 150198
rect 403164 150204 403216 150210
rect 403636 150198 403710 150226
rect 403164 150146 403216 150152
rect 403682 149940 403710 150198
rect 404314 150204 404366 150210
rect 404924 150198 404998 150226
rect 405568 150198 405642 150226
rect 406212 150198 406286 150226
rect 406856 150198 406930 150226
rect 407500 150198 407574 150226
rect 408144 150198 408218 150226
rect 408788 150198 408862 150226
rect 409432 150198 409506 150226
rect 410076 150198 410150 150226
rect 410720 150198 410794 150226
rect 411364 150198 411438 150226
rect 412008 150198 412082 150226
rect 412652 150198 412726 150226
rect 413296 150198 413370 150226
rect 413940 150198 414014 150226
rect 414584 150198 414658 150226
rect 415228 150198 415302 150226
rect 415872 150198 415946 150226
rect 416516 150198 416590 150226
rect 417160 150198 417234 150226
rect 417804 150198 417878 150226
rect 418448 150198 418522 150226
rect 419092 150198 419166 150226
rect 419736 150198 419810 150226
rect 420380 150198 420454 150226
rect 421024 150198 421098 150226
rect 421668 150198 421742 150226
rect 422312 150198 422386 150226
rect 422956 150198 423030 150226
rect 423600 150198 423674 150226
rect 424244 150198 424318 150226
rect 424888 150198 424962 150226
rect 425532 150198 425606 150226
rect 426176 150198 426250 150226
rect 426820 150198 426894 150226
rect 427372 150198 427446 150226
rect 428016 150198 428090 150226
rect 404314 150146 404366 150152
rect 404326 149940 404354 150146
rect 404970 149940 404998 150198
rect 405614 149940 405642 150198
rect 406258 149940 406286 150198
rect 406902 149940 406930 150198
rect 407546 149940 407574 150198
rect 408190 149940 408218 150198
rect 408834 149940 408862 150198
rect 409478 149940 409506 150198
rect 410122 149940 410150 150198
rect 410766 149940 410794 150198
rect 411410 149940 411438 150198
rect 412054 149940 412082 150198
rect 412698 149940 412726 150198
rect 413342 149940 413370 150198
rect 413986 149940 414014 150198
rect 414630 149940 414658 150198
rect 415274 149940 415302 150198
rect 415918 149940 415946 150198
rect 416562 149940 416590 150198
rect 417206 149940 417234 150198
rect 417850 149940 417878 150198
rect 418494 149940 418522 150198
rect 419138 149940 419166 150198
rect 419782 149940 419810 150198
rect 420426 149940 420454 150198
rect 421070 149940 421098 150198
rect 421714 149940 421742 150198
rect 422358 149940 422386 150198
rect 423002 149940 423030 150198
rect 423646 149940 423674 150198
rect 424290 149940 424318 150198
rect 424934 149940 424962 150198
rect 425578 149940 425606 150198
rect 426222 149940 426250 150198
rect 426866 149940 426894 150198
rect 427418 149940 427446 150198
rect 428062 149940 428090 150198
rect 428660 150090 428688 152186
rect 429304 150090 429332 152798
rect 429488 152454 429516 153410
rect 429580 152862 429608 163254
rect 430224 163146 430252 163254
rect 430302 163200 430358 164400
rect 430592 163254 431080 163282
rect 430316 163146 430344 163200
rect 430224 163118 430344 163146
rect 429936 159792 429988 159798
rect 429936 159734 429988 159740
rect 429568 152856 429620 152862
rect 429568 152798 429620 152804
rect 429476 152448 429528 152454
rect 429476 152390 429528 152396
rect 429752 152380 429804 152386
rect 429752 152322 429804 152328
rect 429764 152250 429792 152322
rect 429752 152244 429804 152250
rect 429752 152186 429804 152192
rect 429948 150226 429976 159734
rect 430592 152590 430620 163254
rect 431052 163146 431080 163254
rect 431130 163200 431186 164400
rect 431958 163200 432014 164400
rect 432878 163200 432934 164400
rect 433444 163254 433656 163282
rect 431144 163146 431172 163200
rect 431052 163118 431172 163146
rect 430672 159656 430724 159662
rect 430672 159598 430724 159604
rect 430580 152584 430632 152590
rect 430580 152526 430632 152532
rect 430684 150226 430712 159598
rect 431972 153134 432000 163200
rect 432512 159860 432564 159866
rect 432512 159802 432564 159808
rect 431868 153128 431920 153134
rect 431868 153070 431920 153076
rect 431960 153128 432012 153134
rect 431960 153070 432012 153076
rect 431880 152810 431908 153070
rect 431880 152782 432000 152810
rect 431972 152726 432000 152782
rect 431868 152720 431920 152726
rect 431868 152662 431920 152668
rect 431960 152720 432012 152726
rect 431960 152662 432012 152668
rect 431224 152176 431276 152182
rect 431224 152118 431276 152124
rect 429948 150198 430022 150226
rect 428660 150062 428734 150090
rect 429304 150062 429378 150090
rect 428706 149940 428734 150062
rect 429350 149940 429378 150062
rect 429994 149940 430022 150198
rect 430638 150198 430712 150226
rect 430638 149940 430666 150198
rect 431236 150090 431264 152118
rect 431880 150090 431908 152662
rect 432524 150226 432552 159802
rect 432696 153808 432748 153814
rect 432696 153750 432748 153756
rect 432708 152318 432736 153750
rect 432788 153128 432840 153134
rect 432788 153070 432840 153076
rect 432696 152312 432748 152318
rect 432696 152254 432748 152260
rect 432800 152250 432828 153070
rect 432892 152425 432920 163200
rect 433156 152924 433208 152930
rect 433156 152866 433208 152872
rect 432878 152416 432934 152425
rect 432878 152351 432934 152360
rect 432788 152244 432840 152250
rect 432788 152186 432840 152192
rect 432524 150198 432598 150226
rect 431236 150062 431310 150090
rect 431880 150062 431954 150090
rect 431282 149940 431310 150062
rect 431926 149940 431954 150062
rect 432570 149940 432598 150198
rect 433168 150090 433196 152866
rect 433444 152182 433472 163254
rect 433628 163146 433656 163254
rect 433706 163200 433762 164400
rect 434534 163200 434590 164400
rect 434732 163254 435312 163282
rect 433720 163146 433748 163200
rect 433628 163118 433748 163146
rect 434548 152726 434576 163200
rect 434732 152930 434760 163254
rect 435284 163146 435312 163254
rect 435362 163200 435418 164400
rect 436190 163200 436246 164400
rect 436480 163254 436968 163282
rect 435376 163146 435404 163200
rect 435284 163118 435404 163146
rect 435088 159520 435140 159526
rect 435088 159462 435140 159468
rect 434720 152924 434772 152930
rect 434720 152866 434772 152872
rect 434444 152720 434496 152726
rect 434444 152662 434496 152668
rect 434536 152720 434588 152726
rect 434536 152662 434588 152668
rect 434456 152522 434484 152662
rect 433800 152516 433852 152522
rect 433800 152458 433852 152464
rect 434444 152516 434496 152522
rect 434444 152458 434496 152464
rect 433432 152176 433484 152182
rect 433432 152118 433484 152124
rect 433812 150090 433840 152458
rect 434444 151836 434496 151842
rect 434444 151778 434496 151784
rect 434456 150090 434484 151778
rect 435100 150226 435128 159462
rect 435732 152516 435784 152522
rect 435732 152458 435784 152464
rect 435100 150198 435174 150226
rect 433168 150062 433242 150090
rect 433812 150062 433886 150090
rect 434456 150062 434530 150090
rect 433214 149940 433242 150062
rect 433858 149940 433886 150062
rect 434502 149940 434530 150062
rect 435146 149940 435174 150198
rect 435744 150090 435772 152458
rect 436204 152046 436232 163200
rect 436480 152998 436508 163254
rect 436940 163146 436968 163254
rect 437018 163200 437074 164400
rect 437492 163254 437796 163282
rect 437032 163146 437060 163200
rect 436940 163118 437060 163146
rect 436376 152992 436428 152998
rect 436376 152934 436428 152940
rect 436468 152992 436520 152998
rect 436468 152934 436520 152940
rect 436192 152040 436244 152046
rect 436192 151982 436244 151988
rect 436388 150090 436416 152934
rect 437492 151910 437520 163254
rect 437768 163146 437796 163254
rect 437846 163200 437902 164400
rect 437952 163254 438624 163282
rect 437860 163146 437888 163200
rect 437768 163118 437888 163146
rect 437664 159588 437716 159594
rect 437664 159530 437716 159536
rect 437020 151904 437072 151910
rect 437020 151846 437072 151852
rect 437480 151904 437532 151910
rect 437480 151846 437532 151852
rect 437032 150090 437060 151846
rect 437676 150226 437704 159530
rect 437952 153134 437980 163254
rect 438596 163146 438624 163254
rect 438674 163200 438730 164400
rect 438872 163254 439544 163282
rect 438688 163146 438716 163200
rect 438596 163118 438716 163146
rect 438872 153202 438900 163254
rect 439516 163146 439544 163254
rect 439594 163200 439650 164400
rect 440422 163200 440478 164400
rect 441250 163200 441306 164400
rect 441724 163254 442028 163282
rect 439608 163146 439636 163200
rect 439516 163118 439636 163146
rect 440332 159452 440384 159458
rect 440332 159394 440384 159400
rect 438308 153196 438360 153202
rect 438308 153138 438360 153144
rect 438860 153196 438912 153202
rect 438860 153138 438912 153144
rect 437940 153128 437992 153134
rect 437940 153070 437992 153076
rect 437676 150198 437750 150226
rect 435744 150062 435818 150090
rect 436388 150062 436462 150090
rect 437032 150062 437106 150090
rect 435790 149940 435818 150062
rect 436434 149940 436462 150062
rect 437078 149940 437106 150062
rect 437722 149940 437750 150198
rect 438320 150090 438348 153138
rect 438952 153060 439004 153066
rect 438952 153002 439004 153008
rect 438964 150090 438992 153002
rect 439596 151972 439648 151978
rect 439596 151914 439648 151920
rect 439608 150090 439636 151914
rect 440344 150226 440372 159394
rect 440436 153066 440464 163200
rect 440884 153944 440936 153950
rect 440884 153886 440936 153892
rect 440424 153060 440476 153066
rect 440424 153002 440476 153008
rect 440298 150198 440372 150226
rect 438320 150062 438394 150090
rect 438964 150062 439038 150090
rect 439608 150062 439682 150090
rect 438366 149940 438394 150062
rect 439010 149940 439038 150062
rect 439654 149940 439682 150062
rect 440298 149940 440326 150198
rect 440896 150090 440924 153886
rect 441068 152856 441120 152862
rect 441068 152798 441120 152804
rect 441080 151842 441108 152798
rect 441264 152794 441292 163200
rect 441252 152788 441304 152794
rect 441252 152730 441304 152736
rect 441528 152380 441580 152386
rect 441528 152322 441580 152328
rect 441068 151836 441120 151842
rect 441068 151778 441120 151784
rect 441540 150090 441568 152322
rect 441724 151978 441752 163254
rect 442000 163146 442028 163254
rect 442078 163200 442134 164400
rect 442906 163200 442962 164400
rect 443012 163254 443684 163282
rect 442092 163146 442120 163200
rect 442000 163118 442120 163146
rect 442816 159928 442868 159934
rect 442816 159870 442868 159876
rect 442448 153196 442500 153202
rect 442448 153138 442500 153144
rect 442460 152998 442488 153138
rect 442356 152992 442408 152998
rect 442356 152934 442408 152940
rect 442448 152992 442500 152998
rect 442448 152934 442500 152940
rect 442368 152522 442396 152934
rect 442080 152516 442132 152522
rect 442080 152458 442132 152464
rect 442356 152516 442408 152522
rect 442356 152458 442408 152464
rect 442092 152402 442120 152458
rect 442264 152448 442316 152454
rect 442092 152396 442264 152402
rect 442092 152390 442316 152396
rect 442092 152374 442304 152390
rect 442172 152108 442224 152114
rect 442172 152050 442224 152056
rect 441712 151972 441764 151978
rect 441712 151914 441764 151920
rect 442184 150090 442212 152050
rect 442828 150226 442856 159870
rect 442920 153202 442948 163200
rect 442908 153196 442960 153202
rect 442908 153138 442960 153144
rect 443012 152114 443040 163254
rect 443656 163146 443684 163254
rect 443734 163200 443790 164400
rect 444562 163200 444618 164400
rect 445390 163200 445446 164400
rect 445772 163254 446260 163282
rect 443748 163146 443776 163200
rect 443656 163118 443776 163146
rect 443460 159996 443512 160002
rect 443460 159938 443512 159944
rect 443000 152108 443052 152114
rect 443000 152050 443052 152056
rect 443472 150226 443500 159938
rect 444576 152318 444604 163200
rect 445300 160064 445352 160070
rect 445300 160006 445352 160012
rect 444840 152788 444892 152794
rect 444840 152730 444892 152736
rect 444852 152454 444880 152730
rect 444748 152448 444800 152454
rect 444748 152390 444800 152396
rect 444840 152448 444892 152454
rect 444840 152390 444892 152396
rect 444104 152312 444156 152318
rect 444104 152254 444156 152260
rect 444564 152312 444616 152318
rect 444564 152254 444616 152260
rect 442828 150198 442902 150226
rect 443472 150198 443546 150226
rect 440896 150062 440970 150090
rect 441540 150062 441614 150090
rect 442184 150062 442258 150090
rect 440942 149940 440970 150062
rect 441586 149940 441614 150062
rect 442230 149940 442258 150062
rect 442874 149940 442902 150198
rect 443518 149940 443546 150198
rect 444116 150090 444144 152254
rect 444760 150090 444788 152390
rect 445312 150226 445340 160006
rect 445404 152590 445432 163200
rect 445392 152584 445444 152590
rect 445392 152526 445444 152532
rect 445772 151910 445800 163254
rect 446232 163146 446260 163254
rect 446310 163200 446366 164400
rect 447138 163200 447194 164400
rect 447704 163254 447916 163282
rect 446324 163146 446352 163200
rect 446232 163118 446352 163146
rect 447152 159730 447180 163200
rect 447140 159724 447192 159730
rect 447140 159666 447192 159672
rect 446036 159384 446088 159390
rect 446036 159326 446088 159332
rect 445668 151904 445720 151910
rect 445666 151872 445668 151881
rect 445760 151904 445812 151910
rect 445720 151872 445722 151881
rect 445760 151846 445812 151852
rect 445666 151807 445722 151816
rect 446048 150226 446076 159326
rect 446772 152992 446824 152998
rect 446772 152934 446824 152940
rect 446680 152856 446732 152862
rect 446680 152798 446732 152804
rect 446586 152008 446642 152017
rect 446586 151943 446588 151952
rect 446640 151943 446642 151952
rect 446588 151914 446640 151920
rect 446588 151836 446640 151842
rect 446588 151778 446640 151784
rect 445312 150198 445478 150226
rect 446048 150198 446122 150226
rect 446600 150210 446628 151778
rect 444116 150062 444190 150090
rect 444760 150062 444834 150090
rect 444162 149940 444190 150062
rect 444806 149940 444834 150062
rect 445450 149940 445478 150198
rect 446094 149940 446122 150198
rect 446588 150204 446640 150210
rect 446588 150146 446640 150152
rect 446692 150090 446720 152798
rect 446784 151858 446812 152934
rect 447704 152862 447732 163254
rect 447888 163146 447916 163254
rect 447966 163200 448022 164400
rect 448794 163200 448850 164400
rect 448900 163254 449572 163282
rect 447980 163146 448008 163200
rect 447888 163118 448008 163146
rect 448808 159798 448836 163200
rect 448796 159792 448848 159798
rect 448796 159734 448848 159740
rect 447692 152856 447744 152862
rect 447692 152798 447744 152804
rect 448900 152794 448928 163254
rect 449544 163146 449572 163254
rect 449622 163200 449678 164400
rect 450450 163200 450506 164400
rect 451278 163200 451334 164400
rect 452106 163200 452162 164400
rect 453026 163200 453082 164400
rect 453854 163200 453910 164400
rect 454682 163200 454738 164400
rect 455510 163200 455566 164400
rect 456338 163200 456394 164400
rect 457166 163200 457222 164400
rect 457994 163200 458050 164400
rect 458914 163200 458970 164400
rect 459742 163200 459798 164400
rect 460570 163200 460626 164400
rect 461398 163200 461454 164400
rect 462226 163200 462282 164400
rect 463054 163200 463110 164400
rect 463882 163200 463938 164400
rect 464710 163200 464766 164400
rect 465630 163200 465686 164400
rect 466458 163200 466514 164400
rect 467286 163200 467342 164400
rect 468114 163200 468170 164400
rect 468942 163200 468998 164400
rect 469770 163200 469826 164400
rect 470598 163200 470654 164400
rect 471426 163200 471482 164400
rect 472346 163200 472402 164400
rect 473174 163200 473230 164400
rect 474002 163200 474058 164400
rect 474830 163200 474886 164400
rect 475658 163200 475714 164400
rect 476486 163200 476542 164400
rect 477314 163200 477370 164400
rect 478142 163200 478198 164400
rect 479062 163200 479118 164400
rect 479890 163200 479946 164400
rect 480718 163200 480774 164400
rect 481546 163200 481602 164400
rect 482374 163200 482430 164400
rect 483202 163200 483258 164400
rect 484030 163200 484086 164400
rect 484412 163254 484808 163282
rect 449636 163146 449664 163200
rect 449544 163118 449664 163146
rect 450464 159866 450492 163200
rect 450452 159860 450504 159866
rect 450452 159802 450504 159808
rect 451292 159594 451320 163200
rect 451280 159588 451332 159594
rect 451280 159530 451332 159536
rect 452120 159458 452148 163200
rect 452108 159452 452160 159458
rect 452108 159394 452160 159400
rect 453040 159390 453068 163200
rect 453868 159662 453896 163200
rect 453856 159656 453908 159662
rect 453856 159598 453908 159604
rect 454696 159526 454724 163200
rect 454684 159520 454736 159526
rect 454684 159462 454736 159468
rect 453028 159384 453080 159390
rect 453028 159326 453080 159332
rect 455524 158914 455552 163200
rect 455512 158908 455564 158914
rect 455512 158850 455564 158856
rect 456352 158846 456380 163200
rect 456800 159860 456852 159866
rect 456800 159802 456852 159808
rect 456340 158840 456392 158846
rect 456340 158782 456392 158788
rect 454408 153128 454460 153134
rect 454408 153070 454460 153076
rect 451832 152924 451884 152930
rect 451832 152866 451884 152872
rect 448888 152788 448940 152794
rect 448888 152730 448940 152736
rect 446956 152720 447008 152726
rect 446954 152688 446956 152697
rect 447048 152720 447100 152726
rect 447008 152688 447010 152697
rect 447048 152662 447100 152668
rect 447414 152688 447470 152697
rect 446954 152623 447010 152632
rect 447060 152130 447088 152662
rect 447324 152652 447376 152658
rect 447414 152623 447416 152632
rect 447324 152594 447376 152600
rect 447468 152623 447470 152632
rect 451188 152652 451240 152658
rect 447416 152594 447468 152600
rect 451188 152594 451240 152600
rect 446968 152102 447088 152130
rect 446968 152046 446996 152102
rect 446956 152040 447008 152046
rect 446956 151982 447008 151988
rect 447048 152040 447100 152046
rect 447048 151982 447100 151988
rect 447060 151881 447088 151982
rect 447046 151872 447102 151881
rect 446784 151842 446996 151858
rect 446784 151836 447008 151842
rect 446784 151830 446956 151836
rect 447046 151807 447102 151816
rect 446956 151778 447008 151784
rect 447336 150226 447364 152594
rect 449898 152416 449954 152425
rect 448612 152380 448664 152386
rect 449898 152351 449954 152360
rect 448612 152322 448664 152328
rect 448058 152008 448114 152017
rect 448058 151943 448060 151952
rect 448112 151943 448114 151952
rect 448060 151914 448112 151920
rect 448624 150226 448652 152322
rect 449256 152244 449308 152250
rect 449256 152186 449308 152192
rect 449268 150226 449296 152186
rect 449912 150226 449940 152351
rect 450544 152176 450596 152182
rect 450544 152118 450596 152124
rect 450556 150226 450584 152118
rect 451200 150226 451228 152594
rect 451844 150226 451872 152866
rect 452476 152720 452528 152726
rect 452476 152662 452528 152668
rect 452488 150226 452516 152662
rect 453120 152516 453172 152522
rect 453120 152458 453172 152464
rect 453132 150226 453160 152458
rect 453764 152040 453816 152046
rect 453764 151982 453816 151988
rect 453776 150226 453804 151982
rect 454420 150226 454448 153070
rect 455696 153060 455748 153066
rect 455696 153002 455748 153008
rect 455052 151836 455104 151842
rect 455052 151778 455104 151784
rect 455064 150226 455092 151778
rect 455708 150226 455736 153002
rect 456340 152448 456392 152454
rect 456340 152390 456392 152396
rect 456352 150226 456380 152390
rect 456812 152046 456840 159802
rect 457180 159254 457208 163200
rect 458008 160002 458036 163200
rect 457996 159996 458048 160002
rect 457996 159938 458048 159944
rect 458928 159866 458956 163200
rect 458916 159860 458968 159866
rect 458916 159802 458968 159808
rect 459756 159730 459784 163200
rect 460204 159792 460256 159798
rect 460204 159734 460256 159740
rect 458180 159724 458232 159730
rect 458180 159666 458232 159672
rect 459744 159724 459796 159730
rect 459744 159666 459796 159672
rect 457168 159248 457220 159254
rect 457168 159190 457220 159196
rect 458192 153202 458220 159666
rect 457628 153196 457680 153202
rect 457628 153138 457680 153144
rect 458180 153196 458232 153202
rect 458180 153138 458232 153144
rect 456800 152040 456852 152046
rect 456800 151982 456852 151988
rect 456984 151972 457036 151978
rect 456984 151914 457036 151920
rect 456996 150226 457024 151914
rect 457640 150226 457668 153138
rect 459468 152584 459520 152590
rect 459468 152526 459520 152532
rect 458916 152312 458968 152318
rect 458916 152254 458968 152260
rect 458180 152108 458232 152114
rect 458180 152050 458232 152056
rect 458192 150226 458220 152050
rect 458928 150226 458956 152254
rect 447336 150198 447410 150226
rect 446692 150062 446766 150090
rect 446738 149940 446766 150062
rect 447382 149940 447410 150198
rect 448014 150204 448066 150210
rect 448624 150198 448698 150226
rect 449268 150198 449342 150226
rect 449912 150198 449986 150226
rect 450556 150198 450630 150226
rect 451200 150198 451274 150226
rect 451844 150198 451918 150226
rect 452488 150198 452562 150226
rect 453132 150198 453206 150226
rect 453776 150198 453850 150226
rect 454420 150198 454494 150226
rect 455064 150198 455138 150226
rect 455708 150198 455782 150226
rect 456352 150198 456426 150226
rect 456996 150198 457070 150226
rect 457640 150198 457714 150226
rect 458192 150198 458266 150226
rect 448014 150146 448066 150152
rect 448026 149940 448054 150146
rect 448670 149940 448698 150198
rect 449314 149940 449342 150198
rect 449958 149940 449986 150198
rect 450602 149940 450630 150198
rect 451246 149940 451274 150198
rect 451890 149940 451918 150198
rect 452534 149940 452562 150198
rect 453178 149940 453206 150198
rect 453822 149940 453850 150198
rect 454466 149940 454494 150198
rect 455110 149940 455138 150198
rect 455754 149940 455782 150198
rect 456398 149940 456426 150198
rect 457042 149940 457070 150198
rect 457686 149940 457714 150198
rect 458238 149940 458266 150198
rect 458882 150198 458956 150226
rect 459480 150226 459508 152526
rect 460216 151910 460244 159734
rect 460584 159118 460612 163200
rect 461412 159186 461440 163200
rect 461400 159180 461452 159186
rect 461400 159122 461452 159128
rect 460572 159112 460624 159118
rect 460572 159054 460624 159060
rect 462240 158778 462268 163200
rect 463068 159050 463096 163200
rect 463700 159588 463752 159594
rect 463700 159530 463752 159536
rect 463056 159044 463108 159050
rect 463056 158986 463108 158992
rect 463608 158908 463660 158914
rect 463608 158850 463660 158856
rect 463516 158840 463568 158846
rect 463516 158782 463568 158788
rect 462228 158772 462280 158778
rect 462228 158714 462280 158720
rect 460756 153196 460808 153202
rect 460756 153138 460808 153144
rect 460112 151904 460164 151910
rect 460112 151846 460164 151852
rect 460204 151904 460256 151910
rect 460204 151846 460256 151852
rect 460124 150226 460152 151846
rect 460768 150226 460796 153138
rect 463528 153134 463556 158782
rect 463620 153202 463648 158850
rect 463608 153196 463660 153202
rect 463608 153138 463660 153144
rect 463516 153128 463568 153134
rect 463516 153070 463568 153076
rect 461400 152856 461452 152862
rect 461400 152798 461452 152804
rect 461412 150226 461440 152798
rect 462688 152788 462740 152794
rect 462688 152730 462740 152736
rect 462044 151904 462096 151910
rect 462044 151846 462096 151852
rect 462056 150226 462084 151846
rect 462700 150226 462728 152730
rect 463332 152040 463384 152046
rect 463332 151982 463384 151988
rect 463344 150226 463372 151982
rect 463712 151814 463740 159530
rect 463896 158846 463924 163200
rect 464252 159452 464304 159458
rect 464252 159394 464304 159400
rect 463884 158840 463936 158846
rect 463884 158782 463936 158788
rect 464264 151814 464292 159394
rect 464620 159248 464672 159254
rect 464620 159190 464672 159196
rect 464632 153066 464660 159190
rect 464724 158914 464752 163200
rect 464896 159996 464948 160002
rect 464896 159938 464948 159944
rect 464712 158908 464764 158914
rect 464712 158850 464764 158856
rect 464620 153060 464672 153066
rect 464620 153002 464672 153008
rect 464908 152998 464936 159938
rect 465356 159860 465408 159866
rect 465356 159802 465408 159808
rect 465080 159656 465132 159662
rect 465080 159598 465132 159604
rect 464896 152992 464948 152998
rect 464896 152934 464948 152940
rect 463712 151786 464016 151814
rect 464264 151786 464660 151814
rect 463988 150226 464016 151786
rect 464632 150226 464660 151786
rect 459480 150198 459554 150226
rect 460124 150198 460198 150226
rect 460768 150198 460842 150226
rect 461412 150198 461486 150226
rect 462056 150198 462130 150226
rect 462700 150198 462774 150226
rect 463344 150198 463418 150226
rect 463988 150198 464062 150226
rect 464632 150198 464706 150226
rect 465092 150210 465120 159598
rect 465264 159384 465316 159390
rect 465264 159326 465316 159332
rect 465276 150226 465304 159326
rect 465368 152930 465396 159802
rect 465644 158982 465672 163200
rect 466472 160002 466500 163200
rect 466460 159996 466512 160002
rect 466460 159938 466512 159944
rect 467300 159866 467328 163200
rect 467288 159860 467340 159866
rect 467288 159802 467340 159808
rect 466552 159724 466604 159730
rect 466552 159666 466604 159672
rect 466460 159112 466512 159118
rect 466460 159054 466512 159060
rect 465632 158976 465684 158982
rect 465632 158918 465684 158924
rect 465356 152924 465408 152930
rect 465356 152866 465408 152872
rect 466472 151842 466500 159054
rect 466564 152862 466592 159666
rect 466644 159520 466696 159526
rect 466644 159462 466696 159468
rect 466552 152856 466604 152862
rect 466552 152798 466604 152804
rect 466460 151836 466512 151842
rect 466460 151778 466512 151784
rect 466656 150226 466684 159462
rect 468128 159390 468156 163200
rect 468956 159458 468984 163200
rect 469784 159594 469812 163200
rect 470612 159662 470640 163200
rect 470600 159656 470652 159662
rect 470600 159598 470652 159604
rect 469772 159588 469824 159594
rect 469772 159530 469824 159536
rect 468944 159452 468996 159458
rect 468944 159394 468996 159400
rect 468116 159384 468168 159390
rect 468116 159326 468168 159332
rect 468024 159180 468076 159186
rect 468024 159122 468076 159128
rect 467932 158772 467984 158778
rect 467932 158714 467984 158720
rect 467196 153196 467248 153202
rect 467196 153138 467248 153144
rect 458882 149940 458910 150198
rect 459526 149940 459554 150198
rect 460170 149940 460198 150198
rect 460814 149940 460842 150198
rect 461458 149940 461486 150198
rect 462102 149940 462130 150198
rect 462746 149940 462774 150198
rect 463390 149940 463418 150198
rect 464034 149940 464062 150198
rect 464678 149940 464706 150198
rect 465080 150204 465132 150210
rect 465276 150198 465350 150226
rect 465080 150146 465132 150152
rect 465322 149940 465350 150198
rect 465954 150204 466006 150210
rect 465954 150146 466006 150152
rect 466610 150198 466684 150226
rect 467208 150226 467236 153138
rect 467840 153128 467892 153134
rect 467840 153070 467892 153076
rect 467852 150226 467880 153070
rect 467944 152046 467972 158714
rect 467932 152040 467984 152046
rect 467932 151982 467984 151988
rect 468036 151978 468064 159122
rect 471440 159050 471468 163200
rect 472360 159730 472388 163200
rect 472348 159724 472400 159730
rect 472348 159666 472400 159672
rect 473188 159118 473216 163200
rect 473360 159996 473412 160002
rect 473360 159938 473412 159944
rect 473176 159112 473228 159118
rect 473176 159054 473228 159060
rect 469220 159044 469272 159050
rect 469220 158986 469272 158992
rect 471428 159044 471480 159050
rect 471428 158986 471480 158992
rect 468392 153060 468444 153066
rect 468392 153002 468444 153008
rect 468024 151972 468076 151978
rect 468024 151914 468076 151920
rect 468404 151814 468432 153002
rect 469128 152992 469180 152998
rect 469128 152934 469180 152940
rect 468404 151786 468524 151814
rect 468496 150226 468524 151786
rect 469140 150226 469168 152934
rect 469232 151910 469260 158986
rect 472532 158976 472584 158982
rect 472532 158918 472584 158924
rect 471428 158908 471480 158914
rect 471428 158850 471480 158856
rect 471440 153134 471468 158850
rect 471520 158840 471572 158846
rect 471520 158782 471572 158788
rect 471532 153202 471560 158782
rect 471520 153196 471572 153202
rect 471520 153138 471572 153144
rect 471428 153128 471480 153134
rect 471428 153070 471480 153076
rect 472544 153066 472572 158918
rect 472532 153060 472584 153066
rect 472532 153002 472584 153008
rect 473372 152998 473400 159938
rect 473452 159860 473504 159866
rect 473452 159802 473504 159808
rect 473360 152992 473412 152998
rect 473360 152934 473412 152940
rect 473464 152930 473492 159802
rect 474016 158914 474044 163200
rect 474740 159384 474792 159390
rect 474740 159326 474792 159332
rect 474004 158908 474056 158914
rect 474004 158850 474056 158856
rect 474752 153202 474780 159326
rect 474844 158982 474872 163200
rect 475016 159452 475068 159458
rect 475016 159394 475068 159400
rect 474832 158976 474884 158982
rect 474832 158918 474884 158924
rect 473636 153196 473688 153202
rect 473636 153138 473688 153144
rect 474740 153196 474792 153202
rect 474740 153138 474792 153144
rect 469772 152924 469824 152930
rect 469772 152866 469824 152872
rect 473452 152924 473504 152930
rect 473452 152866 473504 152872
rect 469220 151904 469272 151910
rect 469220 151846 469272 151852
rect 469784 150226 469812 152866
rect 470416 152856 470468 152862
rect 470416 152798 470468 152804
rect 470428 150226 470456 152798
rect 472348 152040 472400 152046
rect 472348 151982 472400 151988
rect 471704 151972 471756 151978
rect 471704 151914 471756 151920
rect 471060 151836 471112 151842
rect 471060 151778 471112 151784
rect 471072 150226 471100 151778
rect 471716 150226 471744 151914
rect 472360 150226 472388 151982
rect 472992 151904 473044 151910
rect 472992 151846 473044 151852
rect 473004 150226 473032 151846
rect 473648 150226 473676 153138
rect 475028 153134 475056 159394
rect 475672 158778 475700 163200
rect 476120 159588 476172 159594
rect 476120 159530 476172 159536
rect 475660 158772 475712 158778
rect 475660 158714 475712 158720
rect 474280 153128 474332 153134
rect 474280 153070 474332 153076
rect 475016 153128 475068 153134
rect 475016 153070 475068 153076
rect 474292 150226 474320 153070
rect 476132 153066 476160 159530
rect 476500 159458 476528 163200
rect 476488 159452 476540 159458
rect 476488 159394 476540 159400
rect 477328 159390 477356 163200
rect 477684 159656 477736 159662
rect 477684 159598 477736 159604
rect 477316 159384 477368 159390
rect 477316 159326 477368 159332
rect 477592 159044 477644 159050
rect 477592 158986 477644 158992
rect 477604 153202 477632 158986
rect 476856 153196 476908 153202
rect 476856 153138 476908 153144
rect 477592 153196 477644 153202
rect 477592 153138 477644 153144
rect 474924 153060 474976 153066
rect 474924 153002 474976 153008
rect 476120 153060 476172 153066
rect 476120 153002 476172 153008
rect 474936 150226 474964 153002
rect 475568 152992 475620 152998
rect 475568 152934 475620 152940
rect 475580 150226 475608 152934
rect 476212 152924 476264 152930
rect 476212 152866 476264 152872
rect 476224 150226 476252 152866
rect 476868 150226 476896 153138
rect 477500 153128 477552 153134
rect 477500 153070 477552 153076
rect 477512 150226 477540 153070
rect 467208 150198 467282 150226
rect 467852 150198 467926 150226
rect 468496 150198 468570 150226
rect 469140 150198 469214 150226
rect 469784 150198 469858 150226
rect 470428 150198 470502 150226
rect 471072 150198 471146 150226
rect 471716 150198 471790 150226
rect 472360 150198 472434 150226
rect 473004 150198 473078 150226
rect 473648 150198 473722 150226
rect 474292 150198 474366 150226
rect 474936 150198 475010 150226
rect 475580 150198 475654 150226
rect 476224 150198 476298 150226
rect 476868 150198 476942 150226
rect 477512 150198 477586 150226
rect 477696 150210 477724 159598
rect 478156 159594 478184 163200
rect 479076 160002 479104 163200
rect 479064 159996 479116 160002
rect 479064 159938 479116 159944
rect 479904 159730 479932 163200
rect 479432 159724 479484 159730
rect 479432 159666 479484 159672
rect 479892 159724 479944 159730
rect 479892 159666 479944 159672
rect 478144 159588 478196 159594
rect 478144 159530 478196 159536
rect 478880 159112 478932 159118
rect 478880 159054 478932 159060
rect 478236 153060 478288 153066
rect 478236 153002 478288 153008
rect 478248 150226 478276 153002
rect 478892 151910 478920 159054
rect 479340 153196 479392 153202
rect 479340 153138 479392 153144
rect 478880 151904 478932 151910
rect 478880 151846 478932 151852
rect 479352 150498 479380 153138
rect 479444 151814 479472 159666
rect 480732 159662 480760 163200
rect 480720 159656 480772 159662
rect 480720 159598 480772 159604
rect 481560 159118 481588 163200
rect 482388 159866 482416 163200
rect 482376 159860 482428 159866
rect 482376 159802 482428 159808
rect 483112 159384 483164 159390
rect 483112 159326 483164 159332
rect 481548 159112 481600 159118
rect 481548 159054 481600 159060
rect 481640 158976 481692 158982
rect 481640 158918 481692 158924
rect 481364 158908 481416 158914
rect 481364 158850 481416 158856
rect 480720 151904 480772 151910
rect 480720 151846 480772 151852
rect 479444 151786 480116 151814
rect 479352 150470 479472 150498
rect 465966 149940 465994 150146
rect 466610 149940 466638 150198
rect 467254 149940 467282 150198
rect 467898 149940 467926 150198
rect 468542 149940 468570 150198
rect 469186 149940 469214 150198
rect 469830 149940 469858 150198
rect 470474 149940 470502 150198
rect 471118 149940 471146 150198
rect 471762 149940 471790 150198
rect 472406 149940 472434 150198
rect 473050 149940 473078 150198
rect 473694 149940 473722 150198
rect 474338 149940 474366 150198
rect 474982 149940 475010 150198
rect 475626 149940 475654 150198
rect 476270 149940 476298 150198
rect 476914 149940 476942 150198
rect 477558 149940 477586 150198
rect 477684 150204 477736 150210
rect 477684 150146 477736 150152
rect 478202 150198 478276 150226
rect 479444 150226 479472 150470
rect 480088 150226 480116 151786
rect 480732 150226 480760 151846
rect 481376 150226 481404 158850
rect 481652 151814 481680 158918
rect 482652 158772 482704 158778
rect 482652 158714 482704 158720
rect 481652 151786 482048 151814
rect 482020 150226 482048 151786
rect 482664 150226 482692 158714
rect 478834 150204 478886 150210
rect 478202 149940 478230 150198
rect 479444 150198 479518 150226
rect 480088 150198 480162 150226
rect 480732 150198 480806 150226
rect 481376 150198 481450 150226
rect 482020 150198 482094 150226
rect 482664 150198 482738 150226
rect 483124 150210 483152 159326
rect 483216 153202 483244 163200
rect 484044 159526 484072 163200
rect 484032 159520 484084 159526
rect 484032 159462 484084 159468
rect 483296 159452 483348 159458
rect 483296 159394 483348 159400
rect 483204 153196 483256 153202
rect 483204 153138 483256 153144
rect 483308 150226 483336 159394
rect 484412 153134 484440 163254
rect 484780 163146 484808 163254
rect 484858 163200 484914 164400
rect 485778 163200 485834 164400
rect 485884 163254 486556 163282
rect 484872 163146 484900 163200
rect 484780 163118 484900 163146
rect 485228 159996 485280 160002
rect 485228 159938 485280 159944
rect 484584 159588 484636 159594
rect 484584 159530 484636 159536
rect 484400 153128 484452 153134
rect 484400 153070 484452 153076
rect 484596 150226 484624 159530
rect 485240 150226 485268 159938
rect 485792 151842 485820 163200
rect 485884 152114 485912 163254
rect 486528 163146 486556 163254
rect 486606 163200 486662 164400
rect 487172 163254 487384 163282
rect 486620 163146 486648 163200
rect 486528 163118 486648 163146
rect 485964 159724 486016 159730
rect 485964 159666 486016 159672
rect 485872 152108 485924 152114
rect 485872 152050 485924 152056
rect 485780 151836 485832 151842
rect 485780 151778 485832 151784
rect 485976 150226 486004 159666
rect 486516 159656 486568 159662
rect 486516 159598 486568 159604
rect 478834 150146 478886 150152
rect 478846 149940 478874 150146
rect 479490 149940 479518 150198
rect 480134 149940 480162 150198
rect 480778 149940 480806 150198
rect 481422 149940 481450 150198
rect 482066 149940 482094 150198
rect 482710 149940 482738 150198
rect 483112 150204 483164 150210
rect 483308 150198 483382 150226
rect 483112 150146 483164 150152
rect 483354 149940 483382 150198
rect 483986 150204 484038 150210
rect 484596 150198 484670 150226
rect 485240 150198 485314 150226
rect 483986 150146 484038 150152
rect 483998 149940 484026 150146
rect 484642 149940 484670 150198
rect 485286 149940 485314 150198
rect 485930 150198 486004 150226
rect 486528 150226 486556 159598
rect 487172 151978 487200 163254
rect 487356 163146 487384 163254
rect 487434 163200 487490 164400
rect 487540 163254 488212 163282
rect 487448 163146 487476 163200
rect 487356 163118 487476 163146
rect 487344 159860 487396 159866
rect 487344 159802 487396 159808
rect 487252 159112 487304 159118
rect 487252 159054 487304 159060
rect 487160 151972 487212 151978
rect 487160 151914 487212 151920
rect 487264 150226 487292 159054
rect 487356 151814 487384 159802
rect 487540 152046 487568 163254
rect 488184 163146 488212 163254
rect 488262 163200 488318 164400
rect 488552 163254 489040 163282
rect 488276 163146 488304 163200
rect 488184 163118 488304 163146
rect 488448 153196 488500 153202
rect 488448 153138 488500 153144
rect 487528 152040 487580 152046
rect 487528 151982 487580 151988
rect 487356 151786 487844 151814
rect 486528 150198 486602 150226
rect 485930 149940 485958 150198
rect 486574 149940 486602 150198
rect 487218 150198 487292 150226
rect 487816 150226 487844 151786
rect 488460 150226 488488 153138
rect 488552 152522 488580 163254
rect 489012 163146 489040 163254
rect 489090 163200 489146 164400
rect 489918 163200 489974 164400
rect 490024 163254 490696 163282
rect 489104 163146 489132 163200
rect 489012 163118 489132 163146
rect 489000 159520 489052 159526
rect 489000 159462 489052 159468
rect 488540 152516 488592 152522
rect 488540 152458 488592 152464
rect 489012 150226 489040 159462
rect 489932 153202 489960 163200
rect 489920 153196 489972 153202
rect 489920 153138 489972 153144
rect 489644 153128 489696 153134
rect 489644 153070 489696 153076
rect 489656 150226 489684 153070
rect 490024 153066 490052 163254
rect 490668 163146 490696 163254
rect 490746 163200 490802 164400
rect 491312 163254 491616 163282
rect 490760 163146 490788 163200
rect 490668 163118 490788 163146
rect 491312 153134 491340 163254
rect 491588 163146 491616 163254
rect 491666 163200 491722 164400
rect 491772 163254 492444 163282
rect 491680 163146 491708 163200
rect 491588 163118 491708 163146
rect 491300 153128 491352 153134
rect 491300 153070 491352 153076
rect 490012 153060 490064 153066
rect 490012 153002 490064 153008
rect 491772 152862 491800 163254
rect 492416 163146 492444 163254
rect 492494 163200 492550 164400
rect 492692 163254 493272 163282
rect 492508 163146 492536 163200
rect 492416 163118 492536 163146
rect 492692 152930 492720 163254
rect 493244 163146 493272 163254
rect 493322 163200 493378 164400
rect 494150 163200 494206 164400
rect 494256 163254 494928 163282
rect 493336 163146 493364 163200
rect 493244 163118 493364 163146
rect 494164 153202 494192 163200
rect 493508 153196 493560 153202
rect 493508 153138 493560 153144
rect 494152 153196 494204 153202
rect 494152 153138 494204 153144
rect 492680 152924 492732 152930
rect 492680 152866 492732 152872
rect 491760 152856 491812 152862
rect 491760 152798 491812 152804
rect 492864 152516 492916 152522
rect 492864 152458 492916 152464
rect 490932 152108 490984 152114
rect 490932 152050 490984 152056
rect 490288 151836 490340 151842
rect 490288 151778 490340 151784
rect 490300 150226 490328 151778
rect 490944 150226 490972 152050
rect 492220 152040 492272 152046
rect 492220 151982 492272 151988
rect 491576 151972 491628 151978
rect 491576 151914 491628 151920
rect 491588 150226 491616 151914
rect 492232 150226 492260 151982
rect 492876 150226 492904 152458
rect 493520 150226 493548 153138
rect 494152 153060 494204 153066
rect 494152 153002 494204 153008
rect 494164 150226 494192 153002
rect 494256 152998 494284 163254
rect 494900 163146 494928 163254
rect 494978 163200 495034 164400
rect 495452 163254 495756 163282
rect 494992 163146 495020 163200
rect 494900 163118 495020 163146
rect 495452 153134 495480 163254
rect 495728 163146 495756 163254
rect 495806 163200 495862 164400
rect 496004 163254 496584 163282
rect 495820 163146 495848 163200
rect 495728 163118 495848 163146
rect 494796 153128 494848 153134
rect 494796 153070 494848 153076
rect 495440 153128 495492 153134
rect 495440 153070 495492 153076
rect 494244 152992 494296 152998
rect 494244 152934 494296 152940
rect 494808 150226 494836 153070
rect 496004 153066 496032 163254
rect 496556 163146 496584 163254
rect 496634 163200 496690 164400
rect 496832 163254 497412 163282
rect 496648 163146 496676 163200
rect 496556 163118 496676 163146
rect 496832 153202 496860 163254
rect 497384 163146 497412 163254
rect 497462 163200 497518 164400
rect 498382 163200 498438 164400
rect 499210 163200 499266 164400
rect 499684 163254 499988 163282
rect 497476 163146 497504 163200
rect 497384 163118 497504 163146
rect 496728 153196 496780 153202
rect 496728 153138 496780 153144
rect 496820 153196 496872 153202
rect 496820 153138 496872 153144
rect 495992 153060 496044 153066
rect 495992 153002 496044 153008
rect 496084 152924 496136 152930
rect 496084 152866 496136 152872
rect 495440 152856 495492 152862
rect 495440 152798 495492 152804
rect 495452 150226 495480 152798
rect 496096 150226 496124 152866
rect 496740 150226 496768 153138
rect 498016 153128 498068 153134
rect 498016 153070 498068 153076
rect 497372 152992 497424 152998
rect 497372 152934 497424 152940
rect 497384 150226 497412 152934
rect 498028 150226 498056 153070
rect 498396 151978 498424 163200
rect 498660 153060 498712 153066
rect 498660 153002 498712 153008
rect 498384 151972 498436 151978
rect 498384 151914 498436 151920
rect 498672 150226 498700 153002
rect 499224 152046 499252 163200
rect 499304 153196 499356 153202
rect 499304 153138 499356 153144
rect 499212 152040 499264 152046
rect 499212 151982 499264 151988
rect 499316 150226 499344 153138
rect 499684 153066 499712 163254
rect 499960 163146 499988 163254
rect 500038 163200 500094 164400
rect 500866 163200 500922 164400
rect 500972 163254 501644 163282
rect 500052 163146 500080 163200
rect 499960 163118 500080 163146
rect 500880 153202 500908 163200
rect 500868 153196 500920 153202
rect 500868 153138 500920 153144
rect 500972 153134 501000 163254
rect 501616 163146 501644 163254
rect 501694 163200 501750 164400
rect 502522 163200 502578 164400
rect 502628 163254 503208 163282
rect 501708 163146 501736 163200
rect 501616 163118 501736 163146
rect 502536 163146 502564 163200
rect 502628 163146 502656 163254
rect 502536 163118 502656 163146
rect 501880 153196 501932 153202
rect 501880 153138 501932 153144
rect 500960 153128 501012 153134
rect 500960 153070 501012 153076
rect 499672 153060 499724 153066
rect 499672 153002 499724 153008
rect 501236 153060 501288 153066
rect 501236 153002 501288 153008
rect 500592 152040 500644 152046
rect 500592 151982 500644 151988
rect 499948 151972 500000 151978
rect 499948 151914 500000 151920
rect 499960 150226 499988 151914
rect 500604 150226 500632 151982
rect 501248 150226 501276 153002
rect 501892 150226 501920 153138
rect 502524 153128 502576 153134
rect 502524 153070 502576 153076
rect 502536 150226 502564 153070
rect 503180 150226 503208 163254
rect 503350 163200 503406 164400
rect 504178 163200 504234 164400
rect 504284 163254 504496 163282
rect 503364 153202 503392 163200
rect 504192 163146 504220 163200
rect 504284 163146 504312 163254
rect 504192 163118 504312 163146
rect 503352 153196 503404 153202
rect 503352 153138 503404 153144
rect 503812 153196 503864 153202
rect 503812 153138 503864 153144
rect 503824 150226 503852 153138
rect 504468 150226 504496 163254
rect 505098 163200 505154 164400
rect 505926 163200 505982 164400
rect 506754 163200 506810 164400
rect 507044 163254 507532 163282
rect 505112 150226 505140 163200
rect 505940 161474 505968 163200
rect 505756 161446 505968 161474
rect 505284 158772 505336 158778
rect 505284 158714 505336 158720
rect 487816 150198 487890 150226
rect 488460 150198 488534 150226
rect 489012 150198 489086 150226
rect 489656 150198 489730 150226
rect 490300 150198 490374 150226
rect 490944 150198 491018 150226
rect 491588 150198 491662 150226
rect 492232 150198 492306 150226
rect 492876 150198 492950 150226
rect 493520 150198 493594 150226
rect 494164 150198 494238 150226
rect 494808 150198 494882 150226
rect 495452 150198 495526 150226
rect 496096 150198 496170 150226
rect 496740 150198 496814 150226
rect 497384 150198 497458 150226
rect 498028 150198 498102 150226
rect 498672 150198 498746 150226
rect 499316 150198 499390 150226
rect 499960 150198 500034 150226
rect 500604 150198 500678 150226
rect 501248 150198 501322 150226
rect 501892 150198 501966 150226
rect 502536 150198 502610 150226
rect 503180 150198 503254 150226
rect 503824 150198 503898 150226
rect 504468 150198 504542 150226
rect 505112 150198 505186 150226
rect 505296 150210 505324 158714
rect 505756 150226 505784 161446
rect 506572 158976 506624 158982
rect 506572 158918 506624 158924
rect 487218 149940 487246 150198
rect 487862 149940 487890 150198
rect 488506 149940 488534 150198
rect 489058 149940 489086 150198
rect 489702 149940 489730 150198
rect 490346 149940 490374 150198
rect 490990 149940 491018 150198
rect 491634 149940 491662 150198
rect 492278 149940 492306 150198
rect 492922 149940 492950 150198
rect 493566 149940 493594 150198
rect 494210 149940 494238 150198
rect 494854 149940 494882 150198
rect 495498 149940 495526 150198
rect 496142 149940 496170 150198
rect 496786 149940 496814 150198
rect 497430 149940 497458 150198
rect 498074 149940 498102 150198
rect 498718 149940 498746 150198
rect 499362 149940 499390 150198
rect 500006 149940 500034 150198
rect 500650 149940 500678 150198
rect 501294 149940 501322 150198
rect 501938 149940 501966 150198
rect 502582 149940 502610 150198
rect 503226 149940 503254 150198
rect 503870 149940 503898 150198
rect 504514 149940 504542 150198
rect 505158 149940 505186 150198
rect 505284 150204 505336 150210
rect 505756 150198 505830 150226
rect 506584 150210 506612 158918
rect 506768 158778 506796 163200
rect 506756 158772 506808 158778
rect 506756 158714 506808 158720
rect 507044 150226 507072 163254
rect 507504 163146 507532 163254
rect 507582 163200 507638 164400
rect 508410 163200 508466 164400
rect 509238 163200 509294 164400
rect 510066 163200 510122 164400
rect 510894 163200 510950 164400
rect 511814 163200 511870 164400
rect 512642 163200 512698 164400
rect 513470 163200 513526 164400
rect 514298 163200 514354 164400
rect 515126 163200 515182 164400
rect 515954 163200 516010 164400
rect 516152 163254 516732 163282
rect 507596 163146 507624 163200
rect 507504 163118 507624 163146
rect 508424 158982 508452 163200
rect 508412 158976 508464 158982
rect 508412 158918 508464 158924
rect 509252 158914 509280 163200
rect 508320 158908 508372 158914
rect 508320 158850 508372 158856
rect 509240 158908 509292 158914
rect 509240 158850 509292 158856
rect 509332 158908 509384 158914
rect 509332 158850 509384 158856
rect 507952 158840 508004 158846
rect 507952 158782 508004 158788
rect 505284 150146 505336 150152
rect 505802 149940 505830 150198
rect 506434 150204 506486 150210
rect 506434 150146 506486 150152
rect 506572 150204 506624 150210
rect 507044 150198 507118 150226
rect 507964 150210 507992 158782
rect 508332 150226 508360 158850
rect 506572 150146 506624 150152
rect 506446 149940 506474 150146
rect 507090 149940 507118 150198
rect 507722 150204 507774 150210
rect 507722 150146 507774 150152
rect 507952 150204 508004 150210
rect 508332 150198 508406 150226
rect 509344 150210 509372 158850
rect 510080 158846 510108 163200
rect 510068 158840 510120 158846
rect 510068 158782 510120 158788
rect 510908 158778 510936 163200
rect 511828 158914 511856 163200
rect 511816 158908 511868 158914
rect 511816 158850 511868 158856
rect 512184 158840 512236 158846
rect 512184 158782 512236 158788
rect 509608 158772 509660 158778
rect 509608 158714 509660 158720
rect 510896 158772 510948 158778
rect 510896 158714 510948 158720
rect 510988 158772 511040 158778
rect 510988 158714 511040 158720
rect 509620 150226 509648 158714
rect 511000 150226 511028 158714
rect 511632 153196 511684 153202
rect 511632 153138 511684 153144
rect 511644 150226 511672 153138
rect 507952 150146 508004 150152
rect 507734 149940 507762 150146
rect 508378 149940 508406 150198
rect 509010 150204 509062 150210
rect 509010 150146 509062 150152
rect 509332 150204 509384 150210
rect 509620 150198 509694 150226
rect 509332 150146 509384 150152
rect 509022 149940 509050 150146
rect 509666 149940 509694 150198
rect 510298 150204 510350 150210
rect 510298 150146 510350 150152
rect 510954 150198 511028 150226
rect 511598 150198 511672 150226
rect 512196 150226 512224 158782
rect 512656 158778 512684 163200
rect 512644 158772 512696 158778
rect 512644 158714 512696 158720
rect 513484 153202 513512 163200
rect 514312 158846 514340 163200
rect 515036 158908 515088 158914
rect 515036 158850 515088 158856
rect 514300 158840 514352 158846
rect 514300 158782 514352 158788
rect 514852 158840 514904 158846
rect 514852 158782 514904 158788
rect 513564 158772 513616 158778
rect 513564 158714 513616 158720
rect 513472 153196 513524 153202
rect 513472 153138 513524 153144
rect 512920 153128 512972 153134
rect 512920 153070 512972 153076
rect 512932 150226 512960 153070
rect 513576 150226 513604 158714
rect 514208 153196 514260 153202
rect 514208 153138 514260 153144
rect 514220 150226 514248 153138
rect 514864 150226 514892 158782
rect 515048 151814 515076 158850
rect 515140 153134 515168 163200
rect 515968 158778 515996 163200
rect 515956 158772 516008 158778
rect 515956 158714 516008 158720
rect 516152 153202 516180 163254
rect 516704 163146 516732 163254
rect 516782 163200 516838 164400
rect 517610 163200 517666 164400
rect 518530 163200 518586 164400
rect 519004 163254 519308 163282
rect 516796 163146 516824 163200
rect 516704 163118 516824 163146
rect 516692 158976 516744 158982
rect 516692 158918 516744 158924
rect 516140 153196 516192 153202
rect 516140 153138 516192 153144
rect 515128 153128 515180 153134
rect 515128 153070 515180 153076
rect 516048 151972 516100 151978
rect 516048 151914 516100 151920
rect 515048 151786 515444 151814
rect 512196 150198 512270 150226
rect 510310 149940 510338 150146
rect 510954 149940 510982 150198
rect 511598 149940 511626 150198
rect 512242 149940 512270 150198
rect 512886 150198 512960 150226
rect 513530 150198 513604 150226
rect 514174 150198 514248 150226
rect 514818 150198 514892 150226
rect 515416 150226 515444 151786
rect 516060 150226 516088 151914
rect 516704 150226 516732 158918
rect 517624 158846 517652 163200
rect 518544 158914 518572 163200
rect 518808 159452 518860 159458
rect 518808 159394 518860 159400
rect 518716 159384 518768 159390
rect 518716 159326 518768 159332
rect 518532 158908 518584 158914
rect 518532 158850 518584 158856
rect 517612 158840 517664 158846
rect 517612 158782 517664 158788
rect 517428 151904 517480 151910
rect 517428 151846 517480 151852
rect 517440 150226 517468 151846
rect 518728 150226 518756 159326
rect 515416 150198 515490 150226
rect 516060 150198 516134 150226
rect 516704 150198 516778 150226
rect 512886 149940 512914 150198
rect 513530 149940 513558 150198
rect 514174 149940 514202 150198
rect 514818 149940 514846 150198
rect 515462 149940 515490 150198
rect 516106 149940 516134 150198
rect 516750 149940 516778 150198
rect 517394 150198 517468 150226
rect 518026 150204 518078 150210
rect 517394 149940 517422 150198
rect 518026 150146 518078 150152
rect 518682 150198 518756 150226
rect 518820 150210 518848 159394
rect 519004 151978 519032 163254
rect 519280 163146 519308 163254
rect 519358 163200 519414 164400
rect 520186 163200 520242 164400
rect 520292 163254 520964 163282
rect 519372 163146 519400 163200
rect 519280 163118 519400 163146
rect 519726 163160 519782 163169
rect 519726 163095 519782 163104
rect 519542 161664 519598 161673
rect 519542 161599 519598 161608
rect 519450 154048 519506 154057
rect 519450 153983 519506 153992
rect 518992 151972 519044 151978
rect 518992 151914 519044 151920
rect 518808 150204 518860 150210
rect 518038 149940 518066 150146
rect 518682 149940 518710 150198
rect 518808 150146 518860 150152
rect 519174 141944 519230 141953
rect 519174 141879 519230 141888
rect 519188 130257 519216 141879
rect 519464 141137 519492 153983
rect 519556 147937 519584 161599
rect 519634 160168 519690 160177
rect 519634 160103 519690 160112
rect 519542 147928 519598 147937
rect 519542 147863 519598 147872
rect 519648 146577 519676 160103
rect 519740 149297 519768 163095
rect 520200 158982 520228 163200
rect 520188 158976 520240 158982
rect 520188 158918 520240 158924
rect 520002 158672 520058 158681
rect 520002 158607 520058 158616
rect 519910 157176 519966 157185
rect 519910 157111 519966 157120
rect 519818 155680 519874 155689
rect 519818 155615 519874 155624
rect 519726 149288 519782 149297
rect 519726 149223 519782 149232
rect 519726 148064 519782 148073
rect 519726 147999 519782 148008
rect 519634 146568 519690 146577
rect 519634 146503 519690 146512
rect 519542 144936 519598 144945
rect 519542 144871 519598 144880
rect 519450 141128 519506 141137
rect 519450 141063 519506 141072
rect 519266 140448 519322 140457
rect 519266 140383 519322 140392
rect 519174 130248 519230 130257
rect 519174 130183 519230 130192
rect 519280 128897 519308 140383
rect 519358 138952 519414 138961
rect 519358 138887 519414 138896
rect 519266 128888 519322 128897
rect 519266 128823 519322 128832
rect 519174 128344 519230 128353
rect 519174 128279 519230 128288
rect 117228 118040 117280 118046
rect 519188 118017 519216 128279
rect 519372 127537 519400 138887
rect 519450 137456 519506 137465
rect 519450 137391 519506 137400
rect 519358 127528 519414 127537
rect 519358 127463 519414 127472
rect 519266 126712 519322 126721
rect 519266 126647 519322 126656
rect 117228 117982 117280 117988
rect 519174 118008 519230 118017
rect 519174 117943 519230 117952
rect 519280 116657 519308 126647
rect 519464 126177 519492 137391
rect 519556 132977 519584 144871
rect 519740 135697 519768 147999
rect 519832 142497 519860 155615
rect 519924 143857 519952 157111
rect 520016 145217 520044 158607
rect 520292 151910 520320 163254
rect 520936 163146 520964 163254
rect 521014 163200 521070 164400
rect 521842 163200 521898 164400
rect 522670 163200 522726 164400
rect 523498 163200 523554 164400
rect 521028 163146 521056 163200
rect 520936 163118 521056 163146
rect 521856 159458 521884 163200
rect 521844 159452 521896 159458
rect 521844 159394 521896 159400
rect 522684 159390 522712 163200
rect 522672 159384 522724 159390
rect 522672 159326 522724 159332
rect 523512 156670 523540 163200
rect 521844 156664 521896 156670
rect 521844 156606 521896 156612
rect 523500 156664 523552 156670
rect 523500 156606 523552 156612
rect 521014 152552 521070 152561
rect 521014 152487 521070 152496
rect 520280 151904 520332 151910
rect 520280 151846 520332 151852
rect 520186 151056 520242 151065
rect 520186 150991 520242 151000
rect 520094 149560 520150 149569
rect 520094 149495 520150 149504
rect 520002 145208 520058 145217
rect 520002 145143 520058 145152
rect 519910 143848 519966 143857
rect 519910 143783 519966 143792
rect 520002 143440 520058 143449
rect 520002 143375 520058 143384
rect 519818 142488 519874 142497
rect 519818 142423 519874 142432
rect 519910 135824 519966 135833
rect 519910 135759 519966 135768
rect 519726 135688 519782 135697
rect 519726 135623 519782 135632
rect 519818 134328 519874 134337
rect 519818 134263 519874 134272
rect 519542 132968 519598 132977
rect 519542 132903 519598 132912
rect 519726 132832 519782 132841
rect 519726 132767 519782 132776
rect 519634 131336 519690 131345
rect 519634 131271 519690 131280
rect 519542 129840 519598 129849
rect 519542 129775 519598 129784
rect 519450 126168 519506 126177
rect 519450 126103 519506 126112
rect 519556 119377 519584 129775
rect 519648 120737 519676 131271
rect 519740 122097 519768 132767
rect 519832 123457 519860 134263
rect 519924 124817 519952 135759
rect 520016 131617 520044 143375
rect 520108 137057 520136 149495
rect 520200 138417 520228 150991
rect 520922 146568 520978 146577
rect 520922 146503 520978 146512
rect 520186 138408 520242 138417
rect 520186 138343 520242 138352
rect 520094 137048 520150 137057
rect 520094 136983 520150 136992
rect 520936 134473 520964 146503
rect 521028 139777 521056 152487
rect 521014 139768 521070 139777
rect 521014 139703 521070 139712
rect 520922 134464 520978 134473
rect 520922 134399 520978 134408
rect 520002 131608 520058 131617
rect 520002 131543 520058 131552
rect 520186 125216 520242 125225
rect 520186 125151 520242 125160
rect 519910 124808 519966 124817
rect 519910 124743 519966 124752
rect 520094 123720 520150 123729
rect 520094 123655 520150 123664
rect 519818 123448 519874 123457
rect 519818 123383 519874 123392
rect 519910 122224 519966 122233
rect 519910 122159 519966 122168
rect 519726 122088 519782 122097
rect 519726 122023 519782 122032
rect 519634 120728 519690 120737
rect 519634 120663 519690 120672
rect 519818 120728 519874 120737
rect 519818 120663 519874 120672
rect 519542 119368 519598 119377
rect 519542 119303 519598 119312
rect 519726 119232 519782 119241
rect 519726 119167 519782 119176
rect 519266 116648 519322 116657
rect 519266 116583 519322 116592
rect 519634 116104 519690 116113
rect 519634 116039 519690 116048
rect 519542 114608 519598 114617
rect 519542 114543 519598 114552
rect 519556 105777 519584 114543
rect 519648 107137 519676 116039
rect 519740 109857 519768 119167
rect 519832 111217 519860 120663
rect 519924 112577 519952 122159
rect 520002 117600 520058 117609
rect 520002 117535 520058 117544
rect 519910 112568 519966 112577
rect 519910 112503 519966 112512
rect 519818 111208 519874 111217
rect 519818 111143 519874 111152
rect 519726 109848 519782 109857
rect 519726 109783 519782 109792
rect 520016 108497 520044 117535
rect 520108 113937 520136 123655
rect 520200 115297 520228 125151
rect 520186 115288 520242 115297
rect 520186 115223 520242 115232
rect 520094 113928 520150 113937
rect 520094 113863 520150 113872
rect 520922 113112 520978 113121
rect 520922 113047 520978 113056
rect 520002 108488 520058 108497
rect 520002 108423 520058 108432
rect 519634 107128 519690 107137
rect 519634 107063 519690 107072
rect 519542 105768 519598 105777
rect 519542 105703 519598 105712
rect 520278 105496 520334 105505
rect 520278 105431 520334 105440
rect 117134 104816 117190 104825
rect 117134 104751 117190 104760
rect 117042 101008 117098 101017
rect 117042 100943 117098 100952
rect 519818 99376 519874 99385
rect 519818 99311 519874 99320
rect 116858 99104 116914 99113
rect 116858 99039 116914 99048
rect 519726 97880 519782 97889
rect 519726 97815 519782 97824
rect 116766 97200 116822 97209
rect 116766 97135 116822 97144
rect 116674 95296 116730 95305
rect 116674 95231 116730 95240
rect 116582 93392 116638 93401
rect 116582 93327 116638 93336
rect 116124 92472 116176 92478
rect 116124 92414 116176 92420
rect 116136 91361 116164 92414
rect 116122 91352 116178 91361
rect 116122 91287 116178 91296
rect 519740 90817 519768 97815
rect 519832 92177 519860 99311
rect 520292 97617 520320 105431
rect 520936 104417 520964 113047
rect 521290 111616 521346 111625
rect 521290 111551 521346 111560
rect 521198 106992 521254 107001
rect 521198 106927 521254 106936
rect 520922 104408 520978 104417
rect 520922 104343 520978 104352
rect 521106 104000 521162 104009
rect 521106 103935 521162 103944
rect 521014 102504 521070 102513
rect 521014 102439 521070 102448
rect 520278 97608 520334 97617
rect 520278 97543 520334 97552
rect 520002 96384 520058 96393
rect 520002 96319 520058 96328
rect 519910 94888 519966 94897
rect 519910 94823 519966 94832
rect 519818 92168 519874 92177
rect 519818 92103 519874 92112
rect 519726 90808 519782 90817
rect 519726 90743 519782 90752
rect 116124 89684 116176 89690
rect 116124 89626 116176 89632
rect 116136 89457 116164 89626
rect 116122 89448 116178 89457
rect 116122 89383 116178 89392
rect 116032 88324 116084 88330
rect 116032 88266 116084 88272
rect 116044 87553 116072 88266
rect 519924 88097 519952 94823
rect 520016 89457 520044 96319
rect 521028 95033 521056 102439
rect 521120 96257 521148 103935
rect 521212 98977 521240 106927
rect 521304 103057 521332 111551
rect 521474 110120 521530 110129
rect 521474 110055 521530 110064
rect 521382 108488 521438 108497
rect 521382 108423 521438 108432
rect 521290 103048 521346 103057
rect 521290 102983 521346 102992
rect 521290 101008 521346 101017
rect 521290 100943 521346 100952
rect 521198 98968 521254 98977
rect 521198 98903 521254 98912
rect 521106 96248 521162 96257
rect 521106 96183 521162 96192
rect 521014 95024 521070 95033
rect 521014 94959 521070 94968
rect 521304 93537 521332 100943
rect 521396 100337 521424 108423
rect 521488 101697 521516 110055
rect 521474 101688 521530 101697
rect 521474 101623 521530 101632
rect 521382 100328 521438 100337
rect 521382 100263 521438 100272
rect 521856 93854 521884 156606
rect 521672 93826 521884 93854
rect 521290 93528 521346 93537
rect 521290 93463 521346 93472
rect 520370 93392 520426 93401
rect 520370 93327 520426 93336
rect 520002 89448 520058 89457
rect 520002 89383 520058 89392
rect 519910 88088 519966 88097
rect 519910 88023 519966 88032
rect 116030 87544 116086 87553
rect 116030 87479 116086 87488
rect 520278 85776 520334 85785
rect 520278 85711 520334 85720
rect 115202 85640 115258 85649
rect 115202 85575 115258 85584
rect 116584 83972 116636 83978
rect 116584 83914 116636 83920
rect 116596 83745 116624 83914
rect 116582 83736 116638 83745
rect 116582 83671 116638 83680
rect 116216 82816 116268 82822
rect 116216 82758 116268 82764
rect 519910 82784 519966 82793
rect 116228 81841 116256 82758
rect 519910 82719 519966 82728
rect 116214 81832 116270 81841
rect 116214 81767 116270 81776
rect 519634 81152 519690 81161
rect 519634 81087 519690 81096
rect 115940 80028 115992 80034
rect 115940 79970 115992 79976
rect 115952 79937 115980 79970
rect 115938 79928 115994 79937
rect 115938 79863 115994 79872
rect 114192 78668 114244 78674
rect 114192 78610 114244 78616
rect 116124 78668 116176 78674
rect 116124 78610 116176 78616
rect 116136 78033 116164 78610
rect 116122 78024 116178 78033
rect 116122 77959 116178 77968
rect 519648 74633 519676 81087
rect 519924 75993 519952 82719
rect 520186 79656 520242 79665
rect 520186 79591 520242 79600
rect 520094 78160 520150 78169
rect 520094 78095 520150 78104
rect 520002 76664 520058 76673
rect 520002 76599 520058 76608
rect 519910 75984 519966 75993
rect 519910 75919 519966 75928
rect 519910 75168 519966 75177
rect 519910 75103 519966 75112
rect 519634 74624 519690 74633
rect 519634 74559 519690 74568
rect 116674 74080 116730 74089
rect 116674 74015 116730 74024
rect 116582 72176 116638 72185
rect 116582 72111 116638 72120
rect 116596 71806 116624 72111
rect 114192 71800 114244 71806
rect 114192 71742 114244 71748
rect 116584 71800 116636 71806
rect 116584 71742 116636 71748
rect 114100 69080 114152 69086
rect 114100 69022 114152 69028
rect 114008 67652 114060 67658
rect 114008 67594 114060 67600
rect 113916 66292 113968 66298
rect 113916 66234 113968 66240
rect 113364 64728 113416 64734
rect 113364 64670 113416 64676
rect 113376 64569 113404 64670
rect 113362 64560 113418 64569
rect 113362 64495 113418 64504
rect 113824 63572 113876 63578
rect 113824 63514 113876 63520
rect 112444 62144 112496 62150
rect 112444 62086 112496 62092
rect 110326 53952 110382 53961
rect 109696 53910 110326 53938
rect 109696 12434 109724 53910
rect 110326 53887 110382 53896
rect 110326 52592 110382 52601
rect 110326 52527 110382 52536
rect 110340 51218 110368 52527
rect 110340 51190 110460 51218
rect 110326 51096 110382 51105
rect 109512 12406 109724 12434
rect 109788 51054 110326 51082
rect 109512 8242 109540 12406
rect 109512 8214 109632 8242
rect 109604 7834 109632 8214
rect 109788 8106 109816 51054
rect 110326 51031 110382 51040
rect 110432 50946 110460 51190
rect 109512 7806 109632 7834
rect 109696 8078 109816 8106
rect 109880 50918 110460 50946
rect 109512 3641 109540 7806
rect 109696 7562 109724 8078
rect 109604 7534 109724 7562
rect 109498 3632 109554 3641
rect 109498 3567 109554 3576
rect 109498 3496 109554 3505
rect 109498 3431 109554 3440
rect 109406 2816 109462 2825
rect 109406 2751 109462 2760
rect 32402 2680 32458 2689
rect 36358 2680 36414 2689
rect 36018 2638 36358 2666
rect 32402 2615 32458 2624
rect 36358 2615 36414 2624
rect 62394 2680 62450 2689
rect 62394 2615 62450 2624
rect 64142 2680 64198 2689
rect 64142 2615 64198 2624
rect 65338 2680 65394 2689
rect 65338 2615 65394 2624
rect 68006 2680 68062 2689
rect 68006 2615 68062 2624
rect 68558 2680 68614 2689
rect 68558 2615 68614 2624
rect 68834 2680 68890 2689
rect 68834 2615 68890 2624
rect 69386 2680 69442 2689
rect 69386 2615 69442 2624
rect 77022 2680 77078 2689
rect 77252 2680 77308 2689
rect 77022 2615 77078 2624
rect 77128 2638 77252 2666
rect 29550 2408 29606 2417
rect 29302 2366 29550 2394
rect 29550 2343 29606 2352
rect 26054 2272 26110 2281
rect 25990 2230 26054 2258
rect 26054 2207 26110 2216
rect 22926 2136 22982 2145
rect 2700 1358 2728 2108
rect 6012 1737 6040 2108
rect 5998 1728 6054 1737
rect 5998 1663 6054 1672
rect 9324 1465 9352 2108
rect 12636 1601 12664 2108
rect 15948 1873 15976 2108
rect 19366 2094 19656 2122
rect 22678 2094 22926 2122
rect 19628 2009 19656 2094
rect 22926 2071 22982 2080
rect 19614 2000 19670 2009
rect 19614 1935 19670 1944
rect 15934 1864 15990 1873
rect 15934 1799 15990 1808
rect 12622 1592 12678 1601
rect 12622 1527 12678 1536
rect 9310 1456 9366 1465
rect 9310 1391 9366 1400
rect 2688 1352 2740 1358
rect 2688 1294 2740 1300
rect 32416 762 32444 2615
rect 33046 2544 33102 2553
rect 32706 2502 33046 2530
rect 33046 2479 33102 2488
rect 39316 1290 39344 2108
rect 42628 1494 42656 2108
rect 42616 1488 42668 1494
rect 42616 1430 42668 1436
rect 46032 1426 46060 2108
rect 46020 1420 46072 1426
rect 46020 1362 46072 1368
rect 39304 1284 39356 1290
rect 39304 1226 39356 1232
rect 49344 1222 49372 2108
rect 49332 1216 49384 1222
rect 49332 1158 49384 1164
rect 52656 1154 52684 2108
rect 52644 1148 52696 1154
rect 52644 1090 52696 1096
rect 55968 1086 55996 2108
rect 59372 1630 59400 2108
rect 62408 1902 62436 2615
rect 62396 1896 62448 1902
rect 62396 1838 62448 1844
rect 62684 1766 62712 2108
rect 64156 1834 64184 2615
rect 65352 1902 65380 2615
rect 65340 1896 65392 1902
rect 65340 1838 65392 1844
rect 64144 1828 64196 1834
rect 64144 1770 64196 1776
rect 62672 1760 62724 1766
rect 62672 1702 62724 1708
rect 59360 1624 59412 1630
rect 59360 1566 59412 1572
rect 55956 1080 56008 1086
rect 55956 1022 56008 1028
rect 65996 1018 66024 2108
rect 68020 1902 68048 2615
rect 68008 1896 68060 1902
rect 68008 1838 68060 1844
rect 68572 1630 68600 2615
rect 68848 1766 68876 2615
rect 68836 1760 68888 1766
rect 68836 1702 68888 1708
rect 69308 1698 69336 2108
rect 69400 1834 69428 2615
rect 69388 1828 69440 1834
rect 69388 1770 69440 1776
rect 69296 1692 69348 1698
rect 69296 1634 69348 1640
rect 68560 1624 68612 1630
rect 68560 1566 68612 1572
rect 72712 1562 72740 2108
rect 72700 1556 72752 1562
rect 72700 1498 72752 1504
rect 65984 1012 66036 1018
rect 65984 954 66036 960
rect 76024 950 76052 2108
rect 77036 1834 77064 2615
rect 77128 1902 77156 2638
rect 77252 2615 77308 2624
rect 77758 2680 77814 2689
rect 77758 2615 77814 2624
rect 77942 2680 77998 2689
rect 77942 2615 77998 2624
rect 78126 2680 78182 2689
rect 78126 2615 78182 2624
rect 78310 2680 78366 2689
rect 78310 2615 78366 2624
rect 95698 2680 95754 2689
rect 96342 2680 96398 2689
rect 96002 2638 96342 2666
rect 95698 2615 95754 2624
rect 96342 2615 96398 2624
rect 103702 2680 103758 2689
rect 103702 2615 103758 2624
rect 104346 2680 104402 2689
rect 104346 2615 104402 2624
rect 105082 2680 105138 2689
rect 105082 2615 105138 2624
rect 106278 2680 106334 2689
rect 107612 2680 107668 2689
rect 106278 2615 106334 2624
rect 107120 2638 107612 2666
rect 77772 1902 77800 2615
rect 77116 1896 77168 1902
rect 77116 1838 77168 1844
rect 77760 1896 77812 1902
rect 77760 1838 77812 1844
rect 77024 1828 77076 1834
rect 77024 1770 77076 1776
rect 77956 1766 77984 2615
rect 77944 1760 77996 1766
rect 77944 1702 77996 1708
rect 78140 1494 78168 2615
rect 78324 1766 78352 2615
rect 95712 2145 95740 2615
rect 96618 2544 96674 2553
rect 96618 2479 96674 2488
rect 97262 2544 97318 2553
rect 97262 2479 97318 2488
rect 94870 2136 94926 2145
rect 78312 1760 78364 1766
rect 78312 1702 78364 1708
rect 79336 1630 79364 2108
rect 82648 1766 82676 2108
rect 86052 1834 86080 2108
rect 89364 1902 89392 2108
rect 88340 1896 88392 1902
rect 88340 1838 88392 1844
rect 89352 1896 89404 1902
rect 89352 1838 89404 1844
rect 85948 1828 86000 1834
rect 85948 1770 86000 1776
rect 86040 1828 86092 1834
rect 86040 1770 86092 1776
rect 82636 1760 82688 1766
rect 82636 1702 82688 1708
rect 79324 1624 79376 1630
rect 79324 1566 79376 1572
rect 78128 1488 78180 1494
rect 78128 1430 78180 1436
rect 85960 1329 85988 1770
rect 85946 1320 86002 1329
rect 85946 1255 86002 1264
rect 88352 1193 88380 1838
rect 88338 1184 88394 1193
rect 88338 1119 88394 1128
rect 76012 944 76064 950
rect 32692 870 32812 898
rect 76012 886 76064 892
rect 32692 762 32720 870
rect 32784 800 32812 870
rect 92676 814 92704 2108
rect 94870 2071 94926 2080
rect 95698 2136 95754 2145
rect 95698 2071 95754 2080
rect 94884 1902 94912 2071
rect 94872 1896 94924 1902
rect 94872 1838 94924 1844
rect 96632 921 96660 2479
rect 97276 2145 97304 2479
rect 97262 2136 97318 2145
rect 100850 2136 100906 2145
rect 97262 2071 97318 2080
rect 99392 1630 99420 2108
rect 100850 2071 100906 2080
rect 100760 1896 100812 1902
rect 100864 1850 100892 2071
rect 102704 1902 102732 2108
rect 102692 1896 102744 1902
rect 100812 1844 100892 1850
rect 100760 1838 100892 1844
rect 100772 1822 100892 1838
rect 100956 1822 101260 1850
rect 102692 1838 102744 1844
rect 100714 1760 100766 1766
rect 100956 1714 100984 1822
rect 100766 1708 100984 1714
rect 100714 1702 100984 1708
rect 100726 1686 100984 1702
rect 101036 1692 101088 1698
rect 101036 1634 101088 1640
rect 97264 1624 97316 1630
rect 97264 1566 97316 1572
rect 99380 1624 99432 1630
rect 99380 1566 99432 1572
rect 100714 1624 100766 1630
rect 100944 1624 100996 1630
rect 100766 1572 100800 1578
rect 100714 1566 100800 1572
rect 100944 1566 100996 1572
rect 97276 1494 97304 1566
rect 100726 1550 100800 1566
rect 97264 1488 97316 1494
rect 97264 1430 97316 1436
rect 100772 1306 100800 1550
rect 100956 1306 100984 1566
rect 100772 1278 100984 1306
rect 101048 1193 101076 1634
rect 101232 1630 101260 1822
rect 101220 1624 101272 1630
rect 101220 1566 101272 1572
rect 101034 1184 101090 1193
rect 101034 1119 101090 1128
rect 96618 912 96674 921
rect 96618 847 96674 856
rect 98288 882 98408 898
rect 98288 876 98420 882
rect 98288 870 98368 876
rect 92664 808 92716 814
rect 32416 734 32720 762
rect 32770 -400 32826 800
rect 98288 800 98316 870
rect 98368 818 98420 824
rect 92664 750 92716 756
rect 98274 -400 98330 800
rect 103716 746 103744 2615
rect 104164 1896 104216 1902
rect 104164 1838 104216 1844
rect 104176 1698 104204 1838
rect 104164 1692 104216 1698
rect 104164 1634 104216 1640
rect 103992 1550 104296 1578
rect 103992 1329 104020 1550
rect 104268 1494 104296 1550
rect 104164 1488 104216 1494
rect 104164 1430 104216 1436
rect 104256 1488 104308 1494
rect 104256 1430 104308 1436
rect 104176 1329 104204 1430
rect 103978 1320 104034 1329
rect 103978 1255 104034 1264
rect 104162 1320 104218 1329
rect 104162 1255 104218 1264
rect 104360 1193 104388 2615
rect 104346 1184 104402 1193
rect 104346 1119 104402 1128
rect 105096 882 105124 2615
rect 106016 1698 106044 2108
rect 106004 1692 106056 1698
rect 106004 1634 106056 1640
rect 106292 1494 106320 2615
rect 106462 2408 106518 2417
rect 106462 2343 106518 2352
rect 106280 1488 106332 1494
rect 106280 1430 106332 1436
rect 106372 1488 106424 1494
rect 106372 1430 106424 1436
rect 105084 876 105136 882
rect 105084 818 105136 824
rect 106384 746 106412 1430
rect 106476 921 106504 2343
rect 106830 2272 106886 2281
rect 107014 2272 107070 2281
rect 106886 2230 107014 2258
rect 106830 2207 106886 2216
rect 107014 2207 107070 2216
rect 107120 2122 107148 2638
rect 107612 2615 107668 2624
rect 107198 2544 107254 2553
rect 107566 2544 107622 2553
rect 107198 2479 107254 2488
rect 107304 2502 107566 2530
rect 107212 2258 107240 2479
rect 107304 2417 107332 2502
rect 107566 2479 107622 2488
rect 107290 2408 107346 2417
rect 107290 2343 107346 2352
rect 107612 2408 107668 2417
rect 107612 2343 107668 2352
rect 107626 2258 107654 2343
rect 107212 2230 107654 2258
rect 107028 2094 107148 2122
rect 107290 2136 107346 2145
rect 107028 1057 107056 2094
rect 107566 2136 107622 2145
rect 107346 2094 107566 2122
rect 107290 2071 107346 2080
rect 107566 2071 107622 2080
rect 107106 2000 107162 2009
rect 107106 1935 107162 1944
rect 107566 2000 107622 2009
rect 107566 1935 107622 1944
rect 107120 1850 107148 1935
rect 107580 1850 107608 1935
rect 109328 1902 109356 2108
rect 107120 1822 107608 1850
rect 109224 1896 109276 1902
rect 109224 1838 109276 1844
rect 109316 1896 109368 1902
rect 109316 1838 109368 1844
rect 109236 1170 109264 1838
rect 109420 1494 109448 2751
rect 109512 1737 109540 3431
rect 109604 1834 109632 7534
rect 109880 3641 109908 50918
rect 110326 48376 110382 48385
rect 109972 48334 110326 48362
rect 109682 3632 109738 3641
rect 109682 3567 109738 3576
rect 109866 3632 109922 3641
rect 109866 3567 109922 3576
rect 109592 1828 109644 1834
rect 109592 1770 109644 1776
rect 109498 1728 109554 1737
rect 109498 1663 109554 1672
rect 109316 1488 109368 1494
rect 109316 1430 109368 1436
rect 109408 1488 109460 1494
rect 109696 1442 109724 3567
rect 109866 2816 109922 2825
rect 109866 2751 109922 2760
rect 109880 1442 109908 2751
rect 109972 1766 110000 48334
rect 110326 48311 110382 48320
rect 110326 47152 110382 47161
rect 110326 47087 110382 47096
rect 110340 45554 110368 47087
rect 110064 45526 110368 45554
rect 110064 7834 110092 45526
rect 110326 44296 110382 44305
rect 110156 44254 110326 44282
rect 110156 7970 110184 44254
rect 110326 44231 110382 44240
rect 110326 41440 110382 41449
rect 110326 41375 110382 41384
rect 110340 35894 110368 41375
rect 110248 35866 110368 35894
rect 110248 8294 110276 35866
rect 110326 34640 110382 34649
rect 110326 34575 110382 34584
rect 110340 8401 110368 34575
rect 110326 8392 110382 8401
rect 110326 8327 110382 8336
rect 110248 8266 110368 8294
rect 110340 8129 110368 8266
rect 110602 8256 110658 8265
rect 110602 8191 110658 8200
rect 110326 8120 110382 8129
rect 110326 8055 110382 8064
rect 110510 8120 110566 8129
rect 110510 8055 110566 8064
rect 110156 7942 110368 7970
rect 110064 7806 110184 7834
rect 110050 3632 110106 3641
rect 110050 3567 110106 3576
rect 109960 1760 110012 1766
rect 109960 1702 110012 1708
rect 109408 1430 109460 1436
rect 109328 1306 109356 1430
rect 109512 1414 109724 1442
rect 109788 1414 109908 1442
rect 109512 1306 109540 1414
rect 109788 1306 109816 1414
rect 109328 1278 109540 1306
rect 109604 1278 109816 1306
rect 109604 1170 109632 1278
rect 109236 1142 109632 1170
rect 107014 1048 107070 1057
rect 107014 983 107070 992
rect 106462 912 106518 921
rect 106462 847 106518 856
rect 110064 814 110092 3567
rect 110156 1630 110184 7806
rect 110234 3904 110290 3913
rect 110234 3839 110290 3848
rect 110248 3505 110276 3839
rect 110234 3496 110290 3505
rect 110234 3431 110290 3440
rect 110144 1624 110196 1630
rect 110144 1566 110196 1572
rect 110340 1329 110368 7942
rect 110524 5794 110552 8055
rect 110432 5766 110552 5794
rect 110432 1562 110460 5766
rect 110510 5672 110566 5681
rect 110510 5607 110566 5616
rect 110524 2825 110552 5607
rect 110616 3233 110644 8191
rect 111062 7032 111118 7041
rect 111062 6967 111118 6976
rect 110602 3224 110658 3233
rect 110602 3159 110658 3168
rect 110510 2816 110566 2825
rect 110510 2751 110566 2760
rect 111076 1970 111104 6967
rect 111706 2952 111762 2961
rect 111706 2887 111708 2896
rect 111760 2887 111762 2896
rect 111708 2858 111760 2864
rect 111800 2848 111852 2854
rect 111800 2790 111852 2796
rect 111064 1964 111116 1970
rect 111064 1906 111116 1912
rect 110420 1556 110472 1562
rect 110420 1498 110472 1504
rect 110326 1320 110382 1329
rect 110326 1255 110382 1264
rect 111812 1086 111840 2790
rect 112456 1766 112484 62086
rect 112536 42832 112588 42838
rect 112536 42774 112588 42780
rect 112444 1760 112496 1766
rect 112444 1702 112496 1708
rect 111800 1080 111852 1086
rect 111800 1022 111852 1028
rect 112548 950 112576 42774
rect 113836 7721 113864 63514
rect 113928 19009 113956 66234
rect 114020 30433 114048 67594
rect 114112 41857 114140 69022
rect 114204 53145 114232 71742
rect 116306 70272 116362 70281
rect 116306 70207 116362 70216
rect 116320 69086 116348 70207
rect 116308 69080 116360 69086
rect 116308 69022 116360 69028
rect 116122 68368 116178 68377
rect 116122 68303 116178 68312
rect 116136 67658 116164 68303
rect 116124 67652 116176 67658
rect 116124 67594 116176 67600
rect 116582 66464 116638 66473
rect 116582 66399 116638 66408
rect 116596 66298 116624 66399
rect 116584 66292 116636 66298
rect 116584 66234 116636 66240
rect 116688 64874 116716 74015
rect 519266 73672 519322 73681
rect 519266 73607 519322 73616
rect 519280 67833 519308 73607
rect 519924 69193 519952 75103
rect 520016 70553 520044 76599
rect 520108 72457 520136 78095
rect 520200 73273 520228 79591
rect 520292 78577 520320 85711
rect 520384 85377 520412 93327
rect 521382 91896 521438 91905
rect 521382 91831 521438 91840
rect 521198 90264 521254 90273
rect 521198 90199 521254 90208
rect 521106 87272 521162 87281
rect 521106 87207 521162 87216
rect 520370 85368 520426 85377
rect 520370 85303 520426 85312
rect 520922 84280 520978 84289
rect 520922 84215 520978 84224
rect 520278 78568 520334 78577
rect 520278 78503 520334 78512
rect 520936 77217 520964 84215
rect 521120 79937 521148 87207
rect 521212 82657 521240 90199
rect 521290 88768 521346 88777
rect 521290 88703 521346 88712
rect 521198 82648 521254 82657
rect 521198 82583 521254 82592
rect 521304 81297 521332 88703
rect 521396 84017 521424 91831
rect 521566 86728 521622 86737
rect 521672 86714 521700 93826
rect 521622 86686 521700 86714
rect 521566 86663 521622 86672
rect 521382 84008 521438 84017
rect 521382 83943 521438 83952
rect 521290 81288 521346 81297
rect 521290 81223 521346 81232
rect 521106 79928 521162 79937
rect 521106 79863 521162 79872
rect 520922 77208 520978 77217
rect 520922 77143 520978 77152
rect 520186 73264 520242 73273
rect 520186 73199 520242 73208
rect 520094 72448 520150 72457
rect 520094 72383 520150 72392
rect 520186 72040 520242 72049
rect 520186 71975 520242 71984
rect 520002 70544 520058 70553
rect 520002 70479 520058 70488
rect 520094 70408 520150 70417
rect 520094 70343 520150 70352
rect 519910 69184 519966 69193
rect 519910 69119 519966 69128
rect 519634 69048 519690 69057
rect 519634 68983 519690 68992
rect 519266 67824 519322 67833
rect 519266 67759 519322 67768
rect 116596 64846 116716 64874
rect 116596 64734 116624 64846
rect 116584 64728 116636 64734
rect 116584 64670 116636 64676
rect 116214 64560 116270 64569
rect 116214 64495 116270 64504
rect 116228 63578 116256 64495
rect 519648 63753 519676 68983
rect 520108 65113 520136 70343
rect 520200 66473 520228 71975
rect 520462 67552 520518 67561
rect 520462 67487 520518 67496
rect 520186 66464 520242 66473
rect 520186 66399 520242 66408
rect 520370 66056 520426 66065
rect 520370 65991 520426 66000
rect 520094 65104 520150 65113
rect 520094 65039 520150 65048
rect 519634 63744 519690 63753
rect 519634 63679 519690 63688
rect 116216 63572 116268 63578
rect 116216 63514 116268 63520
rect 116122 62656 116178 62665
rect 116122 62591 116178 62600
rect 116136 62150 116164 62591
rect 116124 62144 116176 62150
rect 116124 62086 116176 62092
rect 520278 61432 520334 61441
rect 520278 61367 520334 61376
rect 116582 60616 116638 60625
rect 116582 60551 116638 60560
rect 114190 53136 114246 53145
rect 114190 53071 114246 53080
rect 116122 43344 116178 43353
rect 116122 43279 116178 43288
rect 116136 42838 116164 43279
rect 116124 42832 116176 42838
rect 116124 42774 116176 42780
rect 114098 41848 114154 41857
rect 114098 41783 114154 41792
rect 114006 30424 114062 30433
rect 114006 30359 114062 30368
rect 116490 27976 116546 27985
rect 116490 27911 116546 27920
rect 116306 26072 116362 26081
rect 116306 26007 116362 26016
rect 116214 22264 116270 22273
rect 116214 22199 116270 22208
rect 116030 20360 116086 20369
rect 116030 20295 116086 20304
rect 113914 19000 113970 19009
rect 113914 18935 113970 18944
rect 115938 16416 115994 16425
rect 115938 16351 115994 16360
rect 115848 7948 115900 7954
rect 115848 7890 115900 7896
rect 113822 7712 113878 7721
rect 113822 7647 113878 7656
rect 115860 5681 115888 7890
rect 115846 5672 115902 5681
rect 115846 5607 115902 5616
rect 115952 2281 115980 16351
rect 116044 2553 116072 20295
rect 116122 18456 116178 18465
rect 116122 18391 116178 18400
rect 116030 2544 116086 2553
rect 116030 2479 116086 2488
rect 116136 2417 116164 18391
rect 116228 2689 116256 22199
rect 116320 3641 116348 26007
rect 116398 24168 116454 24177
rect 116398 24103 116454 24112
rect 116306 3632 116362 3641
rect 116306 3567 116362 3576
rect 116306 3088 116362 3097
rect 116306 3023 116362 3032
rect 116214 2680 116270 2689
rect 116214 2615 116270 2624
rect 116122 2408 116178 2417
rect 116122 2343 116178 2352
rect 115938 2272 115994 2281
rect 115938 2207 115994 2216
rect 116320 1358 116348 3023
rect 116308 1352 116360 1358
rect 116308 1294 116360 1300
rect 116412 1290 116440 24103
rect 116504 1426 116532 27911
rect 116596 1698 116624 60551
rect 116674 58712 116730 58721
rect 116674 58647 116730 58656
rect 116688 7834 116716 58647
rect 520186 56944 520242 56953
rect 520292 56930 520320 61367
rect 520384 61033 520412 65991
rect 520476 62393 520504 67487
rect 521106 64560 521162 64569
rect 521106 64495 521162 64504
rect 520462 62384 520518 62393
rect 520462 62319 520518 62328
rect 520370 61024 520426 61033
rect 520370 60959 520426 60968
rect 521014 59936 521070 59945
rect 521014 59871 521070 59880
rect 520242 56902 520320 56930
rect 520370 56944 520426 56953
rect 520186 56879 520242 56888
rect 520370 56879 520426 56888
rect 116766 56808 116822 56817
rect 116766 56743 116822 56752
rect 116780 7954 116808 56743
rect 520278 55448 520334 55457
rect 520278 55383 520334 55392
rect 519266 53816 519322 53825
rect 519266 53751 519322 53760
rect 519280 50153 519308 53751
rect 520094 52320 520150 52329
rect 520094 52255 520150 52264
rect 520002 50824 520058 50833
rect 520002 50759 520058 50768
rect 519266 50144 519322 50153
rect 519266 50079 519322 50088
rect 519450 47832 519506 47841
rect 519450 47767 519506 47776
rect 519464 44713 519492 47767
rect 520016 47433 520044 50759
rect 520108 48793 520136 52255
rect 520292 51513 520320 55383
rect 520384 52873 520412 56879
rect 521028 55593 521056 59871
rect 521120 59673 521148 64495
rect 521198 62928 521254 62937
rect 521198 62863 521254 62872
rect 521106 59664 521162 59673
rect 521106 59599 521162 59608
rect 521106 58440 521162 58449
rect 521106 58375 521162 58384
rect 521014 55584 521070 55593
rect 521014 55519 521070 55528
rect 521120 54233 521148 58375
rect 521212 58313 521240 62863
rect 521198 58304 521254 58313
rect 521198 58239 521254 58248
rect 521106 54224 521162 54233
rect 521106 54159 521162 54168
rect 520370 52864 520426 52873
rect 520370 52799 520426 52808
rect 520278 51504 520334 51513
rect 520278 51439 520334 51448
rect 520186 49328 520242 49337
rect 520186 49263 520242 49272
rect 520094 48784 520150 48793
rect 520094 48719 520150 48728
rect 520002 47424 520058 47433
rect 520002 47359 520058 47368
rect 519910 46336 519966 46345
rect 519910 46271 519966 46280
rect 519450 44704 519506 44713
rect 519450 44639 519506 44648
rect 519818 44704 519874 44713
rect 519818 44639 519874 44648
rect 519832 41993 519860 44639
rect 519924 43353 519952 46271
rect 520200 46073 520228 49263
rect 520186 46064 520242 46073
rect 520186 45999 520242 46008
rect 519910 43344 519966 43353
rect 519910 43279 519966 43288
rect 520186 43208 520242 43217
rect 520186 43143 520242 43152
rect 519818 41984 519874 41993
rect 519818 41919 519874 41928
rect 520094 41712 520150 41721
rect 520094 41647 520150 41656
rect 116950 39536 117006 39545
rect 116950 39471 117006 39480
rect 116858 37632 116914 37641
rect 116858 37567 116914 37576
rect 116768 7948 116820 7954
rect 116768 7890 116820 7896
rect 116688 7806 116808 7834
rect 116676 7744 116728 7750
rect 116676 7686 116728 7692
rect 116584 1692 116636 1698
rect 116584 1634 116636 1640
rect 116492 1420 116544 1426
rect 116492 1362 116544 1368
rect 116400 1284 116452 1290
rect 116400 1226 116452 1232
rect 116688 1222 116716 7686
rect 116780 7041 116808 7806
rect 116766 7032 116822 7041
rect 116766 6967 116822 6976
rect 116676 1216 116728 1222
rect 116676 1158 116728 1164
rect 116872 1018 116900 37567
rect 116964 7818 116992 39471
rect 520108 39273 520136 41647
rect 520200 40633 520228 43143
rect 520186 40624 520242 40633
rect 520186 40559 520242 40568
rect 520186 40216 520242 40225
rect 520186 40151 520242 40160
rect 520094 39264 520150 39273
rect 520094 39199 520150 39208
rect 519818 38720 519874 38729
rect 519818 38655 519874 38664
rect 519832 36553 519860 38655
rect 520200 37913 520228 40151
rect 520186 37904 520242 37913
rect 520186 37839 520242 37848
rect 521566 37224 521622 37233
rect 521566 37159 521622 37168
rect 519818 36544 519874 36553
rect 519818 36479 519874 36488
rect 521580 36009 521608 37159
rect 521566 36000 521622 36009
rect 521566 35935 521622 35944
rect 521106 35592 521162 35601
rect 521106 35527 521162 35536
rect 521120 34513 521148 35527
rect 521106 34504 521162 34513
rect 521106 34439 521162 34448
rect 520922 34096 520978 34105
rect 520922 34031 520978 34040
rect 117134 33824 117190 33833
rect 117134 33759 117190 33768
rect 117042 31784 117098 31793
rect 117042 31719 117098 31728
rect 117056 7818 117084 31719
rect 116952 7812 117004 7818
rect 116952 7754 117004 7760
rect 117044 7812 117096 7818
rect 117044 7754 117096 7760
rect 117148 7698 117176 33759
rect 520936 33153 520964 34031
rect 520922 33144 520978 33153
rect 520922 33079 520978 33088
rect 520922 32600 520978 32609
rect 520922 32535 520978 32544
rect 520936 31657 520964 32535
rect 520922 31648 520978 31657
rect 520922 31583 520978 31592
rect 520922 31104 520978 31113
rect 520922 31039 520978 31048
rect 520936 30297 520964 31039
rect 520922 30288 520978 30297
rect 520922 30223 520978 30232
rect 117226 29880 117282 29889
rect 117226 29815 117282 29824
rect 117240 7886 117268 29815
rect 521106 29608 521162 29617
rect 521106 29543 521162 29552
rect 521120 28393 521148 29543
rect 521106 28384 521162 28393
rect 521106 28319 521162 28328
rect 521106 21992 521162 22001
rect 521106 21927 521162 21936
rect 521120 20913 521148 21927
rect 521106 20904 521162 20913
rect 521106 20839 521162 20848
rect 520738 20496 520794 20505
rect 520738 20431 520794 20440
rect 520752 19553 520780 20431
rect 520738 19544 520794 19553
rect 520738 19479 520794 19488
rect 520922 19000 520978 19009
rect 520922 18935 520978 18944
rect 520936 18193 520964 18935
rect 520922 18184 520978 18193
rect 520922 18119 520978 18128
rect 521106 9344 521162 9353
rect 521106 9279 521162 9288
rect 521120 8265 521148 9279
rect 521106 8256 521162 8265
rect 521106 8191 521162 8200
rect 520370 7984 520426 7993
rect 520370 7919 520426 7928
rect 117228 7880 117280 7886
rect 117228 7822 117280 7828
rect 117320 7812 117372 7818
rect 117320 7754 117372 7760
rect 116964 7670 117176 7698
rect 116964 3369 116992 7670
rect 117332 7562 117360 7754
rect 117240 7534 117360 7562
rect 117044 7472 117096 7478
rect 117044 7414 117096 7420
rect 116950 3360 117006 3369
rect 116950 3295 117006 3304
rect 117056 3233 117084 7414
rect 117134 6896 117190 6905
rect 117134 6831 117190 6840
rect 117042 3224 117098 3233
rect 117042 3159 117098 3168
rect 117148 1465 117176 6831
rect 117134 1456 117190 1465
rect 117134 1391 117190 1400
rect 117240 1154 117268 7534
rect 520384 6769 520412 7919
rect 520370 6760 520426 6769
rect 520370 6695 520426 6704
rect 521106 6624 521162 6633
rect 521106 6559 521162 6568
rect 521120 5273 521148 6559
rect 520922 5264 520978 5273
rect 520922 5199 520978 5208
rect 521106 5264 521162 5273
rect 521106 5199 521162 5208
rect 520936 3777 520964 5199
rect 521014 3904 521070 3913
rect 521014 3839 521070 3848
rect 520922 3768 520978 3777
rect 520922 3703 520978 3712
rect 193600 2514 193936 2530
rect 443656 2514 443992 2530
rect 170312 2508 170364 2514
rect 170312 2450 170364 2456
rect 193588 2508 193936 2514
rect 193640 2502 193936 2508
rect 294788 2508 294840 2514
rect 193588 2450 193640 2456
rect 294788 2450 294840 2456
rect 425796 2508 425848 2514
rect 425796 2450 425848 2456
rect 443644 2508 443992 2514
rect 443696 2502 443992 2508
rect 443644 2450 443696 2456
rect 170324 2378 170352 2450
rect 170312 2372 170364 2378
rect 170312 2314 170364 2320
rect 143644 2094 143980 2122
rect 243648 2094 243984 2122
rect 293604 2094 293940 2122
rect 143644 1494 143672 2094
rect 229282 1592 229338 1601
rect 229282 1527 229338 1536
rect 143632 1488 143684 1494
rect 143632 1430 143684 1436
rect 163778 1456 163834 1465
rect 163778 1391 163834 1400
rect 117228 1148 117280 1154
rect 117228 1090 117280 1096
rect 116860 1012 116912 1018
rect 116860 954 116912 960
rect 112536 944 112588 950
rect 112536 886 112588 892
rect 110052 808 110104 814
rect 163792 800 163820 1391
rect 229296 800 229324 1527
rect 243648 1465 243676 2094
rect 293604 1601 293632 2094
rect 293590 1592 293646 1601
rect 293590 1527 293646 1536
rect 243634 1456 243690 1465
rect 294800 1426 294828 2450
rect 343652 2094 343988 2122
rect 393608 2094 393944 2122
rect 343652 1426 343680 2094
rect 393608 1465 393636 2094
rect 360290 1456 360346 1465
rect 243634 1391 243690 1400
rect 294788 1420 294840 1426
rect 294788 1362 294840 1368
rect 343640 1420 343692 1426
rect 360290 1391 360346 1400
rect 393594 1456 393650 1465
rect 393594 1391 393650 1400
rect 343640 1362 343692 1368
rect 294800 800 294828 1362
rect 360304 800 360332 1391
rect 425808 800 425836 2450
rect 521028 2281 521056 3839
rect 521106 2680 521162 2689
rect 521106 2615 521162 2624
rect 521014 2272 521070 2281
rect 521014 2207 521070 2216
rect 493612 2094 493948 2122
rect 493612 1426 493640 2094
rect 491300 1420 491352 1426
rect 491300 1362 491352 1368
rect 493600 1420 493652 1426
rect 493600 1362 493652 1368
rect 491312 800 491340 1362
rect 110052 750 110104 756
rect 103704 740 103756 746
rect 103704 682 103756 688
rect 106372 740 106424 746
rect 106372 682 106424 688
rect 163778 -400 163834 800
rect 229282 -400 229338 800
rect 294786 -400 294842 800
rect 360290 -400 360346 800
rect 425794 -400 425850 800
rect 491298 -400 491354 800
rect 521120 785 521148 2615
rect 521106 776 521162 785
rect 521106 711 521162 720
<< via2 >>
rect 9586 159432 9642 159488
rect 9678 153992 9734 154048
rect 7562 153856 7618 153912
rect 7102 153720 7158 153776
rect 5538 152360 5594 152416
rect 6090 150592 6146 150648
rect 2686 150456 2742 150512
rect 16302 159296 16358 159352
rect 19706 154128 19762 154184
rect 19338 152496 19394 152552
rect 29734 159568 29790 159624
rect 24858 152632 24914 152688
rect 33966 157936 34022 157992
rect 35622 156576 35678 156632
rect 40682 158072 40738 158128
rect 42338 156712 42394 156768
rect 43994 158208 44050 158264
rect 52366 156848 52422 156904
rect 55770 156984 55826 157040
rect 57426 158344 57482 158400
rect 58254 155352 58310 155408
rect 61658 155216 61714 155272
rect 37370 154264 37426 154320
rect 68374 155488 68430 155544
rect 65154 154400 65210 154456
rect 85118 155624 85174 155680
rect 101126 158480 101182 158536
rect 104438 157120 104494 157176
rect 99930 149776 99986 149832
rect 92570 149640 92626 149696
rect 109590 148008 109646 148064
rect 118698 153040 118754 153096
rect 111062 150456 111118 150512
rect 110970 147328 111026 147384
rect 110326 146376 110382 146432
rect 111338 150592 111394 150648
rect 111706 147328 111762 147384
rect 113822 144200 113878 144256
rect 116122 145152 116178 145208
rect 116030 143248 116086 143304
rect 115294 141344 115350 141400
rect 116122 139440 116178 139496
rect 116122 137536 116178 137592
rect 115202 135496 115258 135552
rect 116030 133592 116086 133648
rect 114190 132776 114246 132832
rect 113914 121352 113970 121408
rect 114006 110064 114062 110120
rect 114098 98640 114154 98696
rect 114190 87216 114246 87272
rect 116122 131688 116178 131744
rect 116582 149640 116638 149696
rect 116398 129784 116454 129840
rect 116306 127880 116362 127936
rect 116030 125976 116086 126032
rect 116122 124108 116124 124128
rect 116124 124108 116176 124128
rect 116176 124108 116178 124128
rect 116122 124072 116178 124108
rect 115938 122168 115994 122224
rect 116122 120128 116178 120184
rect 116122 118224 116178 118280
rect 116122 116320 116178 116376
rect 116122 114452 116124 114472
rect 116124 114452 116176 114472
rect 116176 114452 116178 114472
rect 116122 114416 116178 114452
rect 115938 112512 115994 112568
rect 116122 110608 116178 110664
rect 116122 108704 116178 108760
rect 116490 106800 116546 106856
rect 116858 149776 116914 149832
rect 116950 102856 117006 102912
rect 121090 153040 121146 153096
rect 122562 158908 122618 158944
rect 122562 158888 122564 158908
rect 122564 158888 122616 158908
rect 122616 158888 122618 158908
rect 123850 159432 123906 159488
rect 124494 158888 124550 158944
rect 124954 153856 125010 153912
rect 124310 153720 124366 153776
rect 124494 153720 124550 153776
rect 123850 153040 123906 153096
rect 123666 152360 123722 152416
rect 126886 153992 126942 154048
rect 126242 153040 126298 153096
rect 127346 153992 127402 154048
rect 129554 154028 129556 154048
rect 129556 154028 129608 154048
rect 129608 154028 129610 154048
rect 129554 153992 129610 154028
rect 131302 159296 131358 159352
rect 133602 159704 133658 159760
rect 134614 154128 134670 154184
rect 132866 153040 132922 153096
rect 133970 152496 134026 152552
rect 137374 159724 137430 159760
rect 137374 159704 137376 159724
rect 137376 159704 137428 159724
rect 137428 159704 137430 159724
rect 138478 152632 138534 152688
rect 139398 159568 139454 159624
rect 141054 153040 141110 153096
rect 145010 157936 145066 157992
rect 145102 156576 145158 156632
rect 146850 154148 146906 154184
rect 146850 154128 146852 154148
rect 146852 154128 146904 154148
rect 146904 154128 146906 154148
rect 148138 154264 148194 154320
rect 149610 158072 149666 158128
rect 152370 158208 152426 158264
rect 153014 158244 153016 158264
rect 153016 158244 153068 158264
rect 153068 158244 153070 158264
rect 153014 158208 153070 158244
rect 151266 156712 151322 156768
rect 151726 155080 151782 155136
rect 152738 155080 152794 155136
rect 153014 154128 153070 154184
rect 155222 158208 155278 158264
rect 158994 156848 159050 156904
rect 161570 156984 161626 157040
rect 162950 158344 163006 158400
rect 163410 155352 163466 155408
rect 166078 155216 166134 155272
rect 165710 154264 165766 154320
rect 166354 154264 166410 154320
rect 169298 154400 169354 154456
rect 171230 155488 171286 155544
rect 184018 155624 184074 155680
rect 187882 156460 187938 156496
rect 187882 156440 187884 156460
rect 187884 156440 187936 156460
rect 187936 156440 187938 156460
rect 189446 153312 189502 153368
rect 189722 153584 189778 153640
rect 191194 156440 191250 156496
rect 191286 153604 191342 153640
rect 191286 153584 191288 153604
rect 191288 153584 191340 153604
rect 191340 153584 191342 153604
rect 191286 153312 191342 153368
rect 196254 158480 196310 158536
rect 198830 157120 198886 157176
rect 200118 153720 200174 153776
rect 217138 152360 217194 152416
rect 221278 153720 221334 153776
rect 274546 153332 274602 153368
rect 274546 153312 274548 153332
rect 274548 153312 274600 153332
rect 274600 153312 274602 153332
rect 275926 153332 275982 153368
rect 275926 153312 275928 153332
rect 275928 153312 275980 153332
rect 275980 153312 275982 153332
rect 285494 152360 285550 152416
rect 288346 159296 288402 159352
rect 288714 153720 288770 153776
rect 310702 152360 310758 152416
rect 339406 159296 339462 159352
rect 348790 159332 348792 159352
rect 348792 159332 348844 159352
rect 348844 159332 348846 159352
rect 348790 159296 348846 159332
rect 349894 159296 349950 159352
rect 356150 152360 356206 152416
rect 432878 152360 432934 152416
rect 445666 151852 445668 151872
rect 445668 151852 445720 151872
rect 445720 151852 445722 151872
rect 445666 151816 445722 151852
rect 446586 151972 446642 152008
rect 446586 151952 446588 151972
rect 446588 151952 446640 151972
rect 446640 151952 446642 151972
rect 446954 152668 446956 152688
rect 446956 152668 447008 152688
rect 447008 152668 447010 152688
rect 446954 152632 447010 152668
rect 447414 152652 447470 152688
rect 447414 152632 447416 152652
rect 447416 152632 447468 152652
rect 447468 152632 447470 152652
rect 447046 151816 447102 151872
rect 449898 152360 449954 152416
rect 448058 151972 448114 152008
rect 448058 151952 448060 151972
rect 448060 151952 448112 151972
rect 448112 151952 448114 151972
rect 519726 163104 519782 163160
rect 519542 161608 519598 161664
rect 519450 153992 519506 154048
rect 519174 141888 519230 141944
rect 519634 160112 519690 160168
rect 519542 147872 519598 147928
rect 520002 158616 520058 158672
rect 519910 157120 519966 157176
rect 519818 155624 519874 155680
rect 519726 149232 519782 149288
rect 519726 148008 519782 148064
rect 519634 146512 519690 146568
rect 519542 144880 519598 144936
rect 519450 141072 519506 141128
rect 519266 140392 519322 140448
rect 519174 130192 519230 130248
rect 519358 138896 519414 138952
rect 519266 128832 519322 128888
rect 519174 128288 519230 128344
rect 519450 137400 519506 137456
rect 519358 127472 519414 127528
rect 519266 126656 519322 126712
rect 519174 117952 519230 118008
rect 521014 152496 521070 152552
rect 520186 151000 520242 151056
rect 520094 149504 520150 149560
rect 520002 145152 520058 145208
rect 519910 143792 519966 143848
rect 520002 143384 520058 143440
rect 519818 142432 519874 142488
rect 519910 135768 519966 135824
rect 519726 135632 519782 135688
rect 519818 134272 519874 134328
rect 519542 132912 519598 132968
rect 519726 132776 519782 132832
rect 519634 131280 519690 131336
rect 519542 129784 519598 129840
rect 519450 126112 519506 126168
rect 520922 146512 520978 146568
rect 520186 138352 520242 138408
rect 520094 136992 520150 137048
rect 521014 139712 521070 139768
rect 520922 134408 520978 134464
rect 520002 131552 520058 131608
rect 520186 125160 520242 125216
rect 519910 124752 519966 124808
rect 520094 123664 520150 123720
rect 519818 123392 519874 123448
rect 519910 122168 519966 122224
rect 519726 122032 519782 122088
rect 519634 120672 519690 120728
rect 519818 120672 519874 120728
rect 519542 119312 519598 119368
rect 519726 119176 519782 119232
rect 519266 116592 519322 116648
rect 519634 116048 519690 116104
rect 519542 114552 519598 114608
rect 520002 117544 520058 117600
rect 519910 112512 519966 112568
rect 519818 111152 519874 111208
rect 519726 109792 519782 109848
rect 520186 115232 520242 115288
rect 520094 113872 520150 113928
rect 520922 113056 520978 113112
rect 520002 108432 520058 108488
rect 519634 107072 519690 107128
rect 519542 105712 519598 105768
rect 520278 105440 520334 105496
rect 117134 104760 117190 104816
rect 117042 100952 117098 101008
rect 519818 99320 519874 99376
rect 116858 99048 116914 99104
rect 519726 97824 519782 97880
rect 116766 97144 116822 97200
rect 116674 95240 116730 95296
rect 116582 93336 116638 93392
rect 116122 91296 116178 91352
rect 521290 111560 521346 111616
rect 521198 106936 521254 106992
rect 520922 104352 520978 104408
rect 521106 103944 521162 104000
rect 521014 102448 521070 102504
rect 520278 97552 520334 97608
rect 520002 96328 520058 96384
rect 519910 94832 519966 94888
rect 519818 92112 519874 92168
rect 519726 90752 519782 90808
rect 116122 89392 116178 89448
rect 521474 110064 521530 110120
rect 521382 108432 521438 108488
rect 521290 102992 521346 103048
rect 521290 100952 521346 101008
rect 521198 98912 521254 98968
rect 521106 96192 521162 96248
rect 521014 94968 521070 95024
rect 521474 101632 521530 101688
rect 521382 100272 521438 100328
rect 521290 93472 521346 93528
rect 520370 93336 520426 93392
rect 520002 89392 520058 89448
rect 519910 88032 519966 88088
rect 116030 87488 116086 87544
rect 520278 85720 520334 85776
rect 115202 85584 115258 85640
rect 116582 83680 116638 83736
rect 519910 82728 519966 82784
rect 116214 81776 116270 81832
rect 519634 81096 519690 81152
rect 115938 79872 115994 79928
rect 116122 77968 116178 78024
rect 520186 79600 520242 79656
rect 520094 78104 520150 78160
rect 520002 76608 520058 76664
rect 519910 75928 519966 75984
rect 519910 75112 519966 75168
rect 519634 74568 519690 74624
rect 116674 74024 116730 74080
rect 116582 72120 116638 72176
rect 113362 64504 113418 64560
rect 110326 53896 110382 53952
rect 110326 52536 110382 52592
rect 110326 51040 110382 51096
rect 109498 3576 109554 3632
rect 109498 3440 109554 3496
rect 109406 2760 109462 2816
rect 32402 2624 32458 2680
rect 36358 2624 36414 2680
rect 62394 2624 62450 2680
rect 64142 2624 64198 2680
rect 65338 2624 65394 2680
rect 68006 2624 68062 2680
rect 68558 2624 68614 2680
rect 68834 2624 68890 2680
rect 69386 2624 69442 2680
rect 77022 2624 77078 2680
rect 29550 2352 29606 2408
rect 26054 2216 26110 2272
rect 5998 1672 6054 1728
rect 22926 2080 22982 2136
rect 19614 1944 19670 2000
rect 15934 1808 15990 1864
rect 12622 1536 12678 1592
rect 9310 1400 9366 1456
rect 33046 2488 33102 2544
rect 77252 2624 77308 2680
rect 77758 2624 77814 2680
rect 77942 2624 77998 2680
rect 78126 2624 78182 2680
rect 78310 2624 78366 2680
rect 95698 2624 95754 2680
rect 96342 2624 96398 2680
rect 103702 2624 103758 2680
rect 104346 2624 104402 2680
rect 105082 2624 105138 2680
rect 106278 2624 106334 2680
rect 96618 2488 96674 2544
rect 97262 2488 97318 2544
rect 85946 1264 86002 1320
rect 88338 1128 88394 1184
rect 94870 2080 94926 2136
rect 95698 2080 95754 2136
rect 97262 2080 97318 2136
rect 100850 2080 100906 2136
rect 101034 1128 101090 1184
rect 96618 856 96674 912
rect 103978 1264 104034 1320
rect 104162 1264 104218 1320
rect 104346 1128 104402 1184
rect 106462 2352 106518 2408
rect 106830 2216 106886 2272
rect 107014 2216 107070 2272
rect 107612 2624 107668 2680
rect 107198 2488 107254 2544
rect 107566 2488 107622 2544
rect 107290 2352 107346 2408
rect 107612 2352 107668 2408
rect 107290 2080 107346 2136
rect 107566 2080 107622 2136
rect 107106 1944 107162 2000
rect 107566 1944 107622 2000
rect 109682 3576 109738 3632
rect 109866 3576 109922 3632
rect 109498 1672 109554 1728
rect 109866 2760 109922 2816
rect 110326 48320 110382 48376
rect 110326 47096 110382 47152
rect 110326 44240 110382 44296
rect 110326 41384 110382 41440
rect 110326 34584 110382 34640
rect 110326 8336 110382 8392
rect 110602 8200 110658 8256
rect 110326 8064 110382 8120
rect 110510 8064 110566 8120
rect 110050 3576 110106 3632
rect 107014 992 107070 1048
rect 106462 856 106518 912
rect 110234 3848 110290 3904
rect 110234 3440 110290 3496
rect 110510 5616 110566 5672
rect 111062 6976 111118 7032
rect 110602 3168 110658 3224
rect 110510 2760 110566 2816
rect 111706 2916 111762 2952
rect 111706 2896 111708 2916
rect 111708 2896 111760 2916
rect 111760 2896 111762 2916
rect 110326 1264 110382 1320
rect 116306 70216 116362 70272
rect 116122 68312 116178 68368
rect 116582 66408 116638 66464
rect 519266 73616 519322 73672
rect 521382 91840 521438 91896
rect 521198 90208 521254 90264
rect 521106 87216 521162 87272
rect 520370 85312 520426 85368
rect 520922 84224 520978 84280
rect 520278 78512 520334 78568
rect 521290 88712 521346 88768
rect 521198 82592 521254 82648
rect 521566 86672 521622 86728
rect 521382 83952 521438 84008
rect 521290 81232 521346 81288
rect 521106 79872 521162 79928
rect 520922 77152 520978 77208
rect 520186 73208 520242 73264
rect 520094 72392 520150 72448
rect 520186 71984 520242 72040
rect 520002 70488 520058 70544
rect 520094 70352 520150 70408
rect 519910 69128 519966 69184
rect 519634 68992 519690 69048
rect 519266 67768 519322 67824
rect 116214 64504 116270 64560
rect 520462 67496 520518 67552
rect 520186 66408 520242 66464
rect 520370 66000 520426 66056
rect 520094 65048 520150 65104
rect 519634 63688 519690 63744
rect 116122 62600 116178 62656
rect 520278 61376 520334 61432
rect 116582 60560 116638 60616
rect 114190 53080 114246 53136
rect 116122 43288 116178 43344
rect 114098 41792 114154 41848
rect 114006 30368 114062 30424
rect 116490 27920 116546 27976
rect 116306 26016 116362 26072
rect 116214 22208 116270 22264
rect 116030 20304 116086 20360
rect 113914 18944 113970 19000
rect 115938 16360 115994 16416
rect 113822 7656 113878 7712
rect 115846 5616 115902 5672
rect 116122 18400 116178 18456
rect 116030 2488 116086 2544
rect 116398 24112 116454 24168
rect 116306 3576 116362 3632
rect 116306 3032 116362 3088
rect 116214 2624 116270 2680
rect 116122 2352 116178 2408
rect 115938 2216 115994 2272
rect 116674 58656 116730 58712
rect 520186 56888 520242 56944
rect 521106 64504 521162 64560
rect 520462 62328 520518 62384
rect 520370 60968 520426 61024
rect 521014 59880 521070 59936
rect 520370 56888 520426 56944
rect 116766 56752 116822 56808
rect 520278 55392 520334 55448
rect 519266 53760 519322 53816
rect 520094 52264 520150 52320
rect 520002 50768 520058 50824
rect 519266 50088 519322 50144
rect 519450 47776 519506 47832
rect 521198 62872 521254 62928
rect 521106 59608 521162 59664
rect 521106 58384 521162 58440
rect 521014 55528 521070 55584
rect 521198 58248 521254 58304
rect 521106 54168 521162 54224
rect 520370 52808 520426 52864
rect 520278 51448 520334 51504
rect 520186 49272 520242 49328
rect 520094 48728 520150 48784
rect 520002 47368 520058 47424
rect 519910 46280 519966 46336
rect 519450 44648 519506 44704
rect 519818 44648 519874 44704
rect 520186 46008 520242 46064
rect 519910 43288 519966 43344
rect 520186 43152 520242 43208
rect 519818 41928 519874 41984
rect 520094 41656 520150 41712
rect 116950 39480 117006 39536
rect 116858 37576 116914 37632
rect 116766 6976 116822 7032
rect 520186 40568 520242 40624
rect 520186 40160 520242 40216
rect 520094 39208 520150 39264
rect 519818 38664 519874 38720
rect 520186 37848 520242 37904
rect 521566 37168 521622 37224
rect 519818 36488 519874 36544
rect 521566 35944 521622 36000
rect 521106 35536 521162 35592
rect 521106 34448 521162 34504
rect 520922 34040 520978 34096
rect 117134 33768 117190 33824
rect 117042 31728 117098 31784
rect 520922 33088 520978 33144
rect 520922 32544 520978 32600
rect 520922 31592 520978 31648
rect 520922 31048 520978 31104
rect 520922 30232 520978 30288
rect 117226 29824 117282 29880
rect 521106 29552 521162 29608
rect 521106 28328 521162 28384
rect 521106 21936 521162 21992
rect 521106 20848 521162 20904
rect 520738 20440 520794 20496
rect 520738 19488 520794 19544
rect 520922 18944 520978 19000
rect 520922 18128 520978 18184
rect 521106 9288 521162 9344
rect 521106 8200 521162 8256
rect 520370 7928 520426 7984
rect 116950 3304 117006 3360
rect 117134 6840 117190 6896
rect 117042 3168 117098 3224
rect 117134 1400 117190 1456
rect 520370 6704 520426 6760
rect 521106 6568 521162 6624
rect 520922 5208 520978 5264
rect 521106 5208 521162 5264
rect 521014 3848 521070 3904
rect 520922 3712 520978 3768
rect 229282 1536 229338 1592
rect 163778 1400 163834 1456
rect 293590 1536 293646 1592
rect 243634 1400 243690 1456
rect 360290 1400 360346 1456
rect 393594 1400 393650 1456
rect 521106 2624 521162 2680
rect 521014 2216 521070 2272
rect 521106 720 521162 776
<< metal3 >>
rect 519721 163162 519787 163165
rect 523200 163162 524400 163192
rect 519721 163160 524400 163162
rect 519721 163104 519726 163160
rect 519782 163104 524400 163160
rect 519721 163102 524400 163104
rect 519721 163099 519787 163102
rect 523200 163072 524400 163102
rect 519537 161666 519603 161669
rect 523200 161666 524400 161696
rect 519537 161664 524400 161666
rect 519537 161608 519542 161664
rect 519598 161608 524400 161664
rect 519537 161606 524400 161608
rect 519537 161603 519603 161606
rect 523200 161576 524400 161606
rect 519629 160170 519695 160173
rect 523200 160170 524400 160200
rect 519629 160168 524400 160170
rect 519629 160112 519634 160168
rect 519690 160112 524400 160168
rect 519629 160110 524400 160112
rect 519629 160107 519695 160110
rect 523200 160080 524400 160110
rect 133597 159762 133663 159765
rect 137369 159762 137435 159765
rect 133597 159760 137435 159762
rect 133597 159704 133602 159760
rect 133658 159704 137374 159760
rect 137430 159704 137435 159760
rect 133597 159702 137435 159704
rect 133597 159699 133663 159702
rect 137369 159699 137435 159702
rect 29729 159626 29795 159629
rect 139393 159626 139459 159629
rect 29729 159624 139459 159626
rect 29729 159568 29734 159624
rect 29790 159568 139398 159624
rect 139454 159568 139459 159624
rect 29729 159566 139459 159568
rect 29729 159563 29795 159566
rect 139393 159563 139459 159566
rect 9581 159490 9647 159493
rect 123845 159490 123911 159493
rect 9581 159488 123911 159490
rect 9581 159432 9586 159488
rect 9642 159432 123850 159488
rect 123906 159432 123911 159488
rect 9581 159430 123911 159432
rect 9581 159427 9647 159430
rect 123845 159427 123911 159430
rect 16297 159354 16363 159357
rect 131297 159354 131363 159357
rect 16297 159352 131363 159354
rect 16297 159296 16302 159352
rect 16358 159296 131302 159352
rect 131358 159296 131363 159352
rect 16297 159294 131363 159296
rect 16297 159291 16363 159294
rect 131297 159291 131363 159294
rect 288341 159354 288407 159357
rect 339401 159354 339467 159357
rect 288341 159352 339467 159354
rect 288341 159296 288346 159352
rect 288402 159296 339406 159352
rect 339462 159296 339467 159352
rect 288341 159294 339467 159296
rect 288341 159291 288407 159294
rect 339401 159291 339467 159294
rect 348785 159354 348851 159357
rect 349889 159354 349955 159357
rect 348785 159352 349955 159354
rect 348785 159296 348790 159352
rect 348846 159296 349894 159352
rect 349950 159296 349955 159352
rect 348785 159294 349955 159296
rect 348785 159291 348851 159294
rect 349889 159291 349955 159294
rect 122557 158946 122623 158949
rect 124489 158946 124555 158949
rect 122557 158944 124555 158946
rect 122557 158888 122562 158944
rect 122618 158888 124494 158944
rect 124550 158888 124555 158944
rect 122557 158886 124555 158888
rect 122557 158883 122623 158886
rect 124489 158883 124555 158886
rect 519997 158674 520063 158677
rect 523200 158674 524400 158704
rect 519997 158672 524400 158674
rect 519997 158616 520002 158672
rect 520058 158616 524400 158672
rect 519997 158614 524400 158616
rect 519997 158611 520063 158614
rect 523200 158584 524400 158614
rect 101121 158538 101187 158541
rect 196249 158538 196315 158541
rect 101121 158536 196315 158538
rect 101121 158480 101126 158536
rect 101182 158480 196254 158536
rect 196310 158480 196315 158536
rect 101121 158478 196315 158480
rect 101121 158475 101187 158478
rect 196249 158475 196315 158478
rect 57421 158402 57487 158405
rect 162945 158402 163011 158405
rect 57421 158400 163011 158402
rect 57421 158344 57426 158400
rect 57482 158344 162950 158400
rect 163006 158344 163011 158400
rect 57421 158342 163011 158344
rect 57421 158339 57487 158342
rect 162945 158339 163011 158342
rect 43989 158266 44055 158269
rect 152365 158266 152431 158269
rect 43989 158264 152431 158266
rect 43989 158208 43994 158264
rect 44050 158208 152370 158264
rect 152426 158208 152431 158264
rect 43989 158206 152431 158208
rect 43989 158203 44055 158206
rect 152365 158203 152431 158206
rect 153009 158266 153075 158269
rect 155217 158266 155283 158269
rect 153009 158264 155283 158266
rect 153009 158208 153014 158264
rect 153070 158208 155222 158264
rect 155278 158208 155283 158264
rect 153009 158206 155283 158208
rect 153009 158203 153075 158206
rect 155217 158203 155283 158206
rect 40677 158130 40743 158133
rect 149605 158130 149671 158133
rect 40677 158128 149671 158130
rect 40677 158072 40682 158128
rect 40738 158072 149610 158128
rect 149666 158072 149671 158128
rect 40677 158070 149671 158072
rect 40677 158067 40743 158070
rect 149605 158067 149671 158070
rect 33961 157994 34027 157997
rect 145005 157994 145071 157997
rect 33961 157992 145071 157994
rect 33961 157936 33966 157992
rect 34022 157936 145010 157992
rect 145066 157936 145071 157992
rect 33961 157934 145071 157936
rect 33961 157931 34027 157934
rect 145005 157931 145071 157934
rect 104433 157178 104499 157181
rect 198825 157178 198891 157181
rect 104433 157176 198891 157178
rect 104433 157120 104438 157176
rect 104494 157120 198830 157176
rect 198886 157120 198891 157176
rect 104433 157118 198891 157120
rect 104433 157115 104499 157118
rect 198825 157115 198891 157118
rect 519905 157178 519971 157181
rect 523200 157178 524400 157208
rect 519905 157176 524400 157178
rect 519905 157120 519910 157176
rect 519966 157120 524400 157176
rect 519905 157118 524400 157120
rect 519905 157115 519971 157118
rect 523200 157088 524400 157118
rect 55765 157042 55831 157045
rect 161565 157042 161631 157045
rect 55765 157040 161631 157042
rect 55765 156984 55770 157040
rect 55826 156984 161570 157040
rect 161626 156984 161631 157040
rect 55765 156982 161631 156984
rect 55765 156979 55831 156982
rect 161565 156979 161631 156982
rect 52361 156906 52427 156909
rect 158989 156906 159055 156909
rect 52361 156904 159055 156906
rect 52361 156848 52366 156904
rect 52422 156848 158994 156904
rect 159050 156848 159055 156904
rect 52361 156846 159055 156848
rect 52361 156843 52427 156846
rect 158989 156843 159055 156846
rect 42333 156770 42399 156773
rect 151261 156770 151327 156773
rect 42333 156768 151327 156770
rect 42333 156712 42338 156768
rect 42394 156712 151266 156768
rect 151322 156712 151327 156768
rect 42333 156710 151327 156712
rect 42333 156707 42399 156710
rect 151261 156707 151327 156710
rect 35617 156634 35683 156637
rect 145097 156634 145163 156637
rect 35617 156632 145163 156634
rect 35617 156576 35622 156632
rect 35678 156576 145102 156632
rect 145158 156576 145163 156632
rect 35617 156574 145163 156576
rect 35617 156571 35683 156574
rect 145097 156571 145163 156574
rect 187877 156498 187943 156501
rect 191189 156498 191255 156501
rect 187877 156496 191255 156498
rect 187877 156440 187882 156496
rect 187938 156440 191194 156496
rect 191250 156440 191255 156496
rect 187877 156438 191255 156440
rect 187877 156435 187943 156438
rect 191189 156435 191255 156438
rect 85113 155682 85179 155685
rect 184013 155682 184079 155685
rect 85113 155680 184079 155682
rect 85113 155624 85118 155680
rect 85174 155624 184018 155680
rect 184074 155624 184079 155680
rect 85113 155622 184079 155624
rect 85113 155619 85179 155622
rect 184013 155619 184079 155622
rect 519813 155682 519879 155685
rect 523200 155682 524400 155712
rect 519813 155680 524400 155682
rect 519813 155624 519818 155680
rect 519874 155624 524400 155680
rect 519813 155622 524400 155624
rect 519813 155619 519879 155622
rect 523200 155592 524400 155622
rect 68369 155546 68435 155549
rect 171225 155546 171291 155549
rect 68369 155544 171291 155546
rect 68369 155488 68374 155544
rect 68430 155488 171230 155544
rect 171286 155488 171291 155544
rect 68369 155486 171291 155488
rect 68369 155483 68435 155486
rect 171225 155483 171291 155486
rect 58249 155410 58315 155413
rect 163405 155410 163471 155413
rect 58249 155408 163471 155410
rect 58249 155352 58254 155408
rect 58310 155352 163410 155408
rect 163466 155352 163471 155408
rect 58249 155350 163471 155352
rect 58249 155347 58315 155350
rect 163405 155347 163471 155350
rect 61653 155274 61719 155277
rect 166073 155274 166139 155277
rect 61653 155272 166139 155274
rect 61653 155216 61658 155272
rect 61714 155216 166078 155272
rect 166134 155216 166139 155272
rect 61653 155214 166139 155216
rect 61653 155211 61719 155214
rect 166073 155211 166139 155214
rect 151721 155138 151787 155141
rect 152733 155138 152799 155141
rect 151721 155136 152799 155138
rect 151721 155080 151726 155136
rect 151782 155080 152738 155136
rect 152794 155080 152799 155136
rect 151721 155078 152799 155080
rect 151721 155075 151787 155078
rect 152733 155075 152799 155078
rect 65149 154458 65215 154461
rect 169293 154458 169359 154461
rect 65149 154456 169359 154458
rect 65149 154400 65154 154456
rect 65210 154400 169298 154456
rect 169354 154400 169359 154456
rect 65149 154398 169359 154400
rect 65149 154395 65215 154398
rect 169293 154395 169359 154398
rect 37365 154322 37431 154325
rect 148133 154322 148199 154325
rect 37365 154320 148199 154322
rect 37365 154264 37370 154320
rect 37426 154264 148138 154320
rect 148194 154264 148199 154320
rect 37365 154262 148199 154264
rect 37365 154259 37431 154262
rect 148133 154259 148199 154262
rect 165705 154322 165771 154325
rect 166349 154322 166415 154325
rect 165705 154320 166415 154322
rect 165705 154264 165710 154320
rect 165766 154264 166354 154320
rect 166410 154264 166415 154320
rect 165705 154262 166415 154264
rect 165705 154259 165771 154262
rect 166349 154259 166415 154262
rect 19701 154186 19767 154189
rect 134609 154186 134675 154189
rect 19701 154184 134675 154186
rect 19701 154128 19706 154184
rect 19762 154128 134614 154184
rect 134670 154128 134675 154184
rect 19701 154126 134675 154128
rect 19701 154123 19767 154126
rect 134609 154123 134675 154126
rect 146845 154186 146911 154189
rect 153009 154186 153075 154189
rect 146845 154184 153075 154186
rect 146845 154128 146850 154184
rect 146906 154128 153014 154184
rect 153070 154128 153075 154184
rect 146845 154126 153075 154128
rect 146845 154123 146911 154126
rect 153009 154123 153075 154126
rect 9673 154050 9739 154053
rect 126881 154050 126947 154053
rect 9673 154048 126947 154050
rect 9673 153992 9678 154048
rect 9734 153992 126886 154048
rect 126942 153992 126947 154048
rect 9673 153990 126947 153992
rect 9673 153987 9739 153990
rect 126881 153987 126947 153990
rect 127341 154050 127407 154053
rect 129549 154050 129615 154053
rect 127341 154048 129615 154050
rect 127341 153992 127346 154048
rect 127402 153992 129554 154048
rect 129610 153992 129615 154048
rect 127341 153990 129615 153992
rect 127341 153987 127407 153990
rect 129549 153987 129615 153990
rect 519445 154050 519511 154053
rect 523200 154050 524400 154080
rect 519445 154048 524400 154050
rect 519445 153992 519450 154048
rect 519506 153992 524400 154048
rect 519445 153990 524400 153992
rect 519445 153987 519511 153990
rect 523200 153960 524400 153990
rect 7557 153914 7623 153917
rect 124949 153914 125015 153917
rect 7557 153912 125015 153914
rect 7557 153856 7562 153912
rect 7618 153856 124954 153912
rect 125010 153856 125015 153912
rect 7557 153854 125015 153856
rect 7557 153851 7623 153854
rect 124949 153851 125015 153854
rect 7097 153778 7163 153781
rect 124305 153778 124371 153781
rect 7097 153776 124371 153778
rect 7097 153720 7102 153776
rect 7158 153720 124310 153776
rect 124366 153720 124371 153776
rect 7097 153718 124371 153720
rect 7097 153715 7163 153718
rect 124305 153715 124371 153718
rect 124489 153778 124555 153781
rect 200113 153778 200179 153781
rect 124489 153776 200179 153778
rect 124489 153720 124494 153776
rect 124550 153720 200118 153776
rect 200174 153720 200179 153776
rect 124489 153718 200179 153720
rect 124489 153715 124555 153718
rect 200113 153715 200179 153718
rect 221273 153778 221339 153781
rect 288709 153778 288775 153781
rect 221273 153776 288775 153778
rect 221273 153720 221278 153776
rect 221334 153720 288714 153776
rect 288770 153720 288775 153776
rect 221273 153718 288775 153720
rect 221273 153715 221339 153718
rect 288709 153715 288775 153718
rect 189717 153642 189783 153645
rect 191281 153642 191347 153645
rect 189717 153640 191347 153642
rect 189717 153584 189722 153640
rect 189778 153584 191286 153640
rect 191342 153584 191347 153640
rect 189717 153582 191347 153584
rect 189717 153579 189783 153582
rect 191281 153579 191347 153582
rect 189441 153370 189507 153373
rect 191281 153370 191347 153373
rect 189441 153368 191347 153370
rect 189441 153312 189446 153368
rect 189502 153312 191286 153368
rect 191342 153312 191347 153368
rect 189441 153310 191347 153312
rect 189441 153307 189507 153310
rect 191281 153307 191347 153310
rect 274541 153370 274607 153373
rect 275921 153370 275987 153373
rect 274541 153368 275987 153370
rect 274541 153312 274546 153368
rect 274602 153312 275926 153368
rect 275982 153312 275987 153368
rect 274541 153310 275987 153312
rect 274541 153307 274607 153310
rect 275921 153307 275987 153310
rect 118693 153098 118759 153101
rect 121085 153098 121151 153101
rect 118693 153096 121151 153098
rect 118693 153040 118698 153096
rect 118754 153040 121090 153096
rect 121146 153040 121151 153096
rect 118693 153038 121151 153040
rect 118693 153035 118759 153038
rect 121085 153035 121151 153038
rect 123845 153098 123911 153101
rect 126237 153098 126303 153101
rect 123845 153096 126303 153098
rect 123845 153040 123850 153096
rect 123906 153040 126242 153096
rect 126298 153040 126303 153096
rect 123845 153038 126303 153040
rect 123845 153035 123911 153038
rect 126237 153035 126303 153038
rect 132861 153098 132927 153101
rect 141049 153098 141115 153101
rect 132861 153096 141115 153098
rect 132861 153040 132866 153096
rect 132922 153040 141054 153096
rect 141110 153040 141115 153096
rect 132861 153038 141115 153040
rect 132861 153035 132927 153038
rect 141049 153035 141115 153038
rect 24853 152690 24919 152693
rect 138473 152690 138539 152693
rect 24853 152688 138539 152690
rect 24853 152632 24858 152688
rect 24914 152632 138478 152688
rect 138534 152632 138539 152688
rect 24853 152630 138539 152632
rect 24853 152627 24919 152630
rect 138473 152627 138539 152630
rect 446949 152690 447015 152693
rect 447409 152690 447475 152693
rect 446949 152688 447475 152690
rect 446949 152632 446954 152688
rect 447010 152632 447414 152688
rect 447470 152632 447475 152688
rect 446949 152630 447475 152632
rect 446949 152627 447015 152630
rect 447409 152627 447475 152630
rect 19333 152554 19399 152557
rect 133965 152554 134031 152557
rect 19333 152552 134031 152554
rect 19333 152496 19338 152552
rect 19394 152496 133970 152552
rect 134026 152496 134031 152552
rect 19333 152494 134031 152496
rect 19333 152491 19399 152494
rect 133965 152491 134031 152494
rect 521009 152554 521075 152557
rect 523200 152554 524400 152584
rect 521009 152552 524400 152554
rect 521009 152496 521014 152552
rect 521070 152496 524400 152552
rect 521009 152494 524400 152496
rect 521009 152491 521075 152494
rect 523200 152464 524400 152494
rect 5533 152418 5599 152421
rect 123661 152418 123727 152421
rect 5533 152416 123727 152418
rect 5533 152360 5538 152416
rect 5594 152360 123666 152416
rect 123722 152360 123727 152416
rect 5533 152358 123727 152360
rect 5533 152355 5599 152358
rect 123661 152355 123727 152358
rect 217133 152418 217199 152421
rect 285489 152418 285555 152421
rect 217133 152416 285555 152418
rect 217133 152360 217138 152416
rect 217194 152360 285494 152416
rect 285550 152360 285555 152416
rect 217133 152358 285555 152360
rect 217133 152355 217199 152358
rect 285489 152355 285555 152358
rect 310697 152418 310763 152421
rect 356145 152418 356211 152421
rect 310697 152416 356211 152418
rect 310697 152360 310702 152416
rect 310758 152360 356150 152416
rect 356206 152360 356211 152416
rect 310697 152358 356211 152360
rect 310697 152355 310763 152358
rect 356145 152355 356211 152358
rect 432873 152418 432939 152421
rect 449893 152418 449959 152421
rect 432873 152416 449959 152418
rect 432873 152360 432878 152416
rect 432934 152360 449898 152416
rect 449954 152360 449959 152416
rect 432873 152358 449959 152360
rect 432873 152355 432939 152358
rect 449893 152355 449959 152358
rect 446581 152010 446647 152013
rect 448053 152010 448119 152013
rect 446581 152008 448119 152010
rect 446581 151952 446586 152008
rect 446642 151952 448058 152008
rect 448114 151952 448119 152008
rect 446581 151950 448119 151952
rect 446581 151947 446647 151950
rect 448053 151947 448119 151950
rect 445661 151874 445727 151877
rect 447041 151874 447107 151877
rect 445661 151872 447107 151874
rect 445661 151816 445666 151872
rect 445722 151816 447046 151872
rect 447102 151816 447107 151872
rect 445661 151814 447107 151816
rect 445661 151811 445727 151814
rect 447041 151811 447107 151814
rect 520181 151058 520247 151061
rect 523200 151058 524400 151088
rect 520181 151056 524400 151058
rect 520181 151000 520186 151056
rect 520242 151000 524400 151056
rect 520181 150998 524400 151000
rect 520181 150995 520247 150998
rect 523200 150968 524400 150998
rect 6085 150650 6151 150653
rect 111333 150650 111399 150653
rect 6085 150648 111399 150650
rect 6085 150592 6090 150648
rect 6146 150592 111338 150648
rect 111394 150592 111399 150648
rect 6085 150590 111399 150592
rect 6085 150587 6151 150590
rect 111333 150587 111399 150590
rect 2681 150514 2747 150517
rect 111057 150514 111123 150517
rect 2681 150512 111123 150514
rect 2681 150456 2686 150512
rect 2742 150456 111062 150512
rect 111118 150456 111123 150512
rect 2681 150454 111123 150456
rect 2681 150451 2747 150454
rect 111057 150451 111123 150454
rect 99925 149834 99991 149837
rect 116853 149834 116919 149837
rect 99925 149832 116919 149834
rect 99925 149776 99930 149832
rect 99986 149776 116858 149832
rect 116914 149776 116919 149832
rect 99925 149774 116919 149776
rect 99925 149771 99991 149774
rect 116853 149771 116919 149774
rect 92565 149698 92631 149701
rect 116577 149698 116643 149701
rect 92565 149696 116643 149698
rect 92565 149640 92570 149696
rect 92626 149640 116582 149696
rect 116638 149640 116643 149696
rect 92565 149638 116643 149640
rect 92565 149635 92631 149638
rect 116577 149635 116643 149638
rect 520089 149562 520155 149565
rect 523200 149562 524400 149592
rect 520089 149560 524400 149562
rect 520089 149504 520094 149560
rect 520150 149504 524400 149560
rect 520089 149502 524400 149504
rect 520089 149499 520155 149502
rect 523200 149472 524400 149502
rect 519721 149290 519787 149293
rect 518788 149288 519787 149290
rect 518788 149232 519726 149288
rect 519782 149232 519787 149288
rect 518788 149230 519787 149232
rect 519721 149227 519787 149230
rect 109585 148066 109651 148069
rect 119110 148066 119170 148988
rect 109585 148064 119170 148066
rect 109585 148008 109590 148064
rect 109646 148008 119170 148064
rect 109585 148006 119170 148008
rect 519721 148066 519787 148069
rect 523200 148066 524400 148096
rect 519721 148064 524400 148066
rect 519721 148008 519726 148064
rect 519782 148008 524400 148064
rect 519721 148006 524400 148008
rect 109585 148003 109651 148006
rect 519721 148003 519787 148006
rect 523200 147976 524400 148006
rect 519537 147930 519603 147933
rect 518788 147928 519603 147930
rect 518788 147872 519542 147928
rect 519598 147872 519603 147928
rect 518788 147870 519603 147872
rect 519537 147867 519603 147870
rect 110965 147386 111031 147389
rect 111701 147386 111767 147389
rect 110965 147384 111767 147386
rect 110965 147328 110970 147384
rect 111026 147328 111706 147384
rect 111762 147328 111767 147384
rect 110965 147326 111767 147328
rect 110965 147323 111031 147326
rect 111701 147323 111767 147326
rect 110321 146434 110387 146437
rect 119110 146434 119170 147084
rect 519629 146570 519695 146573
rect 518788 146568 519695 146570
rect 518788 146512 519634 146568
rect 519690 146512 519695 146568
rect 518788 146510 519695 146512
rect 519629 146507 519695 146510
rect 520917 146570 520983 146573
rect 523200 146570 524400 146600
rect 520917 146568 524400 146570
rect 520917 146512 520922 146568
rect 520978 146512 524400 146568
rect 520917 146510 524400 146512
rect 520917 146507 520983 146510
rect 523200 146480 524400 146510
rect 110321 146432 119170 146434
rect 110321 146376 110326 146432
rect 110382 146376 119170 146432
rect 110321 146374 119170 146376
rect 110321 146371 110387 146374
rect 116117 145210 116183 145213
rect 519997 145210 520063 145213
rect 116117 145208 119140 145210
rect 116117 145152 116122 145208
rect 116178 145152 119140 145208
rect 116117 145150 119140 145152
rect 518788 145208 520063 145210
rect 518788 145152 520002 145208
rect 520058 145152 520063 145208
rect 518788 145150 520063 145152
rect 116117 145147 116183 145150
rect 519997 145147 520063 145150
rect 519537 144938 519603 144941
rect 523200 144938 524400 144968
rect 519537 144936 524400 144938
rect 519537 144880 519542 144936
rect 519598 144880 524400 144936
rect 519537 144878 524400 144880
rect 519537 144875 519603 144878
rect 523200 144848 524400 144878
rect 113817 144258 113883 144261
rect 110860 144256 113883 144258
rect 110860 144200 113822 144256
rect 113878 144200 113883 144256
rect 110860 144198 113883 144200
rect 113817 144195 113883 144198
rect 519905 143850 519971 143853
rect 518788 143848 519971 143850
rect 518788 143792 519910 143848
rect 519966 143792 519971 143848
rect 518788 143790 519971 143792
rect 519905 143787 519971 143790
rect 519997 143442 520063 143445
rect 523200 143442 524400 143472
rect 519997 143440 524400 143442
rect 519997 143384 520002 143440
rect 520058 143384 524400 143440
rect 519997 143382 524400 143384
rect 519997 143379 520063 143382
rect 523200 143352 524400 143382
rect 116025 143306 116091 143309
rect 116025 143304 119140 143306
rect 116025 143248 116030 143304
rect 116086 143248 119140 143304
rect 116025 143246 119140 143248
rect 116025 143243 116091 143246
rect 519813 142490 519879 142493
rect 518788 142488 519879 142490
rect 518788 142432 519818 142488
rect 519874 142432 519879 142488
rect 518788 142430 519879 142432
rect 519813 142427 519879 142430
rect 519169 141946 519235 141949
rect 523200 141946 524400 141976
rect 519169 141944 524400 141946
rect 519169 141888 519174 141944
rect 519230 141888 524400 141944
rect 519169 141886 524400 141888
rect 519169 141883 519235 141886
rect 523200 141856 524400 141886
rect 115289 141402 115355 141405
rect 115289 141400 119140 141402
rect 115289 141344 115294 141400
rect 115350 141344 119140 141400
rect 115289 141342 119140 141344
rect 115289 141339 115355 141342
rect 519445 141130 519511 141133
rect 518788 141128 519511 141130
rect 518788 141072 519450 141128
rect 519506 141072 519511 141128
rect 518788 141070 519511 141072
rect 519445 141067 519511 141070
rect 519261 140450 519327 140453
rect 523200 140450 524400 140480
rect 519261 140448 524400 140450
rect 519261 140392 519266 140448
rect 519322 140392 524400 140448
rect 519261 140390 524400 140392
rect 519261 140387 519327 140390
rect 523200 140360 524400 140390
rect 521009 139770 521075 139773
rect 518788 139768 521075 139770
rect 518788 139712 521014 139768
rect 521070 139712 521075 139768
rect 518788 139710 521075 139712
rect 521009 139707 521075 139710
rect 116117 139498 116183 139501
rect 116117 139496 119140 139498
rect 116117 139440 116122 139496
rect 116178 139440 119140 139496
rect 116117 139438 119140 139440
rect 116117 139435 116183 139438
rect 519353 138954 519419 138957
rect 523200 138954 524400 138984
rect 519353 138952 524400 138954
rect 519353 138896 519358 138952
rect 519414 138896 524400 138952
rect 519353 138894 524400 138896
rect 519353 138891 519419 138894
rect 523200 138864 524400 138894
rect 520181 138410 520247 138413
rect 518788 138408 520247 138410
rect 518788 138352 520186 138408
rect 520242 138352 520247 138408
rect 518788 138350 520247 138352
rect 520181 138347 520247 138350
rect 116117 137594 116183 137597
rect 116117 137592 119140 137594
rect 116117 137536 116122 137592
rect 116178 137536 119140 137592
rect 116117 137534 119140 137536
rect 116117 137531 116183 137534
rect 519445 137458 519511 137461
rect 523200 137458 524400 137488
rect 519445 137456 524400 137458
rect 519445 137400 519450 137456
rect 519506 137400 524400 137456
rect 519445 137398 524400 137400
rect 519445 137395 519511 137398
rect 523200 137368 524400 137398
rect 520089 137050 520155 137053
rect 518788 137048 520155 137050
rect 518788 136992 520094 137048
rect 520150 136992 520155 137048
rect 518788 136990 520155 136992
rect 520089 136987 520155 136990
rect 519905 135826 519971 135829
rect 523200 135826 524400 135856
rect 519905 135824 524400 135826
rect 519905 135768 519910 135824
rect 519966 135768 524400 135824
rect 519905 135766 524400 135768
rect 519905 135763 519971 135766
rect 523200 135736 524400 135766
rect 519721 135690 519787 135693
rect 518788 135688 519787 135690
rect 518788 135632 519726 135688
rect 519782 135632 519787 135688
rect 518788 135630 519787 135632
rect 519721 135627 519787 135630
rect 115197 135554 115263 135557
rect 115197 135552 119140 135554
rect 115197 135496 115202 135552
rect 115258 135496 119140 135552
rect 115197 135494 119140 135496
rect 115197 135491 115263 135494
rect 520917 134466 520983 134469
rect 518758 134464 520983 134466
rect 518758 134408 520922 134464
rect 520978 134408 520983 134464
rect 518758 134406 520983 134408
rect 518758 134300 518818 134406
rect 520917 134403 520983 134406
rect 519813 134330 519879 134333
rect 523200 134330 524400 134360
rect 519813 134328 524400 134330
rect 519813 134272 519818 134328
rect 519874 134272 524400 134328
rect 519813 134270 524400 134272
rect 519813 134267 519879 134270
rect 523200 134240 524400 134270
rect 116025 133650 116091 133653
rect 116025 133648 119140 133650
rect 116025 133592 116030 133648
rect 116086 133592 119140 133648
rect 116025 133590 119140 133592
rect 116025 133587 116091 133590
rect 519537 132970 519603 132973
rect 518788 132968 519603 132970
rect 518788 132912 519542 132968
rect 519598 132912 519603 132968
rect 518788 132910 519603 132912
rect 519537 132907 519603 132910
rect 114185 132834 114251 132837
rect 110860 132832 114251 132834
rect 110860 132776 114190 132832
rect 114246 132776 114251 132832
rect 110860 132774 114251 132776
rect 114185 132771 114251 132774
rect 519721 132834 519787 132837
rect 523200 132834 524400 132864
rect 519721 132832 524400 132834
rect 519721 132776 519726 132832
rect 519782 132776 524400 132832
rect 519721 132774 524400 132776
rect 519721 132771 519787 132774
rect 523200 132744 524400 132774
rect 116117 131746 116183 131749
rect 116117 131744 119140 131746
rect 116117 131688 116122 131744
rect 116178 131688 119140 131744
rect 116117 131686 119140 131688
rect 116117 131683 116183 131686
rect 519997 131610 520063 131613
rect 518788 131608 520063 131610
rect 518788 131552 520002 131608
rect 520058 131552 520063 131608
rect 518788 131550 520063 131552
rect 519997 131547 520063 131550
rect 519629 131338 519695 131341
rect 523200 131338 524400 131368
rect 519629 131336 524400 131338
rect 519629 131280 519634 131336
rect 519690 131280 524400 131336
rect 519629 131278 524400 131280
rect 519629 131275 519695 131278
rect 523200 131248 524400 131278
rect 519169 130250 519235 130253
rect 518788 130248 519235 130250
rect 518788 130192 519174 130248
rect 519230 130192 519235 130248
rect 518788 130190 519235 130192
rect 519169 130187 519235 130190
rect 116393 129842 116459 129845
rect 519537 129842 519603 129845
rect 523200 129842 524400 129872
rect 116393 129840 119140 129842
rect 116393 129784 116398 129840
rect 116454 129784 119140 129840
rect 116393 129782 119140 129784
rect 519537 129840 524400 129842
rect 519537 129784 519542 129840
rect 519598 129784 524400 129840
rect 519537 129782 524400 129784
rect 116393 129779 116459 129782
rect 519537 129779 519603 129782
rect 523200 129752 524400 129782
rect 519261 128890 519327 128893
rect 518788 128888 519327 128890
rect 518788 128832 519266 128888
rect 519322 128832 519327 128888
rect 518788 128830 519327 128832
rect 519261 128827 519327 128830
rect 519169 128346 519235 128349
rect 523200 128346 524400 128376
rect 519169 128344 524400 128346
rect 519169 128288 519174 128344
rect 519230 128288 524400 128344
rect 519169 128286 524400 128288
rect 519169 128283 519235 128286
rect 523200 128256 524400 128286
rect 116301 127938 116367 127941
rect 116301 127936 119140 127938
rect 116301 127880 116306 127936
rect 116362 127880 119140 127936
rect 116301 127878 119140 127880
rect 116301 127875 116367 127878
rect 519353 127530 519419 127533
rect 518788 127528 519419 127530
rect 518788 127472 519358 127528
rect 519414 127472 519419 127528
rect 518788 127470 519419 127472
rect 519353 127467 519419 127470
rect 519261 126714 519327 126717
rect 523200 126714 524400 126744
rect 519261 126712 524400 126714
rect 519261 126656 519266 126712
rect 519322 126656 524400 126712
rect 519261 126654 524400 126656
rect 519261 126651 519327 126654
rect 523200 126624 524400 126654
rect 519445 126170 519511 126173
rect 518788 126168 519511 126170
rect 518788 126112 519450 126168
rect 519506 126112 519511 126168
rect 518788 126110 519511 126112
rect 519445 126107 519511 126110
rect 116025 126034 116091 126037
rect 116025 126032 119140 126034
rect 116025 125976 116030 126032
rect 116086 125976 119140 126032
rect 116025 125974 119140 125976
rect 116025 125971 116091 125974
rect 520181 125218 520247 125221
rect 523200 125218 524400 125248
rect 520181 125216 524400 125218
rect 520181 125160 520186 125216
rect 520242 125160 524400 125216
rect 520181 125158 524400 125160
rect 520181 125155 520247 125158
rect 523200 125128 524400 125158
rect 519905 124810 519971 124813
rect 518788 124808 519971 124810
rect 518788 124752 519910 124808
rect 519966 124752 519971 124808
rect 518788 124750 519971 124752
rect 519905 124747 519971 124750
rect 116117 124130 116183 124133
rect 116117 124128 119140 124130
rect 116117 124072 116122 124128
rect 116178 124072 119140 124128
rect 116117 124070 119140 124072
rect 116117 124067 116183 124070
rect 520089 123722 520155 123725
rect 523200 123722 524400 123752
rect 520089 123720 524400 123722
rect 520089 123664 520094 123720
rect 520150 123664 524400 123720
rect 520089 123662 524400 123664
rect 520089 123659 520155 123662
rect 523200 123632 524400 123662
rect 519813 123450 519879 123453
rect 518788 123448 519879 123450
rect 518788 123392 519818 123448
rect 519874 123392 519879 123448
rect 518788 123390 519879 123392
rect 519813 123387 519879 123390
rect 115933 122226 115999 122229
rect 519905 122226 519971 122229
rect 523200 122226 524400 122256
rect 115933 122224 119140 122226
rect 115933 122168 115938 122224
rect 115994 122168 119140 122224
rect 115933 122166 119140 122168
rect 519905 122224 524400 122226
rect 519905 122168 519910 122224
rect 519966 122168 524400 122224
rect 519905 122166 524400 122168
rect 115933 122163 115999 122166
rect 519905 122163 519971 122166
rect 523200 122136 524400 122166
rect 519721 122090 519787 122093
rect 518788 122088 519787 122090
rect 518788 122032 519726 122088
rect 519782 122032 519787 122088
rect 518788 122030 519787 122032
rect 519721 122027 519787 122030
rect 113909 121410 113975 121413
rect 110860 121408 113975 121410
rect 110860 121352 113914 121408
rect 113970 121352 113975 121408
rect 110860 121350 113975 121352
rect 113909 121347 113975 121350
rect 519629 120730 519695 120733
rect 518788 120728 519695 120730
rect 518788 120672 519634 120728
rect 519690 120672 519695 120728
rect 518788 120670 519695 120672
rect 519629 120667 519695 120670
rect 519813 120730 519879 120733
rect 523200 120730 524400 120760
rect 519813 120728 524400 120730
rect 519813 120672 519818 120728
rect 519874 120672 524400 120728
rect 519813 120670 524400 120672
rect 519813 120667 519879 120670
rect 523200 120640 524400 120670
rect 116117 120186 116183 120189
rect 116117 120184 119140 120186
rect 116117 120128 116122 120184
rect 116178 120128 119140 120184
rect 116117 120126 119140 120128
rect 116117 120123 116183 120126
rect 519537 119370 519603 119373
rect 518788 119368 519603 119370
rect 518788 119312 519542 119368
rect 519598 119312 519603 119368
rect 518788 119310 519603 119312
rect 519537 119307 519603 119310
rect 519721 119234 519787 119237
rect 523200 119234 524400 119264
rect 519721 119232 524400 119234
rect 519721 119176 519726 119232
rect 519782 119176 524400 119232
rect 519721 119174 524400 119176
rect 519721 119171 519787 119174
rect 523200 119144 524400 119174
rect 116117 118282 116183 118285
rect 116117 118280 119140 118282
rect 116117 118224 116122 118280
rect 116178 118224 119140 118280
rect 116117 118222 119140 118224
rect 116117 118219 116183 118222
rect 519169 118010 519235 118013
rect 518788 118008 519235 118010
rect 518788 117952 519174 118008
rect 519230 117952 519235 118008
rect 518788 117950 519235 117952
rect 519169 117947 519235 117950
rect 519997 117602 520063 117605
rect 523200 117602 524400 117632
rect 519997 117600 524400 117602
rect 519997 117544 520002 117600
rect 520058 117544 524400 117600
rect 519997 117542 524400 117544
rect 519997 117539 520063 117542
rect 523200 117512 524400 117542
rect 519261 116650 519327 116653
rect 518788 116648 519327 116650
rect 518788 116592 519266 116648
rect 519322 116592 519327 116648
rect 518788 116590 519327 116592
rect 519261 116587 519327 116590
rect 116117 116378 116183 116381
rect 116117 116376 119140 116378
rect 116117 116320 116122 116376
rect 116178 116320 119140 116376
rect 116117 116318 119140 116320
rect 116117 116315 116183 116318
rect 519629 116106 519695 116109
rect 523200 116106 524400 116136
rect 519629 116104 524400 116106
rect 519629 116048 519634 116104
rect 519690 116048 524400 116104
rect 519629 116046 524400 116048
rect 519629 116043 519695 116046
rect 523200 116016 524400 116046
rect 520181 115290 520247 115293
rect 518788 115288 520247 115290
rect 518788 115232 520186 115288
rect 520242 115232 520247 115288
rect 518788 115230 520247 115232
rect 520181 115227 520247 115230
rect 519537 114610 519603 114613
rect 523200 114610 524400 114640
rect 519537 114608 524400 114610
rect 519537 114552 519542 114608
rect 519598 114552 524400 114608
rect 519537 114550 524400 114552
rect 519537 114547 519603 114550
rect 523200 114520 524400 114550
rect 116117 114474 116183 114477
rect 116117 114472 119140 114474
rect 116117 114416 116122 114472
rect 116178 114416 119140 114472
rect 116117 114414 119140 114416
rect 116117 114411 116183 114414
rect 520089 113930 520155 113933
rect 518788 113928 520155 113930
rect 518788 113872 520094 113928
rect 520150 113872 520155 113928
rect 518788 113870 520155 113872
rect 520089 113867 520155 113870
rect 520917 113114 520983 113117
rect 523200 113114 524400 113144
rect 520917 113112 524400 113114
rect 520917 113056 520922 113112
rect 520978 113056 524400 113112
rect 520917 113054 524400 113056
rect 520917 113051 520983 113054
rect 523200 113024 524400 113054
rect 115933 112570 115999 112573
rect 519905 112570 519971 112573
rect 115933 112568 119140 112570
rect 115933 112512 115938 112568
rect 115994 112512 119140 112568
rect 115933 112510 119140 112512
rect 518788 112568 519971 112570
rect 518788 112512 519910 112568
rect 519966 112512 519971 112568
rect 518788 112510 519971 112512
rect 115933 112507 115999 112510
rect 519905 112507 519971 112510
rect 521285 111618 521351 111621
rect 523200 111618 524400 111648
rect 521285 111616 524400 111618
rect 521285 111560 521290 111616
rect 521346 111560 524400 111616
rect 521285 111558 524400 111560
rect 521285 111555 521351 111558
rect 523200 111528 524400 111558
rect 519813 111210 519879 111213
rect 518788 111208 519879 111210
rect 518788 111152 519818 111208
rect 519874 111152 519879 111208
rect 518788 111150 519879 111152
rect 519813 111147 519879 111150
rect 116117 110666 116183 110669
rect 116117 110664 119140 110666
rect 116117 110608 116122 110664
rect 116178 110608 119140 110664
rect 116117 110606 119140 110608
rect 116117 110603 116183 110606
rect 114001 110122 114067 110125
rect 110860 110120 114067 110122
rect 110860 110064 114006 110120
rect 114062 110064 114067 110120
rect 110860 110062 114067 110064
rect 114001 110059 114067 110062
rect 521469 110122 521535 110125
rect 523200 110122 524400 110152
rect 521469 110120 524400 110122
rect 521469 110064 521474 110120
rect 521530 110064 524400 110120
rect 521469 110062 524400 110064
rect 521469 110059 521535 110062
rect 523200 110032 524400 110062
rect 519721 109850 519787 109853
rect 518788 109848 519787 109850
rect 518788 109792 519726 109848
rect 519782 109792 519787 109848
rect 518788 109790 519787 109792
rect 519721 109787 519787 109790
rect 116117 108762 116183 108765
rect 116117 108760 119140 108762
rect 116117 108704 116122 108760
rect 116178 108704 119140 108760
rect 116117 108702 119140 108704
rect 116117 108699 116183 108702
rect 519997 108490 520063 108493
rect 518788 108488 520063 108490
rect 518788 108432 520002 108488
rect 520058 108432 520063 108488
rect 518788 108430 520063 108432
rect 519997 108427 520063 108430
rect 521377 108490 521443 108493
rect 523200 108490 524400 108520
rect 521377 108488 524400 108490
rect 521377 108432 521382 108488
rect 521438 108432 524400 108488
rect 521377 108430 524400 108432
rect 521377 108427 521443 108430
rect 523200 108400 524400 108430
rect 519629 107130 519695 107133
rect 518788 107128 519695 107130
rect 518788 107072 519634 107128
rect 519690 107072 519695 107128
rect 518788 107070 519695 107072
rect 519629 107067 519695 107070
rect 521193 106994 521259 106997
rect 523200 106994 524400 107024
rect 521193 106992 524400 106994
rect 521193 106936 521198 106992
rect 521254 106936 524400 106992
rect 521193 106934 524400 106936
rect 521193 106931 521259 106934
rect 523200 106904 524400 106934
rect 116485 106858 116551 106861
rect 116485 106856 119140 106858
rect 116485 106800 116490 106856
rect 116546 106800 119140 106856
rect 116485 106798 119140 106800
rect 116485 106795 116551 106798
rect 519537 105770 519603 105773
rect 518788 105768 519603 105770
rect 518788 105712 519542 105768
rect 519598 105712 519603 105768
rect 518788 105710 519603 105712
rect 519537 105707 519603 105710
rect 520273 105498 520339 105501
rect 523200 105498 524400 105528
rect 520273 105496 524400 105498
rect 520273 105440 520278 105496
rect 520334 105440 524400 105496
rect 520273 105438 524400 105440
rect 520273 105435 520339 105438
rect 523200 105408 524400 105438
rect 117129 104818 117195 104821
rect 117129 104816 119140 104818
rect 117129 104760 117134 104816
rect 117190 104760 119140 104816
rect 117129 104758 119140 104760
rect 117129 104755 117195 104758
rect 520917 104410 520983 104413
rect 518788 104408 520983 104410
rect 518788 104352 520922 104408
rect 520978 104352 520983 104408
rect 518788 104350 520983 104352
rect 520917 104347 520983 104350
rect 521101 104002 521167 104005
rect 523200 104002 524400 104032
rect 521101 104000 524400 104002
rect 521101 103944 521106 104000
rect 521162 103944 524400 104000
rect 521101 103942 524400 103944
rect 521101 103939 521167 103942
rect 523200 103912 524400 103942
rect 521285 103050 521351 103053
rect 518788 103048 521351 103050
rect 518788 102992 521290 103048
rect 521346 102992 521351 103048
rect 518788 102990 521351 102992
rect 521285 102987 521351 102990
rect 116945 102914 117011 102917
rect 116945 102912 119140 102914
rect 116945 102856 116950 102912
rect 117006 102856 119140 102912
rect 116945 102854 119140 102856
rect 116945 102851 117011 102854
rect 521009 102506 521075 102509
rect 523200 102506 524400 102536
rect 521009 102504 524400 102506
rect 521009 102448 521014 102504
rect 521070 102448 524400 102504
rect 521009 102446 524400 102448
rect 521009 102443 521075 102446
rect 523200 102416 524400 102446
rect 521469 101690 521535 101693
rect 518788 101688 521535 101690
rect 518788 101632 521474 101688
rect 521530 101632 521535 101688
rect 518788 101630 521535 101632
rect 521469 101627 521535 101630
rect 117037 101010 117103 101013
rect 521285 101010 521351 101013
rect 523200 101010 524400 101040
rect 117037 101008 119140 101010
rect 117037 100952 117042 101008
rect 117098 100952 119140 101008
rect 117037 100950 119140 100952
rect 521285 101008 524400 101010
rect 521285 100952 521290 101008
rect 521346 100952 524400 101008
rect 521285 100950 524400 100952
rect 117037 100947 117103 100950
rect 521285 100947 521351 100950
rect 523200 100920 524400 100950
rect 521377 100330 521443 100333
rect 518788 100328 521443 100330
rect 518788 100272 521382 100328
rect 521438 100272 521443 100328
rect 518788 100270 521443 100272
rect 521377 100267 521443 100270
rect 519813 99378 519879 99381
rect 523200 99378 524400 99408
rect 519813 99376 524400 99378
rect 519813 99320 519818 99376
rect 519874 99320 524400 99376
rect 519813 99318 524400 99320
rect 519813 99315 519879 99318
rect 523200 99288 524400 99318
rect 116853 99106 116919 99109
rect 116853 99104 119140 99106
rect 116853 99048 116858 99104
rect 116914 99048 119140 99104
rect 116853 99046 119140 99048
rect 116853 99043 116919 99046
rect 521193 98970 521259 98973
rect 518788 98968 521259 98970
rect 518788 98912 521198 98968
rect 521254 98912 521259 98968
rect 518788 98910 521259 98912
rect 521193 98907 521259 98910
rect 114093 98698 114159 98701
rect 110860 98696 114159 98698
rect 110860 98640 114098 98696
rect 114154 98640 114159 98696
rect 110860 98638 114159 98640
rect 114093 98635 114159 98638
rect 519721 97882 519787 97885
rect 523200 97882 524400 97912
rect 519721 97880 524400 97882
rect 519721 97824 519726 97880
rect 519782 97824 524400 97880
rect 519721 97822 524400 97824
rect 519721 97819 519787 97822
rect 523200 97792 524400 97822
rect 520273 97610 520339 97613
rect 518788 97608 520339 97610
rect 518788 97552 520278 97608
rect 520334 97552 520339 97608
rect 518788 97550 520339 97552
rect 520273 97547 520339 97550
rect 116761 97202 116827 97205
rect 116761 97200 119140 97202
rect 116761 97144 116766 97200
rect 116822 97144 119140 97200
rect 116761 97142 119140 97144
rect 116761 97139 116827 97142
rect 519997 96386 520063 96389
rect 523200 96386 524400 96416
rect 519997 96384 524400 96386
rect 519997 96328 520002 96384
rect 520058 96328 524400 96384
rect 519997 96326 524400 96328
rect 519997 96323 520063 96326
rect 523200 96296 524400 96326
rect 521101 96250 521167 96253
rect 518788 96248 521167 96250
rect 518788 96192 521106 96248
rect 521162 96192 521167 96248
rect 518788 96190 521167 96192
rect 521101 96187 521167 96190
rect 116669 95298 116735 95301
rect 116669 95296 119140 95298
rect 116669 95240 116674 95296
rect 116730 95240 119140 95296
rect 116669 95238 119140 95240
rect 116669 95235 116735 95238
rect 521009 95026 521075 95029
rect 518758 95024 521075 95026
rect 518758 94968 521014 95024
rect 521070 94968 521075 95024
rect 518758 94966 521075 94968
rect 518758 94860 518818 94966
rect 521009 94963 521075 94966
rect 519905 94890 519971 94893
rect 523200 94890 524400 94920
rect 519905 94888 524400 94890
rect 519905 94832 519910 94888
rect 519966 94832 524400 94888
rect 519905 94830 524400 94832
rect 519905 94827 519971 94830
rect 523200 94800 524400 94830
rect 521285 93530 521351 93533
rect 518788 93528 521351 93530
rect 518788 93472 521290 93528
rect 521346 93472 521351 93528
rect 518788 93470 521351 93472
rect 521285 93467 521351 93470
rect 116577 93394 116643 93397
rect 520365 93394 520431 93397
rect 523200 93394 524400 93424
rect 116577 93392 119140 93394
rect 116577 93336 116582 93392
rect 116638 93336 119140 93392
rect 116577 93334 119140 93336
rect 520365 93392 524400 93394
rect 520365 93336 520370 93392
rect 520426 93336 524400 93392
rect 520365 93334 524400 93336
rect 116577 93331 116643 93334
rect 520365 93331 520431 93334
rect 523200 93304 524400 93334
rect 519813 92170 519879 92173
rect 518788 92168 519879 92170
rect 518788 92112 519818 92168
rect 519874 92112 519879 92168
rect 518788 92110 519879 92112
rect 519813 92107 519879 92110
rect 521377 91898 521443 91901
rect 523200 91898 524400 91928
rect 521377 91896 524400 91898
rect 521377 91840 521382 91896
rect 521438 91840 524400 91896
rect 521377 91838 524400 91840
rect 521377 91835 521443 91838
rect 523200 91808 524400 91838
rect 116117 91354 116183 91357
rect 116117 91352 119140 91354
rect 116117 91296 116122 91352
rect 116178 91296 119140 91352
rect 116117 91294 119140 91296
rect 116117 91291 116183 91294
rect 519721 90810 519787 90813
rect 518788 90808 519787 90810
rect 518788 90752 519726 90808
rect 519782 90752 519787 90808
rect 518788 90750 519787 90752
rect 519721 90747 519787 90750
rect 521193 90266 521259 90269
rect 523200 90266 524400 90296
rect 521193 90264 524400 90266
rect 521193 90208 521198 90264
rect 521254 90208 524400 90264
rect 521193 90206 524400 90208
rect 521193 90203 521259 90206
rect 523200 90176 524400 90206
rect 116117 89450 116183 89453
rect 519997 89450 520063 89453
rect 116117 89448 119140 89450
rect 116117 89392 116122 89448
rect 116178 89392 119140 89448
rect 116117 89390 119140 89392
rect 518788 89448 520063 89450
rect 518788 89392 520002 89448
rect 520058 89392 520063 89448
rect 518788 89390 520063 89392
rect 116117 89387 116183 89390
rect 519997 89387 520063 89390
rect 521285 88770 521351 88773
rect 523200 88770 524400 88800
rect 521285 88768 524400 88770
rect 521285 88712 521290 88768
rect 521346 88712 524400 88768
rect 521285 88710 524400 88712
rect 521285 88707 521351 88710
rect 523200 88680 524400 88710
rect 519905 88090 519971 88093
rect 518788 88088 519971 88090
rect 518788 88032 519910 88088
rect 519966 88032 519971 88088
rect 518788 88030 519971 88032
rect 519905 88027 519971 88030
rect 116025 87546 116091 87549
rect 116025 87544 119140 87546
rect 116025 87488 116030 87544
rect 116086 87488 119140 87544
rect 116025 87486 119140 87488
rect 116025 87483 116091 87486
rect 114185 87274 114251 87277
rect 110860 87272 114251 87274
rect 110860 87216 114190 87272
rect 114246 87216 114251 87272
rect 110860 87214 114251 87216
rect 114185 87211 114251 87214
rect 521101 87274 521167 87277
rect 523200 87274 524400 87304
rect 521101 87272 524400 87274
rect 521101 87216 521106 87272
rect 521162 87216 524400 87272
rect 521101 87214 524400 87216
rect 521101 87211 521167 87214
rect 523200 87184 524400 87214
rect 521561 86730 521627 86733
rect 518788 86728 521627 86730
rect 518788 86672 521566 86728
rect 521622 86672 521627 86728
rect 518788 86670 521627 86672
rect 521561 86667 521627 86670
rect 520273 85778 520339 85781
rect 523200 85778 524400 85808
rect 520273 85776 524400 85778
rect 520273 85720 520278 85776
rect 520334 85720 524400 85776
rect 520273 85718 524400 85720
rect 520273 85715 520339 85718
rect 523200 85688 524400 85718
rect 115197 85642 115263 85645
rect 115197 85640 119140 85642
rect 115197 85584 115202 85640
rect 115258 85584 119140 85640
rect 115197 85582 119140 85584
rect 115197 85579 115263 85582
rect 520365 85370 520431 85373
rect 518788 85368 520431 85370
rect 518788 85312 520370 85368
rect 520426 85312 520431 85368
rect 518788 85310 520431 85312
rect 520365 85307 520431 85310
rect 520917 84282 520983 84285
rect 523200 84282 524400 84312
rect 520917 84280 524400 84282
rect 520917 84224 520922 84280
rect 520978 84224 524400 84280
rect 520917 84222 524400 84224
rect 520917 84219 520983 84222
rect 523200 84192 524400 84222
rect 521377 84010 521443 84013
rect 518788 84008 521443 84010
rect 518788 83952 521382 84008
rect 521438 83952 521443 84008
rect 518788 83950 521443 83952
rect 521377 83947 521443 83950
rect 116577 83738 116643 83741
rect 116577 83736 119140 83738
rect 116577 83680 116582 83736
rect 116638 83680 119140 83736
rect 116577 83678 119140 83680
rect 116577 83675 116643 83678
rect 519905 82786 519971 82789
rect 523200 82786 524400 82816
rect 519905 82784 524400 82786
rect 519905 82728 519910 82784
rect 519966 82728 524400 82784
rect 519905 82726 524400 82728
rect 519905 82723 519971 82726
rect 523200 82696 524400 82726
rect 521193 82650 521259 82653
rect 518788 82648 521259 82650
rect 518788 82592 521198 82648
rect 521254 82592 521259 82648
rect 518788 82590 521259 82592
rect 521193 82587 521259 82590
rect 116209 81834 116275 81837
rect 116209 81832 119140 81834
rect 116209 81776 116214 81832
rect 116270 81776 119140 81832
rect 116209 81774 119140 81776
rect 116209 81771 116275 81774
rect 521285 81290 521351 81293
rect 518788 81288 521351 81290
rect 518788 81232 521290 81288
rect 521346 81232 521351 81288
rect 518788 81230 521351 81232
rect 521285 81227 521351 81230
rect 519629 81154 519695 81157
rect 523200 81154 524400 81184
rect 519629 81152 524400 81154
rect 519629 81096 519634 81152
rect 519690 81096 524400 81152
rect 519629 81094 524400 81096
rect 519629 81091 519695 81094
rect 523200 81064 524400 81094
rect 115933 79930 115999 79933
rect 521101 79930 521167 79933
rect 115933 79928 119140 79930
rect 115933 79872 115938 79928
rect 115994 79872 119140 79928
rect 115933 79870 119140 79872
rect 518788 79928 521167 79930
rect 518788 79872 521106 79928
rect 521162 79872 521167 79928
rect 518788 79870 521167 79872
rect 115933 79867 115999 79870
rect 521101 79867 521167 79870
rect 520181 79658 520247 79661
rect 523200 79658 524400 79688
rect 520181 79656 524400 79658
rect 520181 79600 520186 79656
rect 520242 79600 524400 79656
rect 520181 79598 524400 79600
rect 520181 79595 520247 79598
rect 523200 79568 524400 79598
rect 520273 78570 520339 78573
rect 518788 78568 520339 78570
rect 518788 78512 520278 78568
rect 520334 78512 520339 78568
rect 518788 78510 520339 78512
rect 520273 78507 520339 78510
rect 520089 78162 520155 78165
rect 523200 78162 524400 78192
rect 520089 78160 524400 78162
rect 520089 78104 520094 78160
rect 520150 78104 524400 78160
rect 520089 78102 524400 78104
rect 520089 78099 520155 78102
rect 523200 78072 524400 78102
rect 116117 78026 116183 78029
rect 116117 78024 119140 78026
rect 116117 77968 116122 78024
rect 116178 77968 119140 78024
rect 116117 77966 119140 77968
rect 116117 77963 116183 77966
rect 520917 77210 520983 77213
rect 518788 77208 520983 77210
rect 518788 77152 520922 77208
rect 520978 77152 520983 77208
rect 518788 77150 520983 77152
rect 520917 77147 520983 77150
rect 519997 76666 520063 76669
rect 523200 76666 524400 76696
rect 519997 76664 524400 76666
rect 519997 76608 520002 76664
rect 520058 76608 524400 76664
rect 519997 76606 524400 76608
rect 519997 76603 520063 76606
rect 523200 76576 524400 76606
rect 519905 75986 519971 75989
rect 110860 75926 119140 75986
rect 518788 75984 519971 75986
rect 518788 75928 519910 75984
rect 519966 75928 519971 75984
rect 518788 75926 519971 75928
rect 519905 75923 519971 75926
rect 519905 75170 519971 75173
rect 523200 75170 524400 75200
rect 519905 75168 524400 75170
rect 519905 75112 519910 75168
rect 519966 75112 524400 75168
rect 519905 75110 524400 75112
rect 519905 75107 519971 75110
rect 523200 75080 524400 75110
rect 519629 74626 519695 74629
rect 518788 74624 519695 74626
rect 518788 74568 519634 74624
rect 519690 74568 519695 74624
rect 518788 74566 519695 74568
rect 519629 74563 519695 74566
rect 116669 74082 116735 74085
rect 116669 74080 119140 74082
rect 116669 74024 116674 74080
rect 116730 74024 119140 74080
rect 116669 74022 119140 74024
rect 116669 74019 116735 74022
rect 519261 73674 519327 73677
rect 523200 73674 524400 73704
rect 519261 73672 524400 73674
rect 519261 73616 519266 73672
rect 519322 73616 524400 73672
rect 519261 73614 524400 73616
rect 519261 73611 519327 73614
rect 523200 73584 524400 73614
rect 520181 73266 520247 73269
rect 518788 73264 520247 73266
rect 518788 73208 520186 73264
rect 520242 73208 520247 73264
rect 518788 73206 520247 73208
rect 520181 73203 520247 73206
rect 520089 72450 520155 72453
rect 518758 72448 520155 72450
rect 518758 72392 520094 72448
rect 520150 72392 520155 72448
rect 518758 72390 520155 72392
rect 116577 72178 116643 72181
rect 116577 72176 119140 72178
rect 116577 72120 116582 72176
rect 116638 72120 119140 72176
rect 116577 72118 119140 72120
rect 116577 72115 116643 72118
rect 518758 71876 518818 72390
rect 520089 72387 520155 72390
rect 520181 72042 520247 72045
rect 523200 72042 524400 72072
rect 520181 72040 524400 72042
rect 520181 71984 520186 72040
rect 520242 71984 524400 72040
rect 520181 71982 524400 71984
rect 520181 71979 520247 71982
rect 523200 71952 524400 71982
rect 519997 70546 520063 70549
rect 523200 70546 524400 70576
rect 518788 70544 520063 70546
rect 518788 70488 520002 70544
rect 520058 70488 520063 70544
rect 518788 70486 520063 70488
rect 519997 70483 520063 70486
rect 520230 70486 524400 70546
rect 520089 70410 520155 70413
rect 520230 70410 520290 70486
rect 523200 70456 524400 70486
rect 520089 70408 520290 70410
rect 520089 70352 520094 70408
rect 520150 70352 520290 70408
rect 520089 70350 520290 70352
rect 520089 70347 520155 70350
rect 116301 70274 116367 70277
rect 116301 70272 119140 70274
rect 116301 70216 116306 70272
rect 116362 70216 119140 70272
rect 116301 70214 119140 70216
rect 116301 70211 116367 70214
rect 519905 69186 519971 69189
rect 518788 69184 519971 69186
rect 518788 69128 519910 69184
rect 519966 69128 519971 69184
rect 518788 69126 519971 69128
rect 519905 69123 519971 69126
rect 519629 69050 519695 69053
rect 523200 69050 524400 69080
rect 519629 69048 524400 69050
rect 519629 68992 519634 69048
rect 519690 68992 524400 69048
rect 519629 68990 524400 68992
rect 519629 68987 519695 68990
rect 523200 68960 524400 68990
rect 116117 68370 116183 68373
rect 116117 68368 119140 68370
rect 116117 68312 116122 68368
rect 116178 68312 119140 68368
rect 116117 68310 119140 68312
rect 116117 68307 116183 68310
rect 519261 67826 519327 67829
rect 518788 67824 519327 67826
rect 518788 67768 519266 67824
rect 519322 67768 519327 67824
rect 518788 67766 519327 67768
rect 519261 67763 519327 67766
rect 520457 67554 520523 67557
rect 523200 67554 524400 67584
rect 520457 67552 524400 67554
rect 520457 67496 520462 67552
rect 520518 67496 524400 67552
rect 520457 67494 524400 67496
rect 520457 67491 520523 67494
rect 523200 67464 524400 67494
rect 116577 66466 116643 66469
rect 520181 66466 520247 66469
rect 116577 66464 119140 66466
rect 116577 66408 116582 66464
rect 116638 66408 119140 66464
rect 116577 66406 119140 66408
rect 518788 66464 520247 66466
rect 518788 66408 520186 66464
rect 520242 66408 520247 66464
rect 518788 66406 520247 66408
rect 116577 66403 116643 66406
rect 520181 66403 520247 66406
rect 520365 66058 520431 66061
rect 523200 66058 524400 66088
rect 520365 66056 524400 66058
rect 520365 66000 520370 66056
rect 520426 66000 524400 66056
rect 520365 65998 524400 66000
rect 520365 65995 520431 65998
rect 523200 65968 524400 65998
rect 520089 65106 520155 65109
rect 518788 65104 520155 65106
rect 518788 65048 520094 65104
rect 520150 65048 520155 65104
rect 518788 65046 520155 65048
rect 520089 65043 520155 65046
rect 113357 64562 113423 64565
rect 110860 64560 113423 64562
rect 110860 64504 113362 64560
rect 113418 64504 113423 64560
rect 110860 64502 113423 64504
rect 113357 64499 113423 64502
rect 116209 64562 116275 64565
rect 521101 64562 521167 64565
rect 523200 64562 524400 64592
rect 116209 64560 119140 64562
rect 116209 64504 116214 64560
rect 116270 64504 119140 64560
rect 116209 64502 119140 64504
rect 521101 64560 524400 64562
rect 521101 64504 521106 64560
rect 521162 64504 524400 64560
rect 521101 64502 524400 64504
rect 116209 64499 116275 64502
rect 521101 64499 521167 64502
rect 523200 64472 524400 64502
rect 519629 63746 519695 63749
rect 518788 63744 519695 63746
rect 518788 63688 519634 63744
rect 519690 63688 519695 63744
rect 518788 63686 519695 63688
rect 519629 63683 519695 63686
rect 521193 62930 521259 62933
rect 523200 62930 524400 62960
rect 521193 62928 524400 62930
rect 521193 62872 521198 62928
rect 521254 62872 524400 62928
rect 521193 62870 524400 62872
rect 521193 62867 521259 62870
rect 523200 62840 524400 62870
rect 116117 62658 116183 62661
rect 116117 62656 119140 62658
rect 116117 62600 116122 62656
rect 116178 62600 119140 62656
rect 116117 62598 119140 62600
rect 116117 62595 116183 62598
rect 520457 62386 520523 62389
rect 518788 62384 520523 62386
rect 518788 62328 520462 62384
rect 520518 62328 520523 62384
rect 518788 62326 520523 62328
rect 520457 62323 520523 62326
rect 520273 61434 520339 61437
rect 523200 61434 524400 61464
rect 520273 61432 524400 61434
rect 520273 61376 520278 61432
rect 520334 61376 524400 61432
rect 520273 61374 524400 61376
rect 520273 61371 520339 61374
rect 523200 61344 524400 61374
rect 520365 61026 520431 61029
rect 518788 61024 520431 61026
rect 518788 60968 520370 61024
rect 520426 60968 520431 61024
rect 518788 60966 520431 60968
rect 520365 60963 520431 60966
rect 116577 60618 116643 60621
rect 116577 60616 119140 60618
rect 116577 60560 116582 60616
rect 116638 60560 119140 60616
rect 116577 60558 119140 60560
rect 116577 60555 116643 60558
rect 521009 59938 521075 59941
rect 523200 59938 524400 59968
rect 521009 59936 524400 59938
rect 521009 59880 521014 59936
rect 521070 59880 524400 59936
rect 521009 59878 524400 59880
rect 521009 59875 521075 59878
rect 523200 59848 524400 59878
rect 521101 59666 521167 59669
rect 518788 59664 521167 59666
rect 518788 59608 521106 59664
rect 521162 59608 521167 59664
rect 518788 59606 521167 59608
rect 521101 59603 521167 59606
rect 116669 58714 116735 58717
rect 116669 58712 119140 58714
rect 116669 58656 116674 58712
rect 116730 58656 119140 58712
rect 116669 58654 119140 58656
rect 116669 58651 116735 58654
rect 521101 58442 521167 58445
rect 523200 58442 524400 58472
rect 521101 58440 524400 58442
rect 521101 58384 521106 58440
rect 521162 58384 524400 58440
rect 521101 58382 524400 58384
rect 521101 58379 521167 58382
rect 523200 58352 524400 58382
rect 521193 58306 521259 58309
rect 518788 58304 521259 58306
rect 518788 58248 521198 58304
rect 521254 58248 521259 58304
rect 518788 58246 521259 58248
rect 521193 58243 521259 58246
rect 520181 56946 520247 56949
rect 518788 56944 520247 56946
rect 518788 56888 520186 56944
rect 520242 56888 520247 56944
rect 518788 56886 520247 56888
rect 520181 56883 520247 56886
rect 520365 56946 520431 56949
rect 523200 56946 524400 56976
rect 520365 56944 524400 56946
rect 520365 56888 520370 56944
rect 520426 56888 524400 56944
rect 520365 56886 524400 56888
rect 520365 56883 520431 56886
rect 523200 56856 524400 56886
rect 116761 56810 116827 56813
rect 116761 56808 119140 56810
rect 116761 56752 116766 56808
rect 116822 56752 119140 56808
rect 116761 56750 119140 56752
rect 116761 56747 116827 56750
rect 521009 55586 521075 55589
rect 518788 55584 521075 55586
rect 518788 55528 521014 55584
rect 521070 55528 521075 55584
rect 518788 55526 521075 55528
rect 521009 55523 521075 55526
rect 520273 55450 520339 55453
rect 523200 55450 524400 55480
rect 520273 55448 524400 55450
rect 520273 55392 520278 55448
rect 520334 55392 524400 55448
rect 520273 55390 524400 55392
rect 520273 55387 520339 55390
rect 523200 55360 524400 55390
rect 110321 53954 110387 53957
rect 119110 53954 119170 54876
rect 521101 54226 521167 54229
rect 518788 54224 521167 54226
rect 518788 54168 521106 54224
rect 521162 54168 521167 54224
rect 518788 54166 521167 54168
rect 521101 54163 521167 54166
rect 110321 53952 119170 53954
rect 110321 53896 110326 53952
rect 110382 53896 119170 53952
rect 110321 53894 119170 53896
rect 110321 53891 110387 53894
rect 519261 53818 519327 53821
rect 523200 53818 524400 53848
rect 519261 53816 524400 53818
rect 519261 53760 519266 53816
rect 519322 53760 524400 53816
rect 519261 53758 524400 53760
rect 519261 53755 519327 53758
rect 523200 53728 524400 53758
rect 114185 53138 114251 53141
rect 110860 53136 114251 53138
rect 110860 53080 114190 53136
rect 114246 53080 114251 53136
rect 110860 53078 114251 53080
rect 114185 53075 114251 53078
rect 110321 52594 110387 52597
rect 119110 52594 119170 52972
rect 520365 52866 520431 52869
rect 518788 52864 520431 52866
rect 518788 52808 520370 52864
rect 520426 52808 520431 52864
rect 518788 52806 520431 52808
rect 520365 52803 520431 52806
rect 110321 52592 119170 52594
rect 110321 52536 110326 52592
rect 110382 52536 119170 52592
rect 110321 52534 119170 52536
rect 110321 52531 110387 52534
rect 520089 52322 520155 52325
rect 523200 52322 524400 52352
rect 520089 52320 524400 52322
rect 520089 52264 520094 52320
rect 520150 52264 524400 52320
rect 520089 52262 524400 52264
rect 520089 52259 520155 52262
rect 523200 52232 524400 52262
rect 520273 51506 520339 51509
rect 518788 51504 520339 51506
rect 518788 51448 520278 51504
rect 520334 51448 520339 51504
rect 518788 51446 520339 51448
rect 520273 51443 520339 51446
rect 110321 51098 110387 51101
rect 110321 51096 119140 51098
rect 110321 51040 110326 51096
rect 110382 51040 119140 51096
rect 110321 51038 119140 51040
rect 110321 51035 110387 51038
rect 519997 50826 520063 50829
rect 523200 50826 524400 50856
rect 519997 50824 524400 50826
rect 519997 50768 520002 50824
rect 520058 50768 524400 50824
rect 519997 50766 524400 50768
rect 519997 50763 520063 50766
rect 523200 50736 524400 50766
rect 519261 50146 519327 50149
rect 518788 50144 519327 50146
rect 518788 50088 519266 50144
rect 519322 50088 519327 50144
rect 518788 50086 519327 50088
rect 519261 50083 519327 50086
rect 520181 49330 520247 49333
rect 523200 49330 524400 49360
rect 520181 49328 524400 49330
rect 520181 49272 520186 49328
rect 520242 49272 524400 49328
rect 520181 49270 524400 49272
rect 520181 49267 520247 49270
rect 523200 49240 524400 49270
rect 110321 48378 110387 48381
rect 119110 48378 119170 49164
rect 520089 48786 520155 48789
rect 518788 48784 520155 48786
rect 518788 48728 520094 48784
rect 520150 48728 520155 48784
rect 518788 48726 520155 48728
rect 520089 48723 520155 48726
rect 110321 48376 119170 48378
rect 110321 48320 110326 48376
rect 110382 48320 119170 48376
rect 110321 48318 119170 48320
rect 110321 48315 110387 48318
rect 519445 47834 519511 47837
rect 523200 47834 524400 47864
rect 519445 47832 524400 47834
rect 519445 47776 519450 47832
rect 519506 47776 524400 47832
rect 519445 47774 524400 47776
rect 519445 47771 519511 47774
rect 523200 47744 524400 47774
rect 519997 47426 520063 47429
rect 518788 47424 520063 47426
rect 518788 47368 520002 47424
rect 520058 47368 520063 47424
rect 518788 47366 520063 47368
rect 519997 47363 520063 47366
rect 110321 47154 110387 47157
rect 110321 47152 119140 47154
rect 110321 47096 110326 47152
rect 110382 47096 119140 47152
rect 110321 47094 119140 47096
rect 110321 47091 110387 47094
rect 519905 46338 519971 46341
rect 523200 46338 524400 46368
rect 519905 46336 524400 46338
rect 519905 46280 519910 46336
rect 519966 46280 524400 46336
rect 519905 46278 524400 46280
rect 519905 46275 519971 46278
rect 523200 46248 524400 46278
rect 520181 46066 520247 46069
rect 518788 46064 520247 46066
rect 518788 46008 520186 46064
rect 520242 46008 520247 46064
rect 518788 46006 520247 46008
rect 520181 46003 520247 46006
rect 110321 44298 110387 44301
rect 119110 44298 119170 45220
rect 519445 44706 519511 44709
rect 518788 44704 519511 44706
rect 518788 44648 519450 44704
rect 519506 44648 519511 44704
rect 518788 44646 519511 44648
rect 519445 44643 519511 44646
rect 519813 44706 519879 44709
rect 523200 44706 524400 44736
rect 519813 44704 524400 44706
rect 519813 44648 519818 44704
rect 519874 44648 524400 44704
rect 519813 44646 524400 44648
rect 519813 44643 519879 44646
rect 523200 44616 524400 44646
rect 110321 44296 119170 44298
rect 110321 44240 110326 44296
rect 110382 44240 119170 44296
rect 110321 44238 119170 44240
rect 110321 44235 110387 44238
rect 116117 43346 116183 43349
rect 519905 43346 519971 43349
rect 116117 43344 119140 43346
rect 116117 43288 116122 43344
rect 116178 43288 119140 43344
rect 116117 43286 119140 43288
rect 518788 43344 519971 43346
rect 518788 43288 519910 43344
rect 519966 43288 519971 43344
rect 518788 43286 519971 43288
rect 116117 43283 116183 43286
rect 519905 43283 519971 43286
rect 520181 43210 520247 43213
rect 523200 43210 524400 43240
rect 520181 43208 524400 43210
rect 520181 43152 520186 43208
rect 520242 43152 524400 43208
rect 520181 43150 524400 43152
rect 520181 43147 520247 43150
rect 523200 43120 524400 43150
rect 519813 41986 519879 41989
rect 518788 41984 519879 41986
rect 518788 41928 519818 41984
rect 519874 41928 519879 41984
rect 518788 41926 519879 41928
rect 519813 41923 519879 41926
rect 114093 41850 114159 41853
rect 110860 41848 114159 41850
rect 110860 41792 114098 41848
rect 114154 41792 114159 41848
rect 110860 41790 114159 41792
rect 114093 41787 114159 41790
rect 520089 41714 520155 41717
rect 523200 41714 524400 41744
rect 520089 41712 524400 41714
rect 520089 41656 520094 41712
rect 520150 41656 524400 41712
rect 520089 41654 524400 41656
rect 520089 41651 520155 41654
rect 523200 41624 524400 41654
rect 110321 41442 110387 41445
rect 110321 41440 119140 41442
rect 110321 41384 110326 41440
rect 110382 41384 119140 41440
rect 110321 41382 119140 41384
rect 110321 41379 110387 41382
rect 520181 40626 520247 40629
rect 518788 40624 520247 40626
rect 518788 40568 520186 40624
rect 520242 40568 520247 40624
rect 518788 40566 520247 40568
rect 520181 40563 520247 40566
rect 520181 40218 520247 40221
rect 523200 40218 524400 40248
rect 520181 40216 524400 40218
rect 520181 40160 520186 40216
rect 520242 40160 524400 40216
rect 520181 40158 524400 40160
rect 520181 40155 520247 40158
rect 523200 40128 524400 40158
rect 116945 39538 117011 39541
rect 116945 39536 119140 39538
rect 116945 39480 116950 39536
rect 117006 39480 119140 39536
rect 116945 39478 119140 39480
rect 116945 39475 117011 39478
rect 520089 39266 520155 39269
rect 518788 39264 520155 39266
rect 518788 39208 520094 39264
rect 520150 39208 520155 39264
rect 518788 39206 520155 39208
rect 520089 39203 520155 39206
rect 519813 38722 519879 38725
rect 523200 38722 524400 38752
rect 519813 38720 524400 38722
rect 519813 38664 519818 38720
rect 519874 38664 524400 38720
rect 519813 38662 524400 38664
rect 519813 38659 519879 38662
rect 523200 38632 524400 38662
rect 520181 37906 520247 37909
rect 518788 37904 520247 37906
rect 518788 37848 520186 37904
rect 520242 37848 520247 37904
rect 518788 37846 520247 37848
rect 520181 37843 520247 37846
rect 116853 37634 116919 37637
rect 116853 37632 119140 37634
rect 116853 37576 116858 37632
rect 116914 37576 119140 37632
rect 116853 37574 119140 37576
rect 116853 37571 116919 37574
rect 521561 37226 521627 37229
rect 523200 37226 524400 37256
rect 521561 37224 524400 37226
rect 521561 37168 521566 37224
rect 521622 37168 524400 37224
rect 521561 37166 524400 37168
rect 521561 37163 521627 37166
rect 523200 37136 524400 37166
rect 519813 36546 519879 36549
rect 518788 36544 519879 36546
rect 518788 36488 519818 36544
rect 519874 36488 519879 36544
rect 518788 36486 519879 36488
rect 519813 36483 519879 36486
rect 521561 36002 521627 36005
rect 521561 36000 521670 36002
rect 521561 35944 521566 36000
rect 521622 35944 521670 36000
rect 521561 35939 521670 35944
rect 521610 35866 521670 35939
rect 518758 35806 521670 35866
rect 110321 34642 110387 34645
rect 119110 34642 119170 35700
rect 518758 35156 518818 35806
rect 521101 35594 521167 35597
rect 523200 35594 524400 35624
rect 521101 35592 524400 35594
rect 521101 35536 521106 35592
rect 521162 35536 524400 35592
rect 521101 35534 524400 35536
rect 521101 35531 521167 35534
rect 523200 35504 524400 35534
rect 110321 34640 119170 34642
rect 110321 34584 110326 34640
rect 110382 34584 119170 34640
rect 110321 34582 119170 34584
rect 110321 34579 110387 34582
rect 521101 34506 521167 34509
rect 518758 34504 521167 34506
rect 518758 34448 521106 34504
rect 521162 34448 521167 34504
rect 518758 34446 521167 34448
rect 117129 33826 117195 33829
rect 117129 33824 119140 33826
rect 117129 33768 117134 33824
rect 117190 33768 119140 33824
rect 518758 33796 518818 34446
rect 521101 34443 521167 34446
rect 520917 34098 520983 34101
rect 523200 34098 524400 34128
rect 520917 34096 524400 34098
rect 520917 34040 520922 34096
rect 520978 34040 524400 34096
rect 520917 34038 524400 34040
rect 520917 34035 520983 34038
rect 523200 34008 524400 34038
rect 117129 33766 119140 33768
rect 117129 33763 117195 33766
rect 520917 33146 520983 33149
rect 518758 33144 520983 33146
rect 518758 33088 520922 33144
rect 520978 33088 520983 33144
rect 518758 33086 520983 33088
rect 518758 32436 518818 33086
rect 520917 33083 520983 33086
rect 520917 32602 520983 32605
rect 523200 32602 524400 32632
rect 520917 32600 524400 32602
rect 520917 32544 520922 32600
rect 520978 32544 524400 32600
rect 520917 32542 524400 32544
rect 520917 32539 520983 32542
rect 523200 32512 524400 32542
rect 117037 31786 117103 31789
rect 117037 31784 119140 31786
rect 117037 31728 117042 31784
rect 117098 31728 119140 31784
rect 117037 31726 119140 31728
rect 117037 31723 117103 31726
rect 520917 31650 520983 31653
rect 518758 31648 520983 31650
rect 518758 31592 520922 31648
rect 520978 31592 520983 31648
rect 518758 31590 520983 31592
rect 518758 31076 518818 31590
rect 520917 31587 520983 31590
rect 520917 31106 520983 31109
rect 523200 31106 524400 31136
rect 520917 31104 524400 31106
rect 520917 31048 520922 31104
rect 520978 31048 524400 31104
rect 520917 31046 524400 31048
rect 520917 31043 520983 31046
rect 523200 31016 524400 31046
rect 114001 30426 114067 30429
rect 110860 30424 114067 30426
rect 110860 30368 114006 30424
rect 114062 30368 114067 30424
rect 110860 30366 114067 30368
rect 114001 30363 114067 30366
rect 520917 30290 520983 30293
rect 518758 30288 520983 30290
rect 518758 30232 520922 30288
rect 520978 30232 520983 30288
rect 518758 30230 520983 30232
rect 117221 29882 117287 29885
rect 117221 29880 119140 29882
rect 117221 29824 117226 29880
rect 117282 29824 119140 29880
rect 117221 29822 119140 29824
rect 117221 29819 117287 29822
rect 518758 29716 518818 30230
rect 520917 30227 520983 30230
rect 521101 29610 521167 29613
rect 523200 29610 524400 29640
rect 521101 29608 524400 29610
rect 521101 29552 521106 29608
rect 521162 29552 524400 29608
rect 521101 29550 524400 29552
rect 521101 29547 521167 29550
rect 523200 29520 524400 29550
rect 521101 28386 521167 28389
rect 518788 28384 521167 28386
rect 518788 28328 521106 28384
rect 521162 28328 521167 28384
rect 518788 28326 521167 28328
rect 521101 28323 521167 28326
rect 523200 28114 524400 28144
rect 518850 28054 524400 28114
rect 116485 27978 116551 27981
rect 116485 27976 119140 27978
rect 116485 27920 116490 27976
rect 116546 27920 119140 27976
rect 116485 27918 119140 27920
rect 116485 27915 116551 27918
rect 518850 27570 518910 28054
rect 523200 28024 524400 28054
rect 518758 27510 518910 27570
rect 518758 26996 518818 27510
rect 523200 26482 524400 26512
rect 521610 26422 524400 26482
rect 521610 26210 521670 26422
rect 523200 26392 524400 26422
rect 518758 26150 521670 26210
rect 116301 26074 116367 26077
rect 116301 26072 119140 26074
rect 116301 26016 116306 26072
rect 116362 26016 119140 26072
rect 116301 26014 119140 26016
rect 116301 26011 116367 26014
rect 518758 25636 518818 26150
rect 523200 24986 524400 25016
rect 518850 24926 524400 24986
rect 518850 24850 518910 24926
rect 523200 24896 524400 24926
rect 518758 24790 518910 24850
rect 518758 24276 518818 24790
rect 116393 24170 116459 24173
rect 116393 24168 119140 24170
rect 116393 24112 116398 24168
rect 116454 24112 119140 24168
rect 116393 24110 119140 24112
rect 116393 24107 116459 24110
rect 523200 23490 524400 23520
rect 518758 23430 524400 23490
rect 518758 22916 518818 23430
rect 523200 23400 524400 23430
rect 116209 22266 116275 22269
rect 116209 22264 119140 22266
rect 116209 22208 116214 22264
rect 116270 22208 119140 22264
rect 116209 22206 119140 22208
rect 116209 22203 116275 22206
rect 521101 21994 521167 21997
rect 523200 21994 524400 22024
rect 521101 21992 524400 21994
rect 521101 21936 521106 21992
rect 521162 21936 524400 21992
rect 521101 21934 524400 21936
rect 521101 21931 521167 21934
rect 523200 21904 524400 21934
rect 518758 20906 518818 21556
rect 521101 20906 521167 20909
rect 518758 20904 521167 20906
rect 518758 20848 521106 20904
rect 521162 20848 521167 20904
rect 518758 20846 521167 20848
rect 521101 20843 521167 20846
rect 520733 20498 520799 20501
rect 523200 20498 524400 20528
rect 520733 20496 524400 20498
rect 520733 20440 520738 20496
rect 520794 20440 524400 20496
rect 520733 20438 524400 20440
rect 520733 20435 520799 20438
rect 523200 20408 524400 20438
rect 116025 20362 116091 20365
rect 116025 20360 119140 20362
rect 116025 20304 116030 20360
rect 116086 20304 119140 20360
rect 116025 20302 119140 20304
rect 116025 20299 116091 20302
rect 518758 19546 518818 20196
rect 520733 19546 520799 19549
rect 518758 19544 520799 19546
rect 518758 19488 520738 19544
rect 520794 19488 520799 19544
rect 518758 19486 520799 19488
rect 520733 19483 520799 19486
rect 113909 19002 113975 19005
rect 110860 19000 113975 19002
rect 110860 18944 113914 19000
rect 113970 18944 113975 19000
rect 110860 18942 113975 18944
rect 113909 18939 113975 18942
rect 520917 19002 520983 19005
rect 523200 19002 524400 19032
rect 520917 19000 524400 19002
rect 520917 18944 520922 19000
rect 520978 18944 524400 19000
rect 520917 18942 524400 18944
rect 520917 18939 520983 18942
rect 523200 18912 524400 18942
rect 116117 18458 116183 18461
rect 116117 18456 119140 18458
rect 116117 18400 116122 18456
rect 116178 18400 119140 18456
rect 116117 18398 119140 18400
rect 116117 18395 116183 18398
rect 518758 18186 518818 18836
rect 520917 18186 520983 18189
rect 518758 18184 520983 18186
rect 518758 18128 520922 18184
rect 520978 18128 520983 18184
rect 518758 18126 520983 18128
rect 520917 18123 520983 18126
rect 518758 16826 518818 17476
rect 523200 17370 524400 17400
rect 521150 17310 524400 17370
rect 521150 16826 521210 17310
rect 523200 17280 524400 17310
rect 518758 16766 521210 16826
rect 115933 16418 115999 16421
rect 115933 16416 119140 16418
rect 115933 16360 115938 16416
rect 115994 16360 119140 16416
rect 115933 16358 119140 16360
rect 115933 16355 115999 16358
rect 518758 15466 518818 16116
rect 523200 15874 524400 15904
rect 521104 15814 524400 15874
rect 521104 15466 521164 15814
rect 523200 15784 524400 15814
rect 518758 15406 521164 15466
rect 116526 14452 116532 14516
rect 116596 14514 116602 14516
rect 116596 14454 119140 14514
rect 116596 14452 116602 14454
rect 518758 14106 518818 14756
rect 523200 14378 524400 14408
rect 521104 14318 524400 14378
rect 521104 14106 521164 14318
rect 523200 14288 524400 14318
rect 518758 14046 521164 14106
rect 518758 12746 518818 13396
rect 523200 12882 524400 12912
rect 521104 12822 524400 12882
rect 521104 12746 521164 12822
rect 523200 12792 524400 12822
rect 518758 12686 521164 12746
rect 116710 12548 116716 12612
rect 116780 12610 116786 12612
rect 116780 12550 119140 12610
rect 116780 12548 116786 12550
rect 518758 11386 518818 12036
rect 523200 11386 524400 11416
rect 518758 11326 524400 11386
rect 523200 11296 524400 11326
rect 116894 10644 116900 10708
rect 116964 10706 116970 10708
rect 116964 10646 119140 10706
rect 116964 10644 116970 10646
rect 518758 10026 518818 10676
rect 518758 9966 518910 10026
rect 518850 9890 518910 9966
rect 523200 9890 524400 9920
rect 518850 9830 524400 9890
rect 523200 9800 524400 9830
rect 521101 9346 521167 9349
rect 518788 9344 521167 9346
rect 518788 9288 521106 9344
rect 521162 9288 521167 9344
rect 518788 9286 521167 9288
rect 521101 9283 521167 9286
rect 117262 8740 117268 8804
rect 117332 8802 117338 8804
rect 117332 8742 119140 8802
rect 117332 8740 117338 8742
rect 110321 8394 110387 8397
rect 110321 8392 110522 8394
rect 110321 8336 110326 8392
rect 110382 8336 110522 8392
rect 110321 8334 110522 8336
rect 110321 8331 110387 8334
rect 110462 8258 110522 8334
rect 110597 8258 110663 8261
rect 110462 8256 110663 8258
rect 110462 8200 110602 8256
rect 110658 8200 110663 8256
rect 110462 8198 110663 8200
rect 110597 8195 110663 8198
rect 521101 8258 521167 8261
rect 523200 8258 524400 8288
rect 521101 8256 524400 8258
rect 521101 8200 521106 8256
rect 521162 8200 524400 8256
rect 521101 8198 524400 8200
rect 521101 8195 521167 8198
rect 523200 8168 524400 8198
rect 110321 8122 110387 8125
rect 110505 8122 110571 8125
rect 110321 8120 110571 8122
rect 110321 8064 110326 8120
rect 110382 8064 110510 8120
rect 110566 8064 110571 8120
rect 110321 8062 110571 8064
rect 110321 8059 110387 8062
rect 110505 8059 110571 8062
rect 520365 7986 520431 7989
rect 518788 7984 520431 7986
rect 518788 7928 520370 7984
rect 520426 7928 520431 7984
rect 518788 7926 520431 7928
rect 520365 7923 520431 7926
rect 113817 7714 113883 7717
rect 110860 7712 113883 7714
rect 110860 7656 113822 7712
rect 113878 7656 113883 7712
rect 110860 7654 113883 7656
rect 113817 7651 113883 7654
rect 111057 7034 111123 7037
rect 116761 7034 116827 7037
rect 111057 7032 116827 7034
rect 111057 6976 111062 7032
rect 111118 6976 116766 7032
rect 116822 6976 116827 7032
rect 111057 6974 116827 6976
rect 111057 6971 111123 6974
rect 116761 6971 116827 6974
rect 117129 6898 117195 6901
rect 117129 6896 119140 6898
rect 117129 6840 117134 6896
rect 117190 6840 119140 6896
rect 117129 6838 119140 6840
rect 117129 6835 117195 6838
rect 520365 6762 520431 6765
rect 523200 6762 524400 6792
rect 520365 6760 524400 6762
rect 520365 6704 520370 6760
rect 520426 6704 524400 6760
rect 520365 6702 524400 6704
rect 520365 6699 520431 6702
rect 523200 6672 524400 6702
rect 521101 6626 521167 6629
rect 518788 6624 521167 6626
rect 518788 6568 521106 6624
rect 521162 6568 521167 6624
rect 518788 6566 521167 6568
rect 521101 6563 521167 6566
rect 110505 5674 110571 5677
rect 115841 5674 115907 5677
rect 110505 5672 115907 5674
rect 110505 5616 110510 5672
rect 110566 5616 115846 5672
rect 115902 5616 115907 5672
rect 110505 5614 115907 5616
rect 110505 5611 110571 5614
rect 115841 5611 115907 5614
rect 520917 5266 520983 5269
rect 518788 5264 520983 5266
rect 518788 5208 520922 5264
rect 520978 5208 520983 5264
rect 518788 5206 520983 5208
rect 520917 5203 520983 5206
rect 521101 5266 521167 5269
rect 523200 5266 524400 5296
rect 521101 5264 524400 5266
rect 521101 5208 521106 5264
rect 521162 5208 524400 5264
rect 521101 5206 524400 5208
rect 521101 5203 521167 5206
rect 523200 5176 524400 5206
rect 119110 4178 119170 4964
rect 110462 4118 119170 4178
rect 68694 3982 83658 4042
rect 55170 3438 59370 3498
rect 55170 3090 55230 3438
rect 45510 3030 55230 3090
rect 45510 2818 45570 3030
rect 32446 2758 45570 2818
rect 59310 2818 59370 3438
rect 59310 2758 63234 2818
rect 32446 2685 32506 2758
rect 32397 2680 32506 2685
rect 32397 2624 32402 2680
rect 32458 2624 32506 2680
rect 32397 2622 32506 2624
rect 36353 2682 36419 2685
rect 62389 2682 62455 2685
rect 36353 2680 62455 2682
rect 36353 2624 36358 2680
rect 36414 2624 62394 2680
rect 62450 2624 62455 2680
rect 36353 2622 62455 2624
rect 63174 2682 63234 2758
rect 64137 2682 64203 2685
rect 63174 2680 64203 2682
rect 63174 2624 64142 2680
rect 64198 2624 64203 2680
rect 63174 2622 64203 2624
rect 32397 2619 32463 2622
rect 36353 2619 36419 2622
rect 62389 2619 62455 2622
rect 64137 2619 64203 2622
rect 65333 2682 65399 2685
rect 68001 2682 68067 2685
rect 65333 2680 68067 2682
rect 65333 2624 65338 2680
rect 65394 2624 68006 2680
rect 68062 2624 68067 2680
rect 65333 2622 68067 2624
rect 65333 2619 65399 2622
rect 68001 2619 68067 2622
rect 68553 2682 68619 2685
rect 68694 2682 68754 3982
rect 83598 3498 83658 3982
rect 88290 3982 89730 4042
rect 83598 3438 83842 3498
rect 83782 3226 83842 3438
rect 88290 3226 88350 3982
rect 89670 3498 89730 3982
rect 91050 3982 92490 4042
rect 91050 3770 91110 3982
rect 90958 3710 91110 3770
rect 90958 3498 91018 3710
rect 92430 3634 92490 3982
rect 93810 3982 95250 4042
rect 93810 3770 93870 3982
rect 93350 3710 93870 3770
rect 93350 3634 93410 3710
rect 92430 3574 93410 3634
rect 89670 3438 91018 3498
rect 95190 3362 95250 3982
rect 99330 3982 109786 4042
rect 96570 3846 98010 3906
rect 96570 3362 96630 3846
rect 95190 3302 96630 3362
rect 83598 3166 83842 3226
rect 84150 3166 88350 3226
rect 83598 2954 83658 3166
rect 84150 2954 84210 3166
rect 92430 3030 93870 3090
rect 83598 2894 88350 2954
rect 84150 2818 84210 2894
rect 68832 2758 77954 2818
rect 68832 2685 68892 2758
rect 77894 2685 77954 2758
rect 78124 2758 84210 2818
rect 88290 2818 88350 2894
rect 89670 2894 91110 2954
rect 89670 2818 89730 2894
rect 88290 2758 89730 2818
rect 91050 2818 91110 2894
rect 92430 2818 92490 3030
rect 91050 2758 92490 2818
rect 93810 2818 93870 3030
rect 95190 3030 96630 3090
rect 95190 2818 95250 3030
rect 93810 2758 95250 2818
rect 96570 2818 96630 3030
rect 97950 2954 98010 3846
rect 99330 2954 99390 3982
rect 109726 3770 109786 3982
rect 110229 3906 110295 3909
rect 110462 3906 110522 4118
rect 521009 3906 521075 3909
rect 110229 3904 110522 3906
rect 110229 3848 110234 3904
rect 110290 3848 110522 3904
rect 110229 3846 110522 3848
rect 518788 3904 521075 3906
rect 518788 3848 521014 3904
rect 521070 3848 521075 3904
rect 518788 3846 521075 3848
rect 110229 3843 110295 3846
rect 521009 3843 521075 3846
rect 520917 3770 520983 3773
rect 523200 3770 524400 3800
rect 109726 3710 113190 3770
rect 109493 3634 109559 3637
rect 109677 3634 109743 3637
rect 109493 3632 109743 3634
rect 109493 3576 109498 3632
rect 109554 3576 109682 3632
rect 109738 3576 109743 3632
rect 109493 3574 109743 3576
rect 109493 3571 109559 3574
rect 109677 3571 109743 3574
rect 109861 3634 109927 3637
rect 110045 3634 110111 3637
rect 109861 3632 110111 3634
rect 109861 3576 109866 3632
rect 109922 3576 110050 3632
rect 110106 3576 110111 3632
rect 109861 3574 110111 3576
rect 113130 3634 113190 3710
rect 520917 3768 524400 3770
rect 520917 3712 520922 3768
rect 520978 3712 524400 3768
rect 520917 3710 524400 3712
rect 520917 3707 520983 3710
rect 523200 3680 524400 3710
rect 116301 3634 116367 3637
rect 113130 3632 116367 3634
rect 113130 3576 116306 3632
rect 116362 3576 116367 3632
rect 113130 3574 116367 3576
rect 109861 3571 109927 3574
rect 110045 3571 110111 3574
rect 116301 3571 116367 3574
rect 109493 3498 109559 3501
rect 110229 3498 110295 3501
rect 109493 3496 110295 3498
rect 109493 3440 109498 3496
rect 109554 3440 110234 3496
rect 110290 3440 110295 3496
rect 109493 3438 110295 3440
rect 109493 3435 109559 3438
rect 110229 3435 110295 3438
rect 116945 3362 117011 3365
rect 97950 2894 99390 2954
rect 102090 3360 117011 3362
rect 102090 3304 116950 3360
rect 117006 3304 117011 3360
rect 102090 3302 117011 3304
rect 102090 2818 102150 3302
rect 116945 3299 117011 3302
rect 110597 3226 110663 3229
rect 117037 3226 117103 3229
rect 104206 3224 110663 3226
rect 104206 3168 110602 3224
rect 110658 3168 110663 3224
rect 104206 3166 110663 3168
rect 104206 3090 104266 3166
rect 110597 3163 110663 3166
rect 113038 3224 117103 3226
rect 113038 3168 117042 3224
rect 117098 3168 117103 3224
rect 113038 3166 117103 3168
rect 113038 3090 113098 3166
rect 117037 3163 117103 3166
rect 96570 2758 102150 2818
rect 103838 3030 104266 3090
rect 104942 3030 113098 3090
rect 116301 3090 116367 3093
rect 116301 3088 119140 3090
rect 116301 3032 116306 3088
rect 116362 3032 119140 3088
rect 116301 3030 119140 3032
rect 78124 2685 78184 2758
rect 68553 2680 68754 2682
rect 68553 2624 68558 2680
rect 68614 2624 68754 2680
rect 68553 2622 68754 2624
rect 68829 2680 68895 2685
rect 68829 2624 68834 2680
rect 68890 2624 68895 2680
rect 68553 2619 68619 2622
rect 68829 2619 68895 2624
rect 69381 2682 69447 2685
rect 77017 2682 77083 2685
rect 69381 2680 77083 2682
rect 69381 2624 69386 2680
rect 69442 2624 77022 2680
rect 77078 2624 77083 2680
rect 69381 2622 77083 2624
rect 69381 2619 69447 2622
rect 77017 2619 77083 2622
rect 77247 2682 77313 2685
rect 77753 2682 77819 2685
rect 77247 2680 77819 2682
rect 77247 2624 77252 2680
rect 77308 2624 77758 2680
rect 77814 2624 77819 2680
rect 77247 2622 77819 2624
rect 77894 2680 78003 2685
rect 77894 2624 77942 2680
rect 77998 2624 78003 2680
rect 77894 2622 78003 2624
rect 77247 2619 77313 2622
rect 77753 2619 77819 2622
rect 77937 2619 78003 2622
rect 78121 2680 78187 2685
rect 78121 2624 78126 2680
rect 78182 2624 78187 2680
rect 78121 2619 78187 2624
rect 78305 2682 78371 2685
rect 95693 2682 95759 2685
rect 78305 2680 95759 2682
rect 78305 2624 78310 2680
rect 78366 2624 95698 2680
rect 95754 2624 95759 2680
rect 78305 2622 95759 2624
rect 78305 2619 78371 2622
rect 95693 2619 95759 2622
rect 96337 2682 96403 2685
rect 103697 2682 103763 2685
rect 96337 2680 103763 2682
rect 96337 2624 96342 2680
rect 96398 2624 103702 2680
rect 103758 2624 103763 2680
rect 96337 2622 103763 2624
rect 96337 2619 96403 2622
rect 103697 2619 103763 2622
rect 33041 2546 33107 2549
rect 96613 2546 96679 2549
rect 33041 2544 96679 2546
rect 33041 2488 33046 2544
rect 33102 2488 96618 2544
rect 96674 2488 96679 2544
rect 33041 2486 96679 2488
rect 33041 2483 33107 2486
rect 96613 2483 96679 2486
rect 97257 2546 97323 2549
rect 103838 2546 103898 3030
rect 104341 2682 104407 2685
rect 104942 2682 105002 3030
rect 116301 3027 116367 3030
rect 111701 2954 111767 2957
rect 105310 2952 111767 2954
rect 105310 2896 111706 2952
rect 111762 2896 111767 2952
rect 105310 2894 111767 2896
rect 104341 2680 105002 2682
rect 104341 2624 104346 2680
rect 104402 2624 105002 2680
rect 104341 2622 105002 2624
rect 105077 2682 105143 2685
rect 105310 2682 105370 2894
rect 111701 2891 111767 2894
rect 109401 2818 109467 2821
rect 106414 2816 109467 2818
rect 106414 2760 109406 2816
rect 109462 2760 109467 2816
rect 106414 2758 109467 2760
rect 105077 2680 105370 2682
rect 105077 2624 105082 2680
rect 105138 2624 105370 2680
rect 105077 2622 105370 2624
rect 106273 2682 106339 2685
rect 106414 2682 106474 2758
rect 109401 2755 109467 2758
rect 109861 2818 109927 2821
rect 110505 2818 110571 2821
rect 109861 2816 110571 2818
rect 109861 2760 109866 2816
rect 109922 2760 110510 2816
rect 110566 2760 110571 2816
rect 109861 2758 110571 2760
rect 109861 2755 109927 2758
rect 110505 2755 110571 2758
rect 106273 2680 106474 2682
rect 106273 2624 106278 2680
rect 106334 2624 106474 2680
rect 106273 2622 106474 2624
rect 107607 2682 107673 2685
rect 116209 2682 116275 2685
rect 521101 2682 521167 2685
rect 107607 2680 116275 2682
rect 107607 2624 107612 2680
rect 107668 2624 116214 2680
rect 116270 2624 116275 2680
rect 107607 2622 116275 2624
rect 518788 2680 521167 2682
rect 518788 2624 521106 2680
rect 521162 2624 521167 2680
rect 518788 2622 521167 2624
rect 104341 2619 104407 2622
rect 105077 2619 105143 2622
rect 106273 2619 106339 2622
rect 107607 2619 107673 2622
rect 116209 2619 116275 2622
rect 521101 2619 521167 2622
rect 107193 2546 107259 2549
rect 97257 2544 103898 2546
rect 97257 2488 97262 2544
rect 97318 2488 103898 2544
rect 97257 2486 103898 2488
rect 104206 2544 107259 2546
rect 104206 2488 107198 2544
rect 107254 2488 107259 2544
rect 104206 2486 107259 2488
rect 97257 2483 97323 2486
rect 29545 2410 29611 2413
rect 104206 2410 104266 2486
rect 107193 2483 107259 2486
rect 107561 2546 107627 2549
rect 116025 2546 116091 2549
rect 107561 2544 116091 2546
rect 107561 2488 107566 2544
rect 107622 2488 116030 2544
rect 116086 2488 116091 2544
rect 107561 2486 116091 2488
rect 107561 2483 107627 2486
rect 116025 2483 116091 2486
rect 29545 2408 104266 2410
rect 29545 2352 29550 2408
rect 29606 2352 104266 2408
rect 29545 2350 104266 2352
rect 106457 2410 106523 2413
rect 107285 2410 107351 2413
rect 106457 2408 107351 2410
rect 106457 2352 106462 2408
rect 106518 2352 107290 2408
rect 107346 2352 107351 2408
rect 106457 2350 107351 2352
rect 29545 2347 29611 2350
rect 106457 2347 106523 2350
rect 107285 2347 107351 2350
rect 107607 2410 107673 2413
rect 116117 2410 116183 2413
rect 107607 2408 116183 2410
rect 107607 2352 107612 2408
rect 107668 2352 116122 2408
rect 116178 2352 116183 2408
rect 107607 2350 116183 2352
rect 107607 2347 107673 2350
rect 116117 2347 116183 2350
rect 26049 2274 26115 2277
rect 106825 2274 106891 2277
rect 26049 2272 106891 2274
rect 26049 2216 26054 2272
rect 26110 2216 106830 2272
rect 106886 2216 106891 2272
rect 26049 2214 106891 2216
rect 26049 2211 26115 2214
rect 106825 2211 106891 2214
rect 107009 2274 107075 2277
rect 115933 2274 115999 2277
rect 107009 2272 115999 2274
rect 107009 2216 107014 2272
rect 107070 2216 115938 2272
rect 115994 2216 115999 2272
rect 107009 2214 115999 2216
rect 107009 2211 107075 2214
rect 115933 2211 115999 2214
rect 521009 2274 521075 2277
rect 523200 2274 524400 2304
rect 521009 2272 524400 2274
rect 521009 2216 521014 2272
rect 521070 2216 524400 2272
rect 521009 2214 524400 2216
rect 521009 2211 521075 2214
rect 523200 2184 524400 2214
rect 22921 2138 22987 2141
rect 94865 2138 94931 2141
rect 22921 2136 94931 2138
rect 22921 2080 22926 2136
rect 22982 2080 94870 2136
rect 94926 2080 94931 2136
rect 22921 2078 94931 2080
rect 22921 2075 22987 2078
rect 94865 2075 94931 2078
rect 95693 2138 95759 2141
rect 97257 2138 97323 2141
rect 95693 2136 97323 2138
rect 95693 2080 95698 2136
rect 95754 2080 97262 2136
rect 97318 2080 97323 2136
rect 95693 2078 97323 2080
rect 95693 2075 95759 2078
rect 97257 2075 97323 2078
rect 100845 2138 100911 2141
rect 107285 2138 107351 2141
rect 100845 2136 107351 2138
rect 100845 2080 100850 2136
rect 100906 2080 107290 2136
rect 107346 2080 107351 2136
rect 100845 2078 107351 2080
rect 100845 2075 100911 2078
rect 107285 2075 107351 2078
rect 107561 2138 107627 2141
rect 116526 2138 116532 2140
rect 107561 2136 116532 2138
rect 107561 2080 107566 2136
rect 107622 2080 116532 2136
rect 107561 2078 116532 2080
rect 107561 2075 107627 2078
rect 116526 2076 116532 2078
rect 116596 2076 116602 2140
rect 19609 2002 19675 2005
rect 107101 2002 107167 2005
rect 19609 2000 107167 2002
rect 19609 1944 19614 2000
rect 19670 1944 107106 2000
rect 107162 1944 107167 2000
rect 19609 1942 107167 1944
rect 19609 1939 19675 1942
rect 107101 1939 107167 1942
rect 107561 2002 107627 2005
rect 116710 2002 116716 2004
rect 107561 2000 116716 2002
rect 107561 1944 107566 2000
rect 107622 1944 116716 2000
rect 107561 1942 116716 1944
rect 107561 1939 107627 1942
rect 116710 1940 116716 1942
rect 116780 1940 116786 2004
rect 15929 1866 15995 1869
rect 106774 1866 106780 1868
rect 15929 1864 106780 1866
rect 15929 1808 15934 1864
rect 15990 1808 106780 1864
rect 15929 1806 106780 1808
rect 15929 1803 15995 1806
rect 106774 1804 106780 1806
rect 106844 1804 106850 1868
rect 107602 1804 107608 1868
rect 107672 1866 107678 1868
rect 116894 1866 116900 1868
rect 107672 1806 116900 1866
rect 107672 1804 107678 1806
rect 116894 1804 116900 1806
rect 116964 1804 116970 1868
rect 5993 1730 6059 1733
rect 109493 1730 109559 1733
rect 5993 1728 109559 1730
rect 5993 1672 5998 1728
rect 6054 1672 109498 1728
rect 109554 1672 109559 1728
rect 5993 1670 109559 1672
rect 5993 1667 6059 1670
rect 109493 1667 109559 1670
rect 12617 1594 12683 1597
rect 117262 1594 117268 1596
rect 12617 1592 117268 1594
rect 12617 1536 12622 1592
rect 12678 1536 117268 1592
rect 12617 1534 117268 1536
rect 12617 1531 12683 1534
rect 117262 1532 117268 1534
rect 117332 1532 117338 1596
rect 229277 1594 229343 1597
rect 293585 1594 293651 1597
rect 229277 1592 293651 1594
rect 229277 1536 229282 1592
rect 229338 1536 293590 1592
rect 293646 1536 293651 1592
rect 229277 1534 293651 1536
rect 229277 1531 229343 1534
rect 293585 1531 293651 1534
rect 9305 1458 9371 1461
rect 117129 1458 117195 1461
rect 9305 1456 117195 1458
rect 9305 1400 9310 1456
rect 9366 1400 117134 1456
rect 117190 1400 117195 1456
rect 9305 1398 117195 1400
rect 9305 1395 9371 1398
rect 117129 1395 117195 1398
rect 163773 1458 163839 1461
rect 243629 1458 243695 1461
rect 163773 1456 243695 1458
rect 163773 1400 163778 1456
rect 163834 1400 243634 1456
rect 243690 1400 243695 1456
rect 163773 1398 243695 1400
rect 163773 1395 163839 1398
rect 243629 1395 243695 1398
rect 360285 1458 360351 1461
rect 393589 1458 393655 1461
rect 360285 1456 393655 1458
rect 360285 1400 360290 1456
rect 360346 1400 393594 1456
rect 393650 1400 393655 1456
rect 360285 1398 393655 1400
rect 360285 1395 360351 1398
rect 393589 1395 393655 1398
rect 85941 1322 86007 1325
rect 103973 1322 104039 1325
rect 85941 1320 104039 1322
rect 85941 1264 85946 1320
rect 86002 1264 103978 1320
rect 104034 1264 104039 1320
rect 85941 1262 104039 1264
rect 85941 1259 86007 1262
rect 103973 1259 104039 1262
rect 104157 1322 104223 1325
rect 110321 1322 110387 1325
rect 104157 1320 110387 1322
rect 104157 1264 104162 1320
rect 104218 1264 110326 1320
rect 110382 1264 110387 1320
rect 104157 1262 110387 1264
rect 104157 1259 104223 1262
rect 110321 1259 110387 1262
rect 88333 1186 88399 1189
rect 101029 1186 101095 1189
rect 104341 1186 104407 1189
rect 88333 1184 100770 1186
rect 88333 1128 88338 1184
rect 88394 1128 100770 1184
rect 88333 1126 100770 1128
rect 88333 1123 88399 1126
rect 100710 1050 100770 1126
rect 101029 1184 104407 1186
rect 101029 1128 101034 1184
rect 101090 1128 104346 1184
rect 104402 1128 104407 1184
rect 101029 1126 104407 1128
rect 101029 1123 101095 1126
rect 104341 1123 104407 1126
rect 107009 1050 107075 1053
rect 100710 1048 107075 1050
rect 100710 992 107014 1048
rect 107070 992 107075 1048
rect 100710 990 107075 992
rect 107009 987 107075 990
rect 96613 914 96679 917
rect 106457 914 106523 917
rect 96613 912 106523 914
rect 96613 856 96618 912
rect 96674 856 106462 912
rect 106518 856 106523 912
rect 96613 854 106523 856
rect 96613 851 96679 854
rect 106457 851 106523 854
rect 521101 778 521167 781
rect 523200 778 524400 808
rect 521101 776 524400 778
rect 521101 720 521106 776
rect 521162 720 524400 776
rect 521101 718 524400 720
rect 521101 715 521167 718
rect 523200 688 524400 718
<< via3 >>
rect 116532 14452 116596 14516
rect 116716 12548 116780 12612
rect 116900 10644 116964 10708
rect 117268 8740 117332 8804
rect 116532 2076 116596 2140
rect 116716 1940 116780 2004
rect 106780 1804 106844 1868
rect 107608 1804 107672 1868
rect 116900 1804 116964 1868
rect 117268 1532 117332 1596
<< metal4 >>
rect 1664 144454 1984 144496
rect 1664 144218 1706 144454
rect 1942 144218 1984 144454
rect 1664 144134 1984 144218
rect 1664 143898 1706 144134
rect 1942 143898 1984 144134
rect 1664 143856 1984 143898
rect 109956 144454 110276 144496
rect 109956 144218 109998 144454
rect 110234 144218 110276 144454
rect 109956 144134 110276 144218
rect 109956 143898 109998 144134
rect 110234 143898 110276 144134
rect 109956 143856 110276 143898
rect 119664 144454 119984 144496
rect 119664 144218 119706 144454
rect 119942 144218 119984 144454
rect 119664 144134 119984 144218
rect 119664 143898 119706 144134
rect 119942 143898 119984 144134
rect 119664 143856 119984 143898
rect 517940 144454 518260 144496
rect 517940 144218 517982 144454
rect 518218 144218 518260 144454
rect 517940 144134 518260 144218
rect 517940 143898 517982 144134
rect 518218 143898 518260 144134
rect 517940 143856 518260 143898
rect 1096 131454 1332 131496
rect 1096 131134 1332 131218
rect 1096 130856 1332 130898
rect 110616 131454 110936 131496
rect 110616 131218 110658 131454
rect 110894 131218 110936 131454
rect 110616 131134 110936 131218
rect 110616 130898 110658 131134
rect 110894 130898 110936 131134
rect 110616 130856 110936 130898
rect 119004 131454 119324 131496
rect 119004 131218 119046 131454
rect 119282 131218 119324 131454
rect 119004 131134 119324 131218
rect 119004 130898 119046 131134
rect 119282 130898 119324 131134
rect 119004 130856 119324 130898
rect 518600 131454 518920 131496
rect 518600 131218 518642 131454
rect 518878 131218 518920 131454
rect 518600 131134 518920 131218
rect 518600 130898 518642 131134
rect 518878 130898 518920 131134
rect 518600 130856 518920 130898
rect 1664 118454 1984 118496
rect 1664 118218 1706 118454
rect 1942 118218 1984 118454
rect 1664 118134 1984 118218
rect 1664 117898 1706 118134
rect 1942 117898 1984 118134
rect 1664 117856 1984 117898
rect 109956 118454 110276 118496
rect 109956 118218 109998 118454
rect 110234 118218 110276 118454
rect 109956 118134 110276 118218
rect 109956 117898 109998 118134
rect 110234 117898 110276 118134
rect 109956 117856 110276 117898
rect 119664 118454 119984 118496
rect 119664 118218 119706 118454
rect 119942 118218 119984 118454
rect 119664 118134 119984 118218
rect 119664 117898 119706 118134
rect 119942 117898 119984 118134
rect 119664 117856 119984 117898
rect 517940 118454 518260 118496
rect 517940 118218 517982 118454
rect 518218 118218 518260 118454
rect 517940 118134 518260 118218
rect 517940 117898 517982 118134
rect 518218 117898 518260 118134
rect 517940 117856 518260 117898
rect 1096 105454 1332 105496
rect 1096 105134 1332 105218
rect 1096 104856 1332 104898
rect 110616 105454 110936 105496
rect 110616 105218 110658 105454
rect 110894 105218 110936 105454
rect 110616 105134 110936 105218
rect 110616 104898 110658 105134
rect 110894 104898 110936 105134
rect 110616 104856 110936 104898
rect 119004 105454 119324 105496
rect 119004 105218 119046 105454
rect 119282 105218 119324 105454
rect 119004 105134 119324 105218
rect 119004 104898 119046 105134
rect 119282 104898 119324 105134
rect 119004 104856 119324 104898
rect 518600 105454 518920 105496
rect 518600 105218 518642 105454
rect 518878 105218 518920 105454
rect 518600 105134 518920 105218
rect 518600 104898 518642 105134
rect 518878 104898 518920 105134
rect 518600 104856 518920 104898
rect 1664 92454 1984 92496
rect 1664 92218 1706 92454
rect 1942 92218 1984 92454
rect 1664 92134 1984 92218
rect 1664 91898 1706 92134
rect 1942 91898 1984 92134
rect 1664 91856 1984 91898
rect 109956 92454 110276 92496
rect 109956 92218 109998 92454
rect 110234 92218 110276 92454
rect 109956 92134 110276 92218
rect 109956 91898 109998 92134
rect 110234 91898 110276 92134
rect 109956 91856 110276 91898
rect 119664 92454 119984 92496
rect 119664 92218 119706 92454
rect 119942 92218 119984 92454
rect 119664 92134 119984 92218
rect 119664 91898 119706 92134
rect 119942 91898 119984 92134
rect 119664 91856 119984 91898
rect 517940 92454 518260 92496
rect 517940 92218 517982 92454
rect 518218 92218 518260 92454
rect 517940 92134 518260 92218
rect 517940 91898 517982 92134
rect 518218 91898 518260 92134
rect 517940 91856 518260 91898
rect 1096 79454 1332 79496
rect 1096 79134 1332 79218
rect 1096 78856 1332 78898
rect 110616 79454 110936 79496
rect 110616 79218 110658 79454
rect 110894 79218 110936 79454
rect 110616 79134 110936 79218
rect 110616 78898 110658 79134
rect 110894 78898 110936 79134
rect 110616 78856 110936 78898
rect 119004 79454 119324 79496
rect 119004 79218 119046 79454
rect 119282 79218 119324 79454
rect 119004 79134 119324 79218
rect 119004 78898 119046 79134
rect 119282 78898 119324 79134
rect 119004 78856 119324 78898
rect 518600 79454 518920 79496
rect 518600 79218 518642 79454
rect 518878 79218 518920 79454
rect 518600 79134 518920 79218
rect 518600 78898 518642 79134
rect 518878 78898 518920 79134
rect 518600 78856 518920 78898
rect 1664 66454 1984 66496
rect 1664 66218 1706 66454
rect 1942 66218 1984 66454
rect 1664 66134 1984 66218
rect 1664 65898 1706 66134
rect 1942 65898 1984 66134
rect 1664 65856 1984 65898
rect 109956 66454 110276 66496
rect 109956 66218 109998 66454
rect 110234 66218 110276 66454
rect 109956 66134 110276 66218
rect 109956 65898 109998 66134
rect 110234 65898 110276 66134
rect 109956 65856 110276 65898
rect 119664 66454 119984 66496
rect 119664 66218 119706 66454
rect 119942 66218 119984 66454
rect 119664 66134 119984 66218
rect 119664 65898 119706 66134
rect 119942 65898 119984 66134
rect 119664 65856 119984 65898
rect 517940 66454 518260 66496
rect 517940 66218 517982 66454
rect 518218 66218 518260 66454
rect 517940 66134 518260 66218
rect 517940 65898 517982 66134
rect 518218 65898 518260 66134
rect 517940 65856 518260 65898
rect 1096 53454 1332 53496
rect 1096 53134 1332 53218
rect 1096 52856 1332 52898
rect 110616 53454 110936 53496
rect 110616 53218 110658 53454
rect 110894 53218 110936 53454
rect 110616 53134 110936 53218
rect 110616 52898 110658 53134
rect 110894 52898 110936 53134
rect 110616 52856 110936 52898
rect 119004 53454 119324 53496
rect 119004 53218 119046 53454
rect 119282 53218 119324 53454
rect 119004 53134 119324 53218
rect 119004 52898 119046 53134
rect 119282 52898 119324 53134
rect 119004 52856 119324 52898
rect 518600 53454 518920 53496
rect 518600 53218 518642 53454
rect 518878 53218 518920 53454
rect 518600 53134 518920 53218
rect 518600 52898 518642 53134
rect 518878 52898 518920 53134
rect 518600 52856 518920 52898
rect 1664 40454 1984 40496
rect 1664 40218 1706 40454
rect 1942 40218 1984 40454
rect 1664 40134 1984 40218
rect 1664 39898 1706 40134
rect 1942 39898 1984 40134
rect 1664 39856 1984 39898
rect 109956 40454 110276 40496
rect 109956 40218 109998 40454
rect 110234 40218 110276 40454
rect 109956 40134 110276 40218
rect 109956 39898 109998 40134
rect 110234 39898 110276 40134
rect 109956 39856 110276 39898
rect 119664 40454 119984 40496
rect 119664 40218 119706 40454
rect 119942 40218 119984 40454
rect 119664 40134 119984 40218
rect 119664 39898 119706 40134
rect 119942 39898 119984 40134
rect 119664 39856 119984 39898
rect 517940 40454 518260 40496
rect 517940 40218 517982 40454
rect 518218 40218 518260 40454
rect 517940 40134 518260 40218
rect 517940 39898 517982 40134
rect 518218 39898 518260 40134
rect 517940 39856 518260 39898
rect 1096 27454 1332 27496
rect 1096 27134 1332 27218
rect 1096 26856 1332 26898
rect 110616 27454 110936 27496
rect 110616 27218 110658 27454
rect 110894 27218 110936 27454
rect 110616 27134 110936 27218
rect 110616 26898 110658 27134
rect 110894 26898 110936 27134
rect 110616 26856 110936 26898
rect 119004 27454 119324 27496
rect 119004 27218 119046 27454
rect 119282 27218 119324 27454
rect 119004 27134 119324 27218
rect 119004 26898 119046 27134
rect 119282 26898 119324 27134
rect 119004 26856 119324 26898
rect 518600 27454 518920 27496
rect 518600 27218 518642 27454
rect 518878 27218 518920 27454
rect 518600 27134 518920 27218
rect 518600 26898 518642 27134
rect 518878 26898 518920 27134
rect 518600 26856 518920 26898
rect 116531 14516 116597 14517
rect 1664 14454 1984 14496
rect 1664 14218 1706 14454
rect 1942 14218 1984 14454
rect 1664 14134 1984 14218
rect 1664 13898 1706 14134
rect 1942 13898 1984 14134
rect 1664 13856 1984 13898
rect 109956 14454 110276 14496
rect 109956 14218 109998 14454
rect 110234 14218 110276 14454
rect 116531 14452 116532 14516
rect 116596 14452 116597 14516
rect 116531 14451 116597 14452
rect 119664 14454 119984 14496
rect 109956 14134 110276 14218
rect 109956 13898 109998 14134
rect 110234 13898 110276 14134
rect 109956 13856 110276 13898
rect 116534 2141 116594 14451
rect 119664 14218 119706 14454
rect 119942 14218 119984 14454
rect 119664 14134 119984 14218
rect 119664 13898 119706 14134
rect 119942 13898 119984 14134
rect 119664 13856 119984 13898
rect 517940 14454 518260 14496
rect 517940 14218 517982 14454
rect 518218 14218 518260 14454
rect 517940 14134 518260 14218
rect 517940 13898 517982 14134
rect 518218 13898 518260 14134
rect 517940 13856 518260 13898
rect 116715 12612 116781 12613
rect 116715 12548 116716 12612
rect 116780 12548 116781 12612
rect 116715 12547 116781 12548
rect 116531 2140 116597 2141
rect 116531 2076 116532 2140
rect 116596 2076 116597 2140
rect 116531 2075 116597 2076
rect 116718 2005 116778 12547
rect 116899 10708 116965 10709
rect 116899 10644 116900 10708
rect 116964 10644 116965 10708
rect 116899 10643 116965 10644
rect 116715 2004 116781 2005
rect 116715 1940 116716 2004
rect 116780 1940 116781 2004
rect 116715 1939 116781 1940
rect 116902 1869 116962 10643
rect 117267 8804 117333 8805
rect 117267 8740 117268 8804
rect 117332 8740 117333 8804
rect 117267 8739 117333 8740
rect 106779 1868 106845 1869
rect 106779 1804 106780 1868
rect 106844 1804 106845 1868
rect 106779 1803 106845 1804
rect 107607 1868 107673 1869
rect 107607 1804 107608 1868
rect 107672 1804 107673 1868
rect 107607 1803 107673 1804
rect 116899 1868 116965 1869
rect 116899 1804 116900 1868
rect 116964 1804 116965 1868
rect 116899 1803 116965 1804
rect 106782 1730 106842 1803
rect 107610 1730 107670 1803
rect 106782 1670 107670 1730
rect 117270 1597 117330 8739
rect 117267 1596 117333 1597
rect 117267 1532 117268 1596
rect 117332 1532 117333 1596
rect 117267 1531 117333 1532
<< via4 >>
rect 1706 144218 1942 144454
rect 1706 143898 1942 144134
rect 109998 144218 110234 144454
rect 109998 143898 110234 144134
rect 119706 144218 119942 144454
rect 119706 143898 119942 144134
rect 517982 144218 518218 144454
rect 517982 143898 518218 144134
rect 1096 131218 1332 131454
rect 1096 130898 1332 131134
rect 110658 131218 110894 131454
rect 110658 130898 110894 131134
rect 119046 131218 119282 131454
rect 119046 130898 119282 131134
rect 518642 131218 518878 131454
rect 518642 130898 518878 131134
rect 1706 118218 1942 118454
rect 1706 117898 1942 118134
rect 109998 118218 110234 118454
rect 109998 117898 110234 118134
rect 119706 118218 119942 118454
rect 119706 117898 119942 118134
rect 517982 118218 518218 118454
rect 517982 117898 518218 118134
rect 1096 105218 1332 105454
rect 1096 104898 1332 105134
rect 110658 105218 110894 105454
rect 110658 104898 110894 105134
rect 119046 105218 119282 105454
rect 119046 104898 119282 105134
rect 518642 105218 518878 105454
rect 518642 104898 518878 105134
rect 1706 92218 1942 92454
rect 1706 91898 1942 92134
rect 109998 92218 110234 92454
rect 109998 91898 110234 92134
rect 119706 92218 119942 92454
rect 119706 91898 119942 92134
rect 517982 92218 518218 92454
rect 517982 91898 518218 92134
rect 1096 79218 1332 79454
rect 1096 78898 1332 79134
rect 110658 79218 110894 79454
rect 110658 78898 110894 79134
rect 119046 79218 119282 79454
rect 119046 78898 119282 79134
rect 518642 79218 518878 79454
rect 518642 78898 518878 79134
rect 1706 66218 1942 66454
rect 1706 65898 1942 66134
rect 109998 66218 110234 66454
rect 109998 65898 110234 66134
rect 119706 66218 119942 66454
rect 119706 65898 119942 66134
rect 517982 66218 518218 66454
rect 517982 65898 518218 66134
rect 1096 53218 1332 53454
rect 1096 52898 1332 53134
rect 110658 53218 110894 53454
rect 110658 52898 110894 53134
rect 119046 53218 119282 53454
rect 119046 52898 119282 53134
rect 518642 53218 518878 53454
rect 518642 52898 518878 53134
rect 1706 40218 1942 40454
rect 1706 39898 1942 40134
rect 109998 40218 110234 40454
rect 109998 39898 110234 40134
rect 119706 40218 119942 40454
rect 119706 39898 119942 40134
rect 517982 40218 518218 40454
rect 517982 39898 518218 40134
rect 1096 27218 1332 27454
rect 1096 26898 1332 27134
rect 110658 27218 110894 27454
rect 110658 26898 110894 27134
rect 119046 27218 119282 27454
rect 119046 26898 119282 27134
rect 518642 27218 518878 27454
rect 518642 26898 518878 27134
rect 1706 14218 1942 14454
rect 1706 13898 1942 14134
rect 109998 14218 110234 14454
rect 109998 13898 110234 14134
rect 119706 14218 119942 14454
rect 119706 13898 119942 14134
rect 517982 14218 518218 14454
rect 517982 13898 518218 14134
<< metal5 >>
rect 1104 156856 522836 157496
rect 1104 144454 2200 144496
rect 1104 144218 1706 144454
rect 1942 144218 2200 144454
rect 1104 144134 2200 144218
rect 1104 143898 1706 144134
rect 1942 143898 2200 144134
rect 1104 143856 2200 143898
rect 109800 144454 120200 144496
rect 109800 144218 109998 144454
rect 110234 144218 119706 144454
rect 119942 144218 120200 144454
rect 109800 144134 120200 144218
rect 109800 143898 109998 144134
rect 110234 143898 119706 144134
rect 119942 143898 120200 144134
rect 109800 143856 120200 143898
rect 517800 144454 522836 144496
rect 517800 144218 517982 144454
rect 518218 144218 522836 144454
rect 517800 144134 522836 144218
rect 517800 143898 517982 144134
rect 518218 143898 522836 144134
rect 517800 143856 522836 143898
rect 1072 131454 2200 131496
rect 1072 131218 1096 131454
rect 1332 131218 2200 131454
rect 1072 131134 2200 131218
rect 1072 130898 1096 131134
rect 1332 130898 2200 131134
rect 1072 130856 2200 130898
rect 109800 131454 120200 131496
rect 109800 131218 110658 131454
rect 110894 131218 119046 131454
rect 119282 131218 120200 131454
rect 109800 131134 120200 131218
rect 109800 130898 110658 131134
rect 110894 130898 119046 131134
rect 119282 130898 120200 131134
rect 109800 130856 120200 130898
rect 517800 131454 522836 131496
rect 517800 131218 518642 131454
rect 518878 131218 522836 131454
rect 517800 131134 522836 131218
rect 517800 130898 518642 131134
rect 518878 130898 522836 131134
rect 517800 130856 522836 130898
rect 1104 118454 2200 118496
rect 1104 118218 1706 118454
rect 1942 118218 2200 118454
rect 1104 118134 2200 118218
rect 1104 117898 1706 118134
rect 1942 117898 2200 118134
rect 1104 117856 2200 117898
rect 109800 118454 120200 118496
rect 109800 118218 109998 118454
rect 110234 118218 119706 118454
rect 119942 118218 120200 118454
rect 109800 118134 120200 118218
rect 109800 117898 109998 118134
rect 110234 117898 119706 118134
rect 119942 117898 120200 118134
rect 109800 117856 120200 117898
rect 517800 118454 522836 118496
rect 517800 118218 517982 118454
rect 518218 118218 522836 118454
rect 517800 118134 522836 118218
rect 517800 117898 517982 118134
rect 518218 117898 522836 118134
rect 517800 117856 522836 117898
rect 1072 105454 2200 105496
rect 1072 105218 1096 105454
rect 1332 105218 2200 105454
rect 1072 105134 2200 105218
rect 1072 104898 1096 105134
rect 1332 104898 2200 105134
rect 1072 104856 2200 104898
rect 109800 105454 120200 105496
rect 109800 105218 110658 105454
rect 110894 105218 119046 105454
rect 119282 105218 120200 105454
rect 109800 105134 120200 105218
rect 109800 104898 110658 105134
rect 110894 104898 119046 105134
rect 119282 104898 120200 105134
rect 109800 104856 120200 104898
rect 517800 105454 522836 105496
rect 517800 105218 518642 105454
rect 518878 105218 522836 105454
rect 517800 105134 522836 105218
rect 517800 104898 518642 105134
rect 518878 104898 522836 105134
rect 517800 104856 522836 104898
rect 1104 92454 2200 92496
rect 1104 92218 1706 92454
rect 1942 92218 2200 92454
rect 1104 92134 2200 92218
rect 1104 91898 1706 92134
rect 1942 91898 2200 92134
rect 1104 91856 2200 91898
rect 109800 92454 120200 92496
rect 109800 92218 109998 92454
rect 110234 92218 119706 92454
rect 119942 92218 120200 92454
rect 109800 92134 120200 92218
rect 109800 91898 109998 92134
rect 110234 91898 119706 92134
rect 119942 91898 120200 92134
rect 109800 91856 120200 91898
rect 517800 92454 522836 92496
rect 517800 92218 517982 92454
rect 518218 92218 522836 92454
rect 517800 92134 522836 92218
rect 517800 91898 517982 92134
rect 518218 91898 522836 92134
rect 517800 91856 522836 91898
rect 1072 79454 2200 79496
rect 1072 79218 1096 79454
rect 1332 79218 2200 79454
rect 1072 79134 2200 79218
rect 1072 78898 1096 79134
rect 1332 78898 2200 79134
rect 1072 78856 2200 78898
rect 109800 79454 120200 79496
rect 109800 79218 110658 79454
rect 110894 79218 119046 79454
rect 119282 79218 120200 79454
rect 109800 79134 120200 79218
rect 109800 78898 110658 79134
rect 110894 78898 119046 79134
rect 119282 78898 120200 79134
rect 109800 78856 120200 78898
rect 517800 79454 522836 79496
rect 517800 79218 518642 79454
rect 518878 79218 522836 79454
rect 517800 79134 522836 79218
rect 517800 78898 518642 79134
rect 518878 78898 522836 79134
rect 517800 78856 522836 78898
rect 1104 66454 2200 66496
rect 1104 66218 1706 66454
rect 1942 66218 2200 66454
rect 1104 66134 2200 66218
rect 1104 65898 1706 66134
rect 1942 65898 2200 66134
rect 1104 65856 2200 65898
rect 109800 66454 120200 66496
rect 109800 66218 109998 66454
rect 110234 66218 119706 66454
rect 119942 66218 120200 66454
rect 109800 66134 120200 66218
rect 109800 65898 109998 66134
rect 110234 65898 119706 66134
rect 119942 65898 120200 66134
rect 109800 65856 120200 65898
rect 517800 66454 522836 66496
rect 517800 66218 517982 66454
rect 518218 66218 522836 66454
rect 517800 66134 522836 66218
rect 517800 65898 517982 66134
rect 518218 65898 522836 66134
rect 517800 65856 522836 65898
rect 1072 53454 2200 53496
rect 1072 53218 1096 53454
rect 1332 53218 2200 53454
rect 1072 53134 2200 53218
rect 1072 52898 1096 53134
rect 1332 52898 2200 53134
rect 1072 52856 2200 52898
rect 109800 53454 120200 53496
rect 109800 53218 110658 53454
rect 110894 53218 119046 53454
rect 119282 53218 120200 53454
rect 109800 53134 120200 53218
rect 109800 52898 110658 53134
rect 110894 52898 119046 53134
rect 119282 52898 120200 53134
rect 109800 52856 120200 52898
rect 517800 53454 522836 53496
rect 517800 53218 518642 53454
rect 518878 53218 522836 53454
rect 517800 53134 522836 53218
rect 517800 52898 518642 53134
rect 518878 52898 522836 53134
rect 517800 52856 522836 52898
rect 1104 40454 2200 40496
rect 1104 40218 1706 40454
rect 1942 40218 2200 40454
rect 1104 40134 2200 40218
rect 1104 39898 1706 40134
rect 1942 39898 2200 40134
rect 1104 39856 2200 39898
rect 109800 40454 120200 40496
rect 109800 40218 109998 40454
rect 110234 40218 119706 40454
rect 119942 40218 120200 40454
rect 109800 40134 120200 40218
rect 109800 39898 109998 40134
rect 110234 39898 119706 40134
rect 119942 39898 120200 40134
rect 109800 39856 120200 39898
rect 517800 40454 522836 40496
rect 517800 40218 517982 40454
rect 518218 40218 522836 40454
rect 517800 40134 522836 40218
rect 517800 39898 517982 40134
rect 518218 39898 522836 40134
rect 517800 39856 522836 39898
rect 1072 27454 2200 27496
rect 1072 27218 1096 27454
rect 1332 27218 2200 27454
rect 1072 27134 2200 27218
rect 1072 26898 1096 27134
rect 1332 26898 2200 27134
rect 1072 26856 2200 26898
rect 109800 27454 120200 27496
rect 109800 27218 110658 27454
rect 110894 27218 119046 27454
rect 119282 27218 120200 27454
rect 109800 27134 120200 27218
rect 109800 26898 110658 27134
rect 110894 26898 119046 27134
rect 119282 26898 120200 27134
rect 109800 26856 120200 26898
rect 517800 27454 522836 27496
rect 517800 27218 518642 27454
rect 518878 27218 522836 27454
rect 517800 27134 522836 27218
rect 517800 26898 518642 27134
rect 518878 26898 522836 27134
rect 517800 26856 522836 26898
rect 1104 14454 2200 14496
rect 1104 14218 1706 14454
rect 1942 14218 2200 14454
rect 1104 14134 2200 14218
rect 1104 13898 1706 14134
rect 1942 13898 2200 14134
rect 1104 13856 2200 13898
rect 109800 14454 120200 14496
rect 109800 14218 109998 14454
rect 110234 14218 119706 14454
rect 119942 14218 120200 14454
rect 109800 14134 120200 14218
rect 109800 13898 109998 14134
rect 110234 13898 119706 14134
rect 119942 13898 120200 14134
rect 109800 13856 120200 13898
rect 517800 14454 522836 14496
rect 517800 14218 517982 14454
rect 518218 14218 522836 14454
rect 517800 14134 522836 14218
rect 517800 13898 517982 14134
rect 518218 13898 522836 14134
rect 517800 13856 522836 13898
use mgmt_core  core
timestamp 1638404839
transform 1 0 119000 0 1 2000
box 0 0 400000 148000
use DFFRAM  DFFRAM
timestamp 1638404839
transform 1 0 1000 0 1 2000
box 4 0 110000 148000
<< labels >>
rlabel metal5 s 1104 26856 2200 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 26856 120200 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 26856 522836 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 52856 2200 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 52856 120200 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 52856 522836 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 78856 2200 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 78856 120200 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 78856 522836 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 104856 2200 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 104856 120200 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 104856 522836 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 130856 2200 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 130856 120200 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 130856 522836 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 156856 522836 157496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 13856 2200 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 13856 120200 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 13856 522836 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 39856 2200 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 39856 120200 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 39856 522836 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 65856 2200 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 65856 120200 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 65856 522836 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 91856 2200 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 91856 120200 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 91856 522836 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 117856 2200 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 117856 120200 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 117856 522836 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 143856 2200 144496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 143856 120200 144496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 143856 522836 144496 6 VPWR
port 1 nsew power input
rlabel metal2 s 294786 -400 294842 800 6 core_clk
port 2 nsew signal input
rlabel metal2 s 98274 -400 98330 800 6 core_rstn
port 3 nsew signal input
rlabel metal3 s 523200 64472 524400 64592 6 debug_in
port 4 nsew signal input
rlabel metal3 s 523200 65968 524400 66088 6 debug_mode
port 5 nsew signal tristate
rlabel metal3 s 523200 67464 524400 67584 6 debug_oeb
port 6 nsew signal tristate
rlabel metal3 s 523200 68960 524400 69080 6 debug_out
port 7 nsew signal tristate
rlabel metal3 s 523200 144848 524400 144968 6 flash_clk
port 8 nsew signal tristate
rlabel metal3 s 523200 143352 524400 143472 6 flash_csb
port 9 nsew signal tristate
rlabel metal3 s 523200 146480 524400 146600 6 flash_io0_di
port 10 nsew signal input
rlabel metal3 s 523200 147976 524400 148096 6 flash_io0_do
port 11 nsew signal tristate
rlabel metal3 s 523200 149472 524400 149592 6 flash_io0_oeb
port 12 nsew signal tristate
rlabel metal3 s 523200 150968 524400 151088 6 flash_io1_di
port 13 nsew signal input
rlabel metal3 s 523200 152464 524400 152584 6 flash_io1_do
port 14 nsew signal tristate
rlabel metal3 s 523200 153960 524400 154080 6 flash_io1_oeb
port 15 nsew signal tristate
rlabel metal3 s 523200 155592 524400 155712 6 flash_io2_di
port 16 nsew signal input
rlabel metal3 s 523200 157088 524400 157208 6 flash_io2_do
port 17 nsew signal tristate
rlabel metal3 s 523200 158584 524400 158704 6 flash_io2_oeb
port 18 nsew signal tristate
rlabel metal3 s 523200 160080 524400 160200 6 flash_io3_di
port 19 nsew signal input
rlabel metal3 s 523200 161576 524400 161696 6 flash_io3_do
port 20 nsew signal tristate
rlabel metal3 s 523200 163072 524400 163192 6 flash_io3_oeb
port 21 nsew signal tristate
rlabel metal2 s 32770 -400 32826 800 6 gpio_in_pad
port 22 nsew signal input
rlabel metal2 s 163778 -400 163834 800 6 gpio_inenb_pad
port 23 nsew signal tristate
rlabel metal2 s 229282 -400 229338 800 6 gpio_mode0_pad
port 24 nsew signal tristate
rlabel metal2 s 360290 -400 360346 800 6 gpio_mode1_pad
port 25 nsew signal tristate
rlabel metal2 s 425794 -400 425850 800 6 gpio_out_pad
port 26 nsew signal tristate
rlabel metal2 s 491298 -400 491354 800 6 gpio_outenb_pad
port 27 nsew signal tristate
rlabel metal3 s 523200 91808 524400 91928 6 hk_ack_i
port 28 nsew signal input
rlabel metal2 s 523498 163200 523554 164400 6 hk_cyc_o
port 29 nsew signal tristate
rlabel metal3 s 523200 94800 524400 94920 6 hk_dat_i[0]
port 30 nsew signal input
rlabel metal3 s 523200 110032 524400 110152 6 hk_dat_i[10]
port 31 nsew signal input
rlabel metal3 s 523200 111528 524400 111648 6 hk_dat_i[11]
port 32 nsew signal input
rlabel metal3 s 523200 113024 524400 113144 6 hk_dat_i[12]
port 33 nsew signal input
rlabel metal3 s 523200 114520 524400 114640 6 hk_dat_i[13]
port 34 nsew signal input
rlabel metal3 s 523200 116016 524400 116136 6 hk_dat_i[14]
port 35 nsew signal input
rlabel metal3 s 523200 117512 524400 117632 6 hk_dat_i[15]
port 36 nsew signal input
rlabel metal3 s 523200 119144 524400 119264 6 hk_dat_i[16]
port 37 nsew signal input
rlabel metal3 s 523200 120640 524400 120760 6 hk_dat_i[17]
port 38 nsew signal input
rlabel metal3 s 523200 122136 524400 122256 6 hk_dat_i[18]
port 39 nsew signal input
rlabel metal3 s 523200 123632 524400 123752 6 hk_dat_i[19]
port 40 nsew signal input
rlabel metal3 s 523200 96296 524400 96416 6 hk_dat_i[1]
port 41 nsew signal input
rlabel metal3 s 523200 125128 524400 125248 6 hk_dat_i[20]
port 42 nsew signal input
rlabel metal3 s 523200 126624 524400 126744 6 hk_dat_i[21]
port 43 nsew signal input
rlabel metal3 s 523200 128256 524400 128376 6 hk_dat_i[22]
port 44 nsew signal input
rlabel metal3 s 523200 129752 524400 129872 6 hk_dat_i[23]
port 45 nsew signal input
rlabel metal3 s 523200 131248 524400 131368 6 hk_dat_i[24]
port 46 nsew signal input
rlabel metal3 s 523200 132744 524400 132864 6 hk_dat_i[25]
port 47 nsew signal input
rlabel metal3 s 523200 134240 524400 134360 6 hk_dat_i[26]
port 48 nsew signal input
rlabel metal3 s 523200 135736 524400 135856 6 hk_dat_i[27]
port 49 nsew signal input
rlabel metal3 s 523200 137368 524400 137488 6 hk_dat_i[28]
port 50 nsew signal input
rlabel metal3 s 523200 138864 524400 138984 6 hk_dat_i[29]
port 51 nsew signal input
rlabel metal3 s 523200 97792 524400 97912 6 hk_dat_i[2]
port 52 nsew signal input
rlabel metal3 s 523200 140360 524400 140480 6 hk_dat_i[30]
port 53 nsew signal input
rlabel metal3 s 523200 141856 524400 141976 6 hk_dat_i[31]
port 54 nsew signal input
rlabel metal3 s 523200 99288 524400 99408 6 hk_dat_i[3]
port 55 nsew signal input
rlabel metal3 s 523200 100920 524400 101040 6 hk_dat_i[4]
port 56 nsew signal input
rlabel metal3 s 523200 102416 524400 102536 6 hk_dat_i[5]
port 57 nsew signal input
rlabel metal3 s 523200 103912 524400 104032 6 hk_dat_i[6]
port 58 nsew signal input
rlabel metal3 s 523200 105408 524400 105528 6 hk_dat_i[7]
port 59 nsew signal input
rlabel metal3 s 523200 106904 524400 107024 6 hk_dat_i[8]
port 60 nsew signal input
rlabel metal3 s 523200 108400 524400 108520 6 hk_dat_i[9]
port 61 nsew signal input
rlabel metal3 s 523200 93304 524400 93424 6 hk_stb_o
port 62 nsew signal tristate
rlabel metal2 s 521014 163200 521070 164400 6 irq[0]
port 63 nsew signal input
rlabel metal2 s 521842 163200 521898 164400 6 irq[1]
port 64 nsew signal input
rlabel metal2 s 522670 163200 522726 164400 6 irq[2]
port 65 nsew signal input
rlabel metal3 s 523200 75080 524400 75200 6 irq[3]
port 66 nsew signal input
rlabel metal3 s 523200 73584 524400 73704 6 irq[4]
port 67 nsew signal input
rlabel metal3 s 523200 71952 524400 72072 6 irq[5]
port 68 nsew signal input
rlabel metal2 s 386 163200 442 164400 6 la_iena[0]
port 69 nsew signal tristate
rlabel metal2 s 336278 163200 336334 164400 6 la_iena[100]
port 70 nsew signal tristate
rlabel metal2 s 339590 163200 339646 164400 6 la_iena[101]
port 71 nsew signal tristate
rlabel metal2 s 342994 163200 343050 164400 6 la_iena[102]
port 72 nsew signal tristate
rlabel metal2 s 346306 163200 346362 164400 6 la_iena[103]
port 73 nsew signal tristate
rlabel metal2 s 349710 163200 349766 164400 6 la_iena[104]
port 74 nsew signal tristate
rlabel metal2 s 353022 163200 353078 164400 6 la_iena[105]
port 75 nsew signal tristate
rlabel metal2 s 356426 163200 356482 164400 6 la_iena[106]
port 76 nsew signal tristate
rlabel metal2 s 359738 163200 359794 164400 6 la_iena[107]
port 77 nsew signal tristate
rlabel metal2 s 363142 163200 363198 164400 6 la_iena[108]
port 78 nsew signal tristate
rlabel metal2 s 366454 163200 366510 164400 6 la_iena[109]
port 79 nsew signal tristate
rlabel metal2 s 33966 163200 34022 164400 6 la_iena[10]
port 80 nsew signal tristate
rlabel metal2 s 369858 163200 369914 164400 6 la_iena[110]
port 81 nsew signal tristate
rlabel metal2 s 373170 163200 373226 164400 6 la_iena[111]
port 82 nsew signal tristate
rlabel metal2 s 376574 163200 376630 164400 6 la_iena[112]
port 83 nsew signal tristate
rlabel metal2 s 379886 163200 379942 164400 6 la_iena[113]
port 84 nsew signal tristate
rlabel metal2 s 383290 163200 383346 164400 6 la_iena[114]
port 85 nsew signal tristate
rlabel metal2 s 386602 163200 386658 164400 6 la_iena[115]
port 86 nsew signal tristate
rlabel metal2 s 390006 163200 390062 164400 6 la_iena[116]
port 87 nsew signal tristate
rlabel metal2 s 393410 163200 393466 164400 6 la_iena[117]
port 88 nsew signal tristate
rlabel metal2 s 396722 163200 396778 164400 6 la_iena[118]
port 89 nsew signal tristate
rlabel metal2 s 400126 163200 400182 164400 6 la_iena[119]
port 90 nsew signal tristate
rlabel metal2 s 37278 163200 37334 164400 6 la_iena[11]
port 91 nsew signal tristate
rlabel metal2 s 403438 163200 403494 164400 6 la_iena[120]
port 92 nsew signal tristate
rlabel metal2 s 406842 163200 406898 164400 6 la_iena[121]
port 93 nsew signal tristate
rlabel metal2 s 410154 163200 410210 164400 6 la_iena[122]
port 94 nsew signal tristate
rlabel metal2 s 413558 163200 413614 164400 6 la_iena[123]
port 95 nsew signal tristate
rlabel metal2 s 416870 163200 416926 164400 6 la_iena[124]
port 96 nsew signal tristate
rlabel metal2 s 420274 163200 420330 164400 6 la_iena[125]
port 97 nsew signal tristate
rlabel metal2 s 423586 163200 423642 164400 6 la_iena[126]
port 98 nsew signal tristate
rlabel metal2 s 426990 163200 427046 164400 6 la_iena[127]
port 99 nsew signal tristate
rlabel metal2 s 40682 163200 40738 164400 6 la_iena[12]
port 100 nsew signal tristate
rlabel metal2 s 43994 163200 44050 164400 6 la_iena[13]
port 101 nsew signal tristate
rlabel metal2 s 47398 163200 47454 164400 6 la_iena[14]
port 102 nsew signal tristate
rlabel metal2 s 50710 163200 50766 164400 6 la_iena[15]
port 103 nsew signal tristate
rlabel metal2 s 54114 163200 54170 164400 6 la_iena[16]
port 104 nsew signal tristate
rlabel metal2 s 57426 163200 57482 164400 6 la_iena[17]
port 105 nsew signal tristate
rlabel metal2 s 60830 163200 60886 164400 6 la_iena[18]
port 106 nsew signal tristate
rlabel metal2 s 64142 163200 64198 164400 6 la_iena[19]
port 107 nsew signal tristate
rlabel metal2 s 3698 163200 3754 164400 6 la_iena[1]
port 108 nsew signal tristate
rlabel metal2 s 67546 163200 67602 164400 6 la_iena[20]
port 109 nsew signal tristate
rlabel metal2 s 70858 163200 70914 164400 6 la_iena[21]
port 110 nsew signal tristate
rlabel metal2 s 74262 163200 74318 164400 6 la_iena[22]
port 111 nsew signal tristate
rlabel metal2 s 77574 163200 77630 164400 6 la_iena[23]
port 112 nsew signal tristate
rlabel metal2 s 80978 163200 81034 164400 6 la_iena[24]
port 113 nsew signal tristate
rlabel metal2 s 84290 163200 84346 164400 6 la_iena[25]
port 114 nsew signal tristate
rlabel metal2 s 87694 163200 87750 164400 6 la_iena[26]
port 115 nsew signal tristate
rlabel metal2 s 91006 163200 91062 164400 6 la_iena[27]
port 116 nsew signal tristate
rlabel metal2 s 94410 163200 94466 164400 6 la_iena[28]
port 117 nsew signal tristate
rlabel metal2 s 97722 163200 97778 164400 6 la_iena[29]
port 118 nsew signal tristate
rlabel metal2 s 7102 163200 7158 164400 6 la_iena[2]
port 119 nsew signal tristate
rlabel metal2 s 101126 163200 101182 164400 6 la_iena[30]
port 120 nsew signal tristate
rlabel metal2 s 104438 163200 104494 164400 6 la_iena[31]
port 121 nsew signal tristate
rlabel metal2 s 107842 163200 107898 164400 6 la_iena[32]
port 122 nsew signal tristate
rlabel metal2 s 111154 163200 111210 164400 6 la_iena[33]
port 123 nsew signal tristate
rlabel metal2 s 114558 163200 114614 164400 6 la_iena[34]
port 124 nsew signal tristate
rlabel metal2 s 117870 163200 117926 164400 6 la_iena[35]
port 125 nsew signal tristate
rlabel metal2 s 121274 163200 121330 164400 6 la_iena[36]
port 126 nsew signal tristate
rlabel metal2 s 124586 163200 124642 164400 6 la_iena[37]
port 127 nsew signal tristate
rlabel metal2 s 127990 163200 128046 164400 6 la_iena[38]
port 128 nsew signal tristate
rlabel metal2 s 131394 163200 131450 164400 6 la_iena[39]
port 129 nsew signal tristate
rlabel metal2 s 10414 163200 10470 164400 6 la_iena[3]
port 130 nsew signal tristate
rlabel metal2 s 134706 163200 134762 164400 6 la_iena[40]
port 131 nsew signal tristate
rlabel metal2 s 138110 163200 138166 164400 6 la_iena[41]
port 132 nsew signal tristate
rlabel metal2 s 141422 163200 141478 164400 6 la_iena[42]
port 133 nsew signal tristate
rlabel metal2 s 144826 163200 144882 164400 6 la_iena[43]
port 134 nsew signal tristate
rlabel metal2 s 148138 163200 148194 164400 6 la_iena[44]
port 135 nsew signal tristate
rlabel metal2 s 151542 163200 151598 164400 6 la_iena[45]
port 136 nsew signal tristate
rlabel metal2 s 154854 163200 154910 164400 6 la_iena[46]
port 137 nsew signal tristate
rlabel metal2 s 158258 163200 158314 164400 6 la_iena[47]
port 138 nsew signal tristate
rlabel metal2 s 161570 163200 161626 164400 6 la_iena[48]
port 139 nsew signal tristate
rlabel metal2 s 164974 163200 165030 164400 6 la_iena[49]
port 140 nsew signal tristate
rlabel metal2 s 13818 163200 13874 164400 6 la_iena[4]
port 141 nsew signal tristate
rlabel metal2 s 168286 163200 168342 164400 6 la_iena[50]
port 142 nsew signal tristate
rlabel metal2 s 171690 163200 171746 164400 6 la_iena[51]
port 143 nsew signal tristate
rlabel metal2 s 175002 163200 175058 164400 6 la_iena[52]
port 144 nsew signal tristate
rlabel metal2 s 178406 163200 178462 164400 6 la_iena[53]
port 145 nsew signal tristate
rlabel metal2 s 181718 163200 181774 164400 6 la_iena[54]
port 146 nsew signal tristate
rlabel metal2 s 185122 163200 185178 164400 6 la_iena[55]
port 147 nsew signal tristate
rlabel metal2 s 188434 163200 188490 164400 6 la_iena[56]
port 148 nsew signal tristate
rlabel metal2 s 191838 163200 191894 164400 6 la_iena[57]
port 149 nsew signal tristate
rlabel metal2 s 195150 163200 195206 164400 6 la_iena[58]
port 150 nsew signal tristate
rlabel metal2 s 198554 163200 198610 164400 6 la_iena[59]
port 151 nsew signal tristate
rlabel metal2 s 17130 163200 17186 164400 6 la_iena[5]
port 152 nsew signal tristate
rlabel metal2 s 201866 163200 201922 164400 6 la_iena[60]
port 153 nsew signal tristate
rlabel metal2 s 205270 163200 205326 164400 6 la_iena[61]
port 154 nsew signal tristate
rlabel metal2 s 208582 163200 208638 164400 6 la_iena[62]
port 155 nsew signal tristate
rlabel metal2 s 211986 163200 212042 164400 6 la_iena[63]
port 156 nsew signal tristate
rlabel metal2 s 215298 163200 215354 164400 6 la_iena[64]
port 157 nsew signal tristate
rlabel metal2 s 218702 163200 218758 164400 6 la_iena[65]
port 158 nsew signal tristate
rlabel metal2 s 222014 163200 222070 164400 6 la_iena[66]
port 159 nsew signal tristate
rlabel metal2 s 225418 163200 225474 164400 6 la_iena[67]
port 160 nsew signal tristate
rlabel metal2 s 228730 163200 228786 164400 6 la_iena[68]
port 161 nsew signal tristate
rlabel metal2 s 232134 163200 232190 164400 6 la_iena[69]
port 162 nsew signal tristate
rlabel metal2 s 20534 163200 20590 164400 6 la_iena[6]
port 163 nsew signal tristate
rlabel metal2 s 235446 163200 235502 164400 6 la_iena[70]
port 164 nsew signal tristate
rlabel metal2 s 238850 163200 238906 164400 6 la_iena[71]
port 165 nsew signal tristate
rlabel metal2 s 242162 163200 242218 164400 6 la_iena[72]
port 166 nsew signal tristate
rlabel metal2 s 245566 163200 245622 164400 6 la_iena[73]
port 167 nsew signal tristate
rlabel metal2 s 248878 163200 248934 164400 6 la_iena[74]
port 168 nsew signal tristate
rlabel metal2 s 252282 163200 252338 164400 6 la_iena[75]
port 169 nsew signal tristate
rlabel metal2 s 255594 163200 255650 164400 6 la_iena[76]
port 170 nsew signal tristate
rlabel metal2 s 258998 163200 259054 164400 6 la_iena[77]
port 171 nsew signal tristate
rlabel metal2 s 262402 163200 262458 164400 6 la_iena[78]
port 172 nsew signal tristate
rlabel metal2 s 265714 163200 265770 164400 6 la_iena[79]
port 173 nsew signal tristate
rlabel metal2 s 23846 163200 23902 164400 6 la_iena[7]
port 174 nsew signal tristate
rlabel metal2 s 269118 163200 269174 164400 6 la_iena[80]
port 175 nsew signal tristate
rlabel metal2 s 272430 163200 272486 164400 6 la_iena[81]
port 176 nsew signal tristate
rlabel metal2 s 275834 163200 275890 164400 6 la_iena[82]
port 177 nsew signal tristate
rlabel metal2 s 279146 163200 279202 164400 6 la_iena[83]
port 178 nsew signal tristate
rlabel metal2 s 282550 163200 282606 164400 6 la_iena[84]
port 179 nsew signal tristate
rlabel metal2 s 285862 163200 285918 164400 6 la_iena[85]
port 180 nsew signal tristate
rlabel metal2 s 289266 163200 289322 164400 6 la_iena[86]
port 181 nsew signal tristate
rlabel metal2 s 292578 163200 292634 164400 6 la_iena[87]
port 182 nsew signal tristate
rlabel metal2 s 295982 163200 296038 164400 6 la_iena[88]
port 183 nsew signal tristate
rlabel metal2 s 299294 163200 299350 164400 6 la_iena[89]
port 184 nsew signal tristate
rlabel metal2 s 27250 163200 27306 164400 6 la_iena[8]
port 185 nsew signal tristate
rlabel metal2 s 302698 163200 302754 164400 6 la_iena[90]
port 186 nsew signal tristate
rlabel metal2 s 306010 163200 306066 164400 6 la_iena[91]
port 187 nsew signal tristate
rlabel metal2 s 309414 163200 309470 164400 6 la_iena[92]
port 188 nsew signal tristate
rlabel metal2 s 312726 163200 312782 164400 6 la_iena[93]
port 189 nsew signal tristate
rlabel metal2 s 316130 163200 316186 164400 6 la_iena[94]
port 190 nsew signal tristate
rlabel metal2 s 319442 163200 319498 164400 6 la_iena[95]
port 191 nsew signal tristate
rlabel metal2 s 322846 163200 322902 164400 6 la_iena[96]
port 192 nsew signal tristate
rlabel metal2 s 326158 163200 326214 164400 6 la_iena[97]
port 193 nsew signal tristate
rlabel metal2 s 329562 163200 329618 164400 6 la_iena[98]
port 194 nsew signal tristate
rlabel metal2 s 332874 163200 332930 164400 6 la_iena[99]
port 195 nsew signal tristate
rlabel metal2 s 30562 163200 30618 164400 6 la_iena[9]
port 196 nsew signal tristate
rlabel metal2 s 1214 163200 1270 164400 6 la_input[0]
port 197 nsew signal input
rlabel metal2 s 337106 163200 337162 164400 6 la_input[100]
port 198 nsew signal input
rlabel metal2 s 340418 163200 340474 164400 6 la_input[101]
port 199 nsew signal input
rlabel metal2 s 343822 163200 343878 164400 6 la_input[102]
port 200 nsew signal input
rlabel metal2 s 347134 163200 347190 164400 6 la_input[103]
port 201 nsew signal input
rlabel metal2 s 350538 163200 350594 164400 6 la_input[104]
port 202 nsew signal input
rlabel metal2 s 353850 163200 353906 164400 6 la_input[105]
port 203 nsew signal input
rlabel metal2 s 357254 163200 357310 164400 6 la_input[106]
port 204 nsew signal input
rlabel metal2 s 360658 163200 360714 164400 6 la_input[107]
port 205 nsew signal input
rlabel metal2 s 363970 163200 364026 164400 6 la_input[108]
port 206 nsew signal input
rlabel metal2 s 367374 163200 367430 164400 6 la_input[109]
port 207 nsew signal input
rlabel metal2 s 34794 163200 34850 164400 6 la_input[10]
port 208 nsew signal input
rlabel metal2 s 370686 163200 370742 164400 6 la_input[110]
port 209 nsew signal input
rlabel metal2 s 374090 163200 374146 164400 6 la_input[111]
port 210 nsew signal input
rlabel metal2 s 377402 163200 377458 164400 6 la_input[112]
port 211 nsew signal input
rlabel metal2 s 380806 163200 380862 164400 6 la_input[113]
port 212 nsew signal input
rlabel metal2 s 384118 163200 384174 164400 6 la_input[114]
port 213 nsew signal input
rlabel metal2 s 387522 163200 387578 164400 6 la_input[115]
port 214 nsew signal input
rlabel metal2 s 390834 163200 390890 164400 6 la_input[116]
port 215 nsew signal input
rlabel metal2 s 394238 163200 394294 164400 6 la_input[117]
port 216 nsew signal input
rlabel metal2 s 397550 163200 397606 164400 6 la_input[118]
port 217 nsew signal input
rlabel metal2 s 400954 163200 401010 164400 6 la_input[119]
port 218 nsew signal input
rlabel metal2 s 38106 163200 38162 164400 6 la_input[11]
port 219 nsew signal input
rlabel metal2 s 404266 163200 404322 164400 6 la_input[120]
port 220 nsew signal input
rlabel metal2 s 407670 163200 407726 164400 6 la_input[121]
port 221 nsew signal input
rlabel metal2 s 410982 163200 411038 164400 6 la_input[122]
port 222 nsew signal input
rlabel metal2 s 414386 163200 414442 164400 6 la_input[123]
port 223 nsew signal input
rlabel metal2 s 417698 163200 417754 164400 6 la_input[124]
port 224 nsew signal input
rlabel metal2 s 421102 163200 421158 164400 6 la_input[125]
port 225 nsew signal input
rlabel metal2 s 424414 163200 424470 164400 6 la_input[126]
port 226 nsew signal input
rlabel metal2 s 427818 163200 427874 164400 6 la_input[127]
port 227 nsew signal input
rlabel metal2 s 41510 163200 41566 164400 6 la_input[12]
port 228 nsew signal input
rlabel metal2 s 44822 163200 44878 164400 6 la_input[13]
port 229 nsew signal input
rlabel metal2 s 48226 163200 48282 164400 6 la_input[14]
port 230 nsew signal input
rlabel metal2 s 51538 163200 51594 164400 6 la_input[15]
port 231 nsew signal input
rlabel metal2 s 54942 163200 54998 164400 6 la_input[16]
port 232 nsew signal input
rlabel metal2 s 58254 163200 58310 164400 6 la_input[17]
port 233 nsew signal input
rlabel metal2 s 61658 163200 61714 164400 6 la_input[18]
port 234 nsew signal input
rlabel metal2 s 64970 163200 65026 164400 6 la_input[19]
port 235 nsew signal input
rlabel metal2 s 4526 163200 4582 164400 6 la_input[1]
port 236 nsew signal input
rlabel metal2 s 68374 163200 68430 164400 6 la_input[20]
port 237 nsew signal input
rlabel metal2 s 71686 163200 71742 164400 6 la_input[21]
port 238 nsew signal input
rlabel metal2 s 75090 163200 75146 164400 6 la_input[22]
port 239 nsew signal input
rlabel metal2 s 78402 163200 78458 164400 6 la_input[23]
port 240 nsew signal input
rlabel metal2 s 81806 163200 81862 164400 6 la_input[24]
port 241 nsew signal input
rlabel metal2 s 85118 163200 85174 164400 6 la_input[25]
port 242 nsew signal input
rlabel metal2 s 88522 163200 88578 164400 6 la_input[26]
port 243 nsew signal input
rlabel metal2 s 91834 163200 91890 164400 6 la_input[27]
port 244 nsew signal input
rlabel metal2 s 95238 163200 95294 164400 6 la_input[28]
port 245 nsew signal input
rlabel metal2 s 98642 163200 98698 164400 6 la_input[29]
port 246 nsew signal input
rlabel metal2 s 7930 163200 7986 164400 6 la_input[2]
port 247 nsew signal input
rlabel metal2 s 101954 163200 102010 164400 6 la_input[30]
port 248 nsew signal input
rlabel metal2 s 105358 163200 105414 164400 6 la_input[31]
port 249 nsew signal input
rlabel metal2 s 108670 163200 108726 164400 6 la_input[32]
port 250 nsew signal input
rlabel metal2 s 112074 163200 112130 164400 6 la_input[33]
port 251 nsew signal input
rlabel metal2 s 115386 163200 115442 164400 6 la_input[34]
port 252 nsew signal input
rlabel metal2 s 118790 163200 118846 164400 6 la_input[35]
port 253 nsew signal input
rlabel metal2 s 122102 163200 122158 164400 6 la_input[36]
port 254 nsew signal input
rlabel metal2 s 125506 163200 125562 164400 6 la_input[37]
port 255 nsew signal input
rlabel metal2 s 128818 163200 128874 164400 6 la_input[38]
port 256 nsew signal input
rlabel metal2 s 132222 163200 132278 164400 6 la_input[39]
port 257 nsew signal input
rlabel metal2 s 11242 163200 11298 164400 6 la_input[3]
port 258 nsew signal input
rlabel metal2 s 135534 163200 135590 164400 6 la_input[40]
port 259 nsew signal input
rlabel metal2 s 138938 163200 138994 164400 6 la_input[41]
port 260 nsew signal input
rlabel metal2 s 142250 163200 142306 164400 6 la_input[42]
port 261 nsew signal input
rlabel metal2 s 145654 163200 145710 164400 6 la_input[43]
port 262 nsew signal input
rlabel metal2 s 148966 163200 149022 164400 6 la_input[44]
port 263 nsew signal input
rlabel metal2 s 152370 163200 152426 164400 6 la_input[45]
port 264 nsew signal input
rlabel metal2 s 155682 163200 155738 164400 6 la_input[46]
port 265 nsew signal input
rlabel metal2 s 159086 163200 159142 164400 6 la_input[47]
port 266 nsew signal input
rlabel metal2 s 162398 163200 162454 164400 6 la_input[48]
port 267 nsew signal input
rlabel metal2 s 165802 163200 165858 164400 6 la_input[49]
port 268 nsew signal input
rlabel metal2 s 14646 163200 14702 164400 6 la_input[4]
port 269 nsew signal input
rlabel metal2 s 169114 163200 169170 164400 6 la_input[50]
port 270 nsew signal input
rlabel metal2 s 172518 163200 172574 164400 6 la_input[51]
port 271 nsew signal input
rlabel metal2 s 175830 163200 175886 164400 6 la_input[52]
port 272 nsew signal input
rlabel metal2 s 179234 163200 179290 164400 6 la_input[53]
port 273 nsew signal input
rlabel metal2 s 182546 163200 182602 164400 6 la_input[54]
port 274 nsew signal input
rlabel metal2 s 185950 163200 186006 164400 6 la_input[55]
port 275 nsew signal input
rlabel metal2 s 189262 163200 189318 164400 6 la_input[56]
port 276 nsew signal input
rlabel metal2 s 192666 163200 192722 164400 6 la_input[57]
port 277 nsew signal input
rlabel metal2 s 195978 163200 196034 164400 6 la_input[58]
port 278 nsew signal input
rlabel metal2 s 199382 163200 199438 164400 6 la_input[59]
port 279 nsew signal input
rlabel metal2 s 17958 163200 18014 164400 6 la_input[5]
port 280 nsew signal input
rlabel metal2 s 202694 163200 202750 164400 6 la_input[60]
port 281 nsew signal input
rlabel metal2 s 206098 163200 206154 164400 6 la_input[61]
port 282 nsew signal input
rlabel metal2 s 209410 163200 209466 164400 6 la_input[62]
port 283 nsew signal input
rlabel metal2 s 212814 163200 212870 164400 6 la_input[63]
port 284 nsew signal input
rlabel metal2 s 216126 163200 216182 164400 6 la_input[64]
port 285 nsew signal input
rlabel metal2 s 219530 163200 219586 164400 6 la_input[65]
port 286 nsew signal input
rlabel metal2 s 222842 163200 222898 164400 6 la_input[66]
port 287 nsew signal input
rlabel metal2 s 226246 163200 226302 164400 6 la_input[67]
port 288 nsew signal input
rlabel metal2 s 229650 163200 229706 164400 6 la_input[68]
port 289 nsew signal input
rlabel metal2 s 232962 163200 233018 164400 6 la_input[69]
port 290 nsew signal input
rlabel metal2 s 21362 163200 21418 164400 6 la_input[6]
port 291 nsew signal input
rlabel metal2 s 236366 163200 236422 164400 6 la_input[70]
port 292 nsew signal input
rlabel metal2 s 239678 163200 239734 164400 6 la_input[71]
port 293 nsew signal input
rlabel metal2 s 243082 163200 243138 164400 6 la_input[72]
port 294 nsew signal input
rlabel metal2 s 246394 163200 246450 164400 6 la_input[73]
port 295 nsew signal input
rlabel metal2 s 249798 163200 249854 164400 6 la_input[74]
port 296 nsew signal input
rlabel metal2 s 253110 163200 253166 164400 6 la_input[75]
port 297 nsew signal input
rlabel metal2 s 256514 163200 256570 164400 6 la_input[76]
port 298 nsew signal input
rlabel metal2 s 259826 163200 259882 164400 6 la_input[77]
port 299 nsew signal input
rlabel metal2 s 263230 163200 263286 164400 6 la_input[78]
port 300 nsew signal input
rlabel metal2 s 266542 163200 266598 164400 6 la_input[79]
port 301 nsew signal input
rlabel metal2 s 24674 163200 24730 164400 6 la_input[7]
port 302 nsew signal input
rlabel metal2 s 269946 163200 270002 164400 6 la_input[80]
port 303 nsew signal input
rlabel metal2 s 273258 163200 273314 164400 6 la_input[81]
port 304 nsew signal input
rlabel metal2 s 276662 163200 276718 164400 6 la_input[82]
port 305 nsew signal input
rlabel metal2 s 279974 163200 280030 164400 6 la_input[83]
port 306 nsew signal input
rlabel metal2 s 283378 163200 283434 164400 6 la_input[84]
port 307 nsew signal input
rlabel metal2 s 286690 163200 286746 164400 6 la_input[85]
port 308 nsew signal input
rlabel metal2 s 290094 163200 290150 164400 6 la_input[86]
port 309 nsew signal input
rlabel metal2 s 293406 163200 293462 164400 6 la_input[87]
port 310 nsew signal input
rlabel metal2 s 296810 163200 296866 164400 6 la_input[88]
port 311 nsew signal input
rlabel metal2 s 300122 163200 300178 164400 6 la_input[89]
port 312 nsew signal input
rlabel metal2 s 28078 163200 28134 164400 6 la_input[8]
port 313 nsew signal input
rlabel metal2 s 303526 163200 303582 164400 6 la_input[90]
port 314 nsew signal input
rlabel metal2 s 306838 163200 306894 164400 6 la_input[91]
port 315 nsew signal input
rlabel metal2 s 310242 163200 310298 164400 6 la_input[92]
port 316 nsew signal input
rlabel metal2 s 313554 163200 313610 164400 6 la_input[93]
port 317 nsew signal input
rlabel metal2 s 316958 163200 317014 164400 6 la_input[94]
port 318 nsew signal input
rlabel metal2 s 320270 163200 320326 164400 6 la_input[95]
port 319 nsew signal input
rlabel metal2 s 323674 163200 323730 164400 6 la_input[96]
port 320 nsew signal input
rlabel metal2 s 326986 163200 327042 164400 6 la_input[97]
port 321 nsew signal input
rlabel metal2 s 330390 163200 330446 164400 6 la_input[98]
port 322 nsew signal input
rlabel metal2 s 333702 163200 333758 164400 6 la_input[99]
port 323 nsew signal input
rlabel metal2 s 31390 163200 31446 164400 6 la_input[9]
port 324 nsew signal input
rlabel metal2 s 2042 163200 2098 164400 6 la_oenb[0]
port 325 nsew signal tristate
rlabel metal2 s 337934 163200 337990 164400 6 la_oenb[100]
port 326 nsew signal tristate
rlabel metal2 s 341338 163200 341394 164400 6 la_oenb[101]
port 327 nsew signal tristate
rlabel metal2 s 344650 163200 344706 164400 6 la_oenb[102]
port 328 nsew signal tristate
rlabel metal2 s 348054 163200 348110 164400 6 la_oenb[103]
port 329 nsew signal tristate
rlabel metal2 s 351366 163200 351422 164400 6 la_oenb[104]
port 330 nsew signal tristate
rlabel metal2 s 354770 163200 354826 164400 6 la_oenb[105]
port 331 nsew signal tristate
rlabel metal2 s 358082 163200 358138 164400 6 la_oenb[106]
port 332 nsew signal tristate
rlabel metal2 s 361486 163200 361542 164400 6 la_oenb[107]
port 333 nsew signal tristate
rlabel metal2 s 364798 163200 364854 164400 6 la_oenb[108]
port 334 nsew signal tristate
rlabel metal2 s 368202 163200 368258 164400 6 la_oenb[109]
port 335 nsew signal tristate
rlabel metal2 s 35622 163200 35678 164400 6 la_oenb[10]
port 336 nsew signal tristate
rlabel metal2 s 371514 163200 371570 164400 6 la_oenb[110]
port 337 nsew signal tristate
rlabel metal2 s 374918 163200 374974 164400 6 la_oenb[111]
port 338 nsew signal tristate
rlabel metal2 s 378230 163200 378286 164400 6 la_oenb[112]
port 339 nsew signal tristate
rlabel metal2 s 381634 163200 381690 164400 6 la_oenb[113]
port 340 nsew signal tristate
rlabel metal2 s 384946 163200 385002 164400 6 la_oenb[114]
port 341 nsew signal tristate
rlabel metal2 s 388350 163200 388406 164400 6 la_oenb[115]
port 342 nsew signal tristate
rlabel metal2 s 391662 163200 391718 164400 6 la_oenb[116]
port 343 nsew signal tristate
rlabel metal2 s 395066 163200 395122 164400 6 la_oenb[117]
port 344 nsew signal tristate
rlabel metal2 s 398378 163200 398434 164400 6 la_oenb[118]
port 345 nsew signal tristate
rlabel metal2 s 401782 163200 401838 164400 6 la_oenb[119]
port 346 nsew signal tristate
rlabel metal2 s 38934 163200 38990 164400 6 la_oenb[11]
port 347 nsew signal tristate
rlabel metal2 s 405094 163200 405150 164400 6 la_oenb[120]
port 348 nsew signal tristate
rlabel metal2 s 408498 163200 408554 164400 6 la_oenb[121]
port 349 nsew signal tristate
rlabel metal2 s 411810 163200 411866 164400 6 la_oenb[122]
port 350 nsew signal tristate
rlabel metal2 s 415214 163200 415270 164400 6 la_oenb[123]
port 351 nsew signal tristate
rlabel metal2 s 418526 163200 418582 164400 6 la_oenb[124]
port 352 nsew signal tristate
rlabel metal2 s 421930 163200 421986 164400 6 la_oenb[125]
port 353 nsew signal tristate
rlabel metal2 s 425242 163200 425298 164400 6 la_oenb[126]
port 354 nsew signal tristate
rlabel metal2 s 428646 163200 428702 164400 6 la_oenb[127]
port 355 nsew signal tristate
rlabel metal2 s 42338 163200 42394 164400 6 la_oenb[12]
port 356 nsew signal tristate
rlabel metal2 s 45650 163200 45706 164400 6 la_oenb[13]
port 357 nsew signal tristate
rlabel metal2 s 49054 163200 49110 164400 6 la_oenb[14]
port 358 nsew signal tristate
rlabel metal2 s 52366 163200 52422 164400 6 la_oenb[15]
port 359 nsew signal tristate
rlabel metal2 s 55770 163200 55826 164400 6 la_oenb[16]
port 360 nsew signal tristate
rlabel metal2 s 59082 163200 59138 164400 6 la_oenb[17]
port 361 nsew signal tristate
rlabel metal2 s 62486 163200 62542 164400 6 la_oenb[18]
port 362 nsew signal tristate
rlabel metal2 s 65890 163200 65946 164400 6 la_oenb[19]
port 363 nsew signal tristate
rlabel metal2 s 5354 163200 5410 164400 6 la_oenb[1]
port 364 nsew signal tristate
rlabel metal2 s 69202 163200 69258 164400 6 la_oenb[20]
port 365 nsew signal tristate
rlabel metal2 s 72606 163200 72662 164400 6 la_oenb[21]
port 366 nsew signal tristate
rlabel metal2 s 75918 163200 75974 164400 6 la_oenb[22]
port 367 nsew signal tristate
rlabel metal2 s 79322 163200 79378 164400 6 la_oenb[23]
port 368 nsew signal tristate
rlabel metal2 s 82634 163200 82690 164400 6 la_oenb[24]
port 369 nsew signal tristate
rlabel metal2 s 86038 163200 86094 164400 6 la_oenb[25]
port 370 nsew signal tristate
rlabel metal2 s 89350 163200 89406 164400 6 la_oenb[26]
port 371 nsew signal tristate
rlabel metal2 s 92754 163200 92810 164400 6 la_oenb[27]
port 372 nsew signal tristate
rlabel metal2 s 96066 163200 96122 164400 6 la_oenb[28]
port 373 nsew signal tristate
rlabel metal2 s 99470 163200 99526 164400 6 la_oenb[29]
port 374 nsew signal tristate
rlabel metal2 s 8758 163200 8814 164400 6 la_oenb[2]
port 375 nsew signal tristate
rlabel metal2 s 102782 163200 102838 164400 6 la_oenb[30]
port 376 nsew signal tristate
rlabel metal2 s 106186 163200 106242 164400 6 la_oenb[31]
port 377 nsew signal tristate
rlabel metal2 s 109498 163200 109554 164400 6 la_oenb[32]
port 378 nsew signal tristate
rlabel metal2 s 112902 163200 112958 164400 6 la_oenb[33]
port 379 nsew signal tristate
rlabel metal2 s 116214 163200 116270 164400 6 la_oenb[34]
port 380 nsew signal tristate
rlabel metal2 s 119618 163200 119674 164400 6 la_oenb[35]
port 381 nsew signal tristate
rlabel metal2 s 122930 163200 122986 164400 6 la_oenb[36]
port 382 nsew signal tristate
rlabel metal2 s 126334 163200 126390 164400 6 la_oenb[37]
port 383 nsew signal tristate
rlabel metal2 s 129646 163200 129702 164400 6 la_oenb[38]
port 384 nsew signal tristate
rlabel metal2 s 133050 163200 133106 164400 6 la_oenb[39]
port 385 nsew signal tristate
rlabel metal2 s 12070 163200 12126 164400 6 la_oenb[3]
port 386 nsew signal tristate
rlabel metal2 s 136362 163200 136418 164400 6 la_oenb[40]
port 387 nsew signal tristate
rlabel metal2 s 139766 163200 139822 164400 6 la_oenb[41]
port 388 nsew signal tristate
rlabel metal2 s 143078 163200 143134 164400 6 la_oenb[42]
port 389 nsew signal tristate
rlabel metal2 s 146482 163200 146538 164400 6 la_oenb[43]
port 390 nsew signal tristate
rlabel metal2 s 149794 163200 149850 164400 6 la_oenb[44]
port 391 nsew signal tristate
rlabel metal2 s 153198 163200 153254 164400 6 la_oenb[45]
port 392 nsew signal tristate
rlabel metal2 s 156510 163200 156566 164400 6 la_oenb[46]
port 393 nsew signal tristate
rlabel metal2 s 159914 163200 159970 164400 6 la_oenb[47]
port 394 nsew signal tristate
rlabel metal2 s 163226 163200 163282 164400 6 la_oenb[48]
port 395 nsew signal tristate
rlabel metal2 s 166630 163200 166686 164400 6 la_oenb[49]
port 396 nsew signal tristate
rlabel metal2 s 15474 163200 15530 164400 6 la_oenb[4]
port 397 nsew signal tristate
rlabel metal2 s 169942 163200 169998 164400 6 la_oenb[50]
port 398 nsew signal tristate
rlabel metal2 s 173346 163200 173402 164400 6 la_oenb[51]
port 399 nsew signal tristate
rlabel metal2 s 176658 163200 176714 164400 6 la_oenb[52]
port 400 nsew signal tristate
rlabel metal2 s 180062 163200 180118 164400 6 la_oenb[53]
port 401 nsew signal tristate
rlabel metal2 s 183374 163200 183430 164400 6 la_oenb[54]
port 402 nsew signal tristate
rlabel metal2 s 186778 163200 186834 164400 6 la_oenb[55]
port 403 nsew signal tristate
rlabel metal2 s 190090 163200 190146 164400 6 la_oenb[56]
port 404 nsew signal tristate
rlabel metal2 s 193494 163200 193550 164400 6 la_oenb[57]
port 405 nsew signal tristate
rlabel metal2 s 196898 163200 196954 164400 6 la_oenb[58]
port 406 nsew signal tristate
rlabel metal2 s 200210 163200 200266 164400 6 la_oenb[59]
port 407 nsew signal tristate
rlabel metal2 s 18786 163200 18842 164400 6 la_oenb[5]
port 408 nsew signal tristate
rlabel metal2 s 203614 163200 203670 164400 6 la_oenb[60]
port 409 nsew signal tristate
rlabel metal2 s 206926 163200 206982 164400 6 la_oenb[61]
port 410 nsew signal tristate
rlabel metal2 s 210330 163200 210386 164400 6 la_oenb[62]
port 411 nsew signal tristate
rlabel metal2 s 213642 163200 213698 164400 6 la_oenb[63]
port 412 nsew signal tristate
rlabel metal2 s 217046 163200 217102 164400 6 la_oenb[64]
port 413 nsew signal tristate
rlabel metal2 s 220358 163200 220414 164400 6 la_oenb[65]
port 414 nsew signal tristate
rlabel metal2 s 223762 163200 223818 164400 6 la_oenb[66]
port 415 nsew signal tristate
rlabel metal2 s 227074 163200 227130 164400 6 la_oenb[67]
port 416 nsew signal tristate
rlabel metal2 s 230478 163200 230534 164400 6 la_oenb[68]
port 417 nsew signal tristate
rlabel metal2 s 233790 163200 233846 164400 6 la_oenb[69]
port 418 nsew signal tristate
rlabel metal2 s 22190 163200 22246 164400 6 la_oenb[6]
port 419 nsew signal tristate
rlabel metal2 s 237194 163200 237250 164400 6 la_oenb[70]
port 420 nsew signal tristate
rlabel metal2 s 240506 163200 240562 164400 6 la_oenb[71]
port 421 nsew signal tristate
rlabel metal2 s 243910 163200 243966 164400 6 la_oenb[72]
port 422 nsew signal tristate
rlabel metal2 s 247222 163200 247278 164400 6 la_oenb[73]
port 423 nsew signal tristate
rlabel metal2 s 250626 163200 250682 164400 6 la_oenb[74]
port 424 nsew signal tristate
rlabel metal2 s 253938 163200 253994 164400 6 la_oenb[75]
port 425 nsew signal tristate
rlabel metal2 s 257342 163200 257398 164400 6 la_oenb[76]
port 426 nsew signal tristate
rlabel metal2 s 260654 163200 260710 164400 6 la_oenb[77]
port 427 nsew signal tristate
rlabel metal2 s 264058 163200 264114 164400 6 la_oenb[78]
port 428 nsew signal tristate
rlabel metal2 s 267370 163200 267426 164400 6 la_oenb[79]
port 429 nsew signal tristate
rlabel metal2 s 25502 163200 25558 164400 6 la_oenb[7]
port 430 nsew signal tristate
rlabel metal2 s 270774 163200 270830 164400 6 la_oenb[80]
port 431 nsew signal tristate
rlabel metal2 s 274086 163200 274142 164400 6 la_oenb[81]
port 432 nsew signal tristate
rlabel metal2 s 277490 163200 277546 164400 6 la_oenb[82]
port 433 nsew signal tristate
rlabel metal2 s 280802 163200 280858 164400 6 la_oenb[83]
port 434 nsew signal tristate
rlabel metal2 s 284206 163200 284262 164400 6 la_oenb[84]
port 435 nsew signal tristate
rlabel metal2 s 287518 163200 287574 164400 6 la_oenb[85]
port 436 nsew signal tristate
rlabel metal2 s 290922 163200 290978 164400 6 la_oenb[86]
port 437 nsew signal tristate
rlabel metal2 s 294234 163200 294290 164400 6 la_oenb[87]
port 438 nsew signal tristate
rlabel metal2 s 297638 163200 297694 164400 6 la_oenb[88]
port 439 nsew signal tristate
rlabel metal2 s 300950 163200 301006 164400 6 la_oenb[89]
port 440 nsew signal tristate
rlabel metal2 s 28906 163200 28962 164400 6 la_oenb[8]
port 441 nsew signal tristate
rlabel metal2 s 304354 163200 304410 164400 6 la_oenb[90]
port 442 nsew signal tristate
rlabel metal2 s 307666 163200 307722 164400 6 la_oenb[91]
port 443 nsew signal tristate
rlabel metal2 s 311070 163200 311126 164400 6 la_oenb[92]
port 444 nsew signal tristate
rlabel metal2 s 314382 163200 314438 164400 6 la_oenb[93]
port 445 nsew signal tristate
rlabel metal2 s 317786 163200 317842 164400 6 la_oenb[94]
port 446 nsew signal tristate
rlabel metal2 s 321098 163200 321154 164400 6 la_oenb[95]
port 447 nsew signal tristate
rlabel metal2 s 324502 163200 324558 164400 6 la_oenb[96]
port 448 nsew signal tristate
rlabel metal2 s 327906 163200 327962 164400 6 la_oenb[97]
port 449 nsew signal tristate
rlabel metal2 s 331218 163200 331274 164400 6 la_oenb[98]
port 450 nsew signal tristate
rlabel metal2 s 334622 163200 334678 164400 6 la_oenb[99]
port 451 nsew signal tristate
rlabel metal2 s 32218 163200 32274 164400 6 la_oenb[9]
port 452 nsew signal tristate
rlabel metal2 s 2870 163200 2926 164400 6 la_output[0]
port 453 nsew signal tristate
rlabel metal2 s 338762 163200 338818 164400 6 la_output[100]
port 454 nsew signal tristate
rlabel metal2 s 342166 163200 342222 164400 6 la_output[101]
port 455 nsew signal tristate
rlabel metal2 s 345478 163200 345534 164400 6 la_output[102]
port 456 nsew signal tristate
rlabel metal2 s 348882 163200 348938 164400 6 la_output[103]
port 457 nsew signal tristate
rlabel metal2 s 352194 163200 352250 164400 6 la_output[104]
port 458 nsew signal tristate
rlabel metal2 s 355598 163200 355654 164400 6 la_output[105]
port 459 nsew signal tristate
rlabel metal2 s 358910 163200 358966 164400 6 la_output[106]
port 460 nsew signal tristate
rlabel metal2 s 362314 163200 362370 164400 6 la_output[107]
port 461 nsew signal tristate
rlabel metal2 s 365626 163200 365682 164400 6 la_output[108]
port 462 nsew signal tristate
rlabel metal2 s 369030 163200 369086 164400 6 la_output[109]
port 463 nsew signal tristate
rlabel metal2 s 36450 163200 36506 164400 6 la_output[10]
port 464 nsew signal tristate
rlabel metal2 s 372342 163200 372398 164400 6 la_output[110]
port 465 nsew signal tristate
rlabel metal2 s 375746 163200 375802 164400 6 la_output[111]
port 466 nsew signal tristate
rlabel metal2 s 379058 163200 379114 164400 6 la_output[112]
port 467 nsew signal tristate
rlabel metal2 s 382462 163200 382518 164400 6 la_output[113]
port 468 nsew signal tristate
rlabel metal2 s 385774 163200 385830 164400 6 la_output[114]
port 469 nsew signal tristate
rlabel metal2 s 389178 163200 389234 164400 6 la_output[115]
port 470 nsew signal tristate
rlabel metal2 s 392490 163200 392546 164400 6 la_output[116]
port 471 nsew signal tristate
rlabel metal2 s 395894 163200 395950 164400 6 la_output[117]
port 472 nsew signal tristate
rlabel metal2 s 399206 163200 399262 164400 6 la_output[118]
port 473 nsew signal tristate
rlabel metal2 s 402610 163200 402666 164400 6 la_output[119]
port 474 nsew signal tristate
rlabel metal2 s 39854 163200 39910 164400 6 la_output[11]
port 475 nsew signal tristate
rlabel metal2 s 405922 163200 405978 164400 6 la_output[120]
port 476 nsew signal tristate
rlabel metal2 s 409326 163200 409382 164400 6 la_output[121]
port 477 nsew signal tristate
rlabel metal2 s 412638 163200 412694 164400 6 la_output[122]
port 478 nsew signal tristate
rlabel metal2 s 416042 163200 416098 164400 6 la_output[123]
port 479 nsew signal tristate
rlabel metal2 s 419354 163200 419410 164400 6 la_output[124]
port 480 nsew signal tristate
rlabel metal2 s 422758 163200 422814 164400 6 la_output[125]
port 481 nsew signal tristate
rlabel metal2 s 426162 163200 426218 164400 6 la_output[126]
port 482 nsew signal tristate
rlabel metal2 s 429474 163200 429530 164400 6 la_output[127]
port 483 nsew signal tristate
rlabel metal2 s 43166 163200 43222 164400 6 la_output[12]
port 484 nsew signal tristate
rlabel metal2 s 46570 163200 46626 164400 6 la_output[13]
port 485 nsew signal tristate
rlabel metal2 s 49882 163200 49938 164400 6 la_output[14]
port 486 nsew signal tristate
rlabel metal2 s 53286 163200 53342 164400 6 la_output[15]
port 487 nsew signal tristate
rlabel metal2 s 56598 163200 56654 164400 6 la_output[16]
port 488 nsew signal tristate
rlabel metal2 s 60002 163200 60058 164400 6 la_output[17]
port 489 nsew signal tristate
rlabel metal2 s 63314 163200 63370 164400 6 la_output[18]
port 490 nsew signal tristate
rlabel metal2 s 66718 163200 66774 164400 6 la_output[19]
port 491 nsew signal tristate
rlabel metal2 s 6182 163200 6238 164400 6 la_output[1]
port 492 nsew signal tristate
rlabel metal2 s 70030 163200 70086 164400 6 la_output[20]
port 493 nsew signal tristate
rlabel metal2 s 73434 163200 73490 164400 6 la_output[21]
port 494 nsew signal tristate
rlabel metal2 s 76746 163200 76802 164400 6 la_output[22]
port 495 nsew signal tristate
rlabel metal2 s 80150 163200 80206 164400 6 la_output[23]
port 496 nsew signal tristate
rlabel metal2 s 83462 163200 83518 164400 6 la_output[24]
port 497 nsew signal tristate
rlabel metal2 s 86866 163200 86922 164400 6 la_output[25]
port 498 nsew signal tristate
rlabel metal2 s 90178 163200 90234 164400 6 la_output[26]
port 499 nsew signal tristate
rlabel metal2 s 93582 163200 93638 164400 6 la_output[27]
port 500 nsew signal tristate
rlabel metal2 s 96894 163200 96950 164400 6 la_output[28]
port 501 nsew signal tristate
rlabel metal2 s 100298 163200 100354 164400 6 la_output[29]
port 502 nsew signal tristate
rlabel metal2 s 9586 163200 9642 164400 6 la_output[2]
port 503 nsew signal tristate
rlabel metal2 s 103610 163200 103666 164400 6 la_output[30]
port 504 nsew signal tristate
rlabel metal2 s 107014 163200 107070 164400 6 la_output[31]
port 505 nsew signal tristate
rlabel metal2 s 110326 163200 110382 164400 6 la_output[32]
port 506 nsew signal tristate
rlabel metal2 s 113730 163200 113786 164400 6 la_output[33]
port 507 nsew signal tristate
rlabel metal2 s 117042 163200 117098 164400 6 la_output[34]
port 508 nsew signal tristate
rlabel metal2 s 120446 163200 120502 164400 6 la_output[35]
port 509 nsew signal tristate
rlabel metal2 s 123758 163200 123814 164400 6 la_output[36]
port 510 nsew signal tristate
rlabel metal2 s 127162 163200 127218 164400 6 la_output[37]
port 511 nsew signal tristate
rlabel metal2 s 130474 163200 130530 164400 6 la_output[38]
port 512 nsew signal tristate
rlabel metal2 s 133878 163200 133934 164400 6 la_output[39]
port 513 nsew signal tristate
rlabel metal2 s 12898 163200 12954 164400 6 la_output[3]
port 514 nsew signal tristate
rlabel metal2 s 137190 163200 137246 164400 6 la_output[40]
port 515 nsew signal tristate
rlabel metal2 s 140594 163200 140650 164400 6 la_output[41]
port 516 nsew signal tristate
rlabel metal2 s 143906 163200 143962 164400 6 la_output[42]
port 517 nsew signal tristate
rlabel metal2 s 147310 163200 147366 164400 6 la_output[43]
port 518 nsew signal tristate
rlabel metal2 s 150622 163200 150678 164400 6 la_output[44]
port 519 nsew signal tristate
rlabel metal2 s 154026 163200 154082 164400 6 la_output[45]
port 520 nsew signal tristate
rlabel metal2 s 157338 163200 157394 164400 6 la_output[46]
port 521 nsew signal tristate
rlabel metal2 s 160742 163200 160798 164400 6 la_output[47]
port 522 nsew signal tristate
rlabel metal2 s 164146 163200 164202 164400 6 la_output[48]
port 523 nsew signal tristate
rlabel metal2 s 167458 163200 167514 164400 6 la_output[49]
port 524 nsew signal tristate
rlabel metal2 s 16302 163200 16358 164400 6 la_output[4]
port 525 nsew signal tristate
rlabel metal2 s 170862 163200 170918 164400 6 la_output[50]
port 526 nsew signal tristate
rlabel metal2 s 174174 163200 174230 164400 6 la_output[51]
port 527 nsew signal tristate
rlabel metal2 s 177578 163200 177634 164400 6 la_output[52]
port 528 nsew signal tristate
rlabel metal2 s 180890 163200 180946 164400 6 la_output[53]
port 529 nsew signal tristate
rlabel metal2 s 184294 163200 184350 164400 6 la_output[54]
port 530 nsew signal tristate
rlabel metal2 s 187606 163200 187662 164400 6 la_output[55]
port 531 nsew signal tristate
rlabel metal2 s 191010 163200 191066 164400 6 la_output[56]
port 532 nsew signal tristate
rlabel metal2 s 194322 163200 194378 164400 6 la_output[57]
port 533 nsew signal tristate
rlabel metal2 s 197726 163200 197782 164400 6 la_output[58]
port 534 nsew signal tristate
rlabel metal2 s 201038 163200 201094 164400 6 la_output[59]
port 535 nsew signal tristate
rlabel metal2 s 19614 163200 19670 164400 6 la_output[5]
port 536 nsew signal tristate
rlabel metal2 s 204442 163200 204498 164400 6 la_output[60]
port 537 nsew signal tristate
rlabel metal2 s 207754 163200 207810 164400 6 la_output[61]
port 538 nsew signal tristate
rlabel metal2 s 211158 163200 211214 164400 6 la_output[62]
port 539 nsew signal tristate
rlabel metal2 s 214470 163200 214526 164400 6 la_output[63]
port 540 nsew signal tristate
rlabel metal2 s 217874 163200 217930 164400 6 la_output[64]
port 541 nsew signal tristate
rlabel metal2 s 221186 163200 221242 164400 6 la_output[65]
port 542 nsew signal tristate
rlabel metal2 s 224590 163200 224646 164400 6 la_output[66]
port 543 nsew signal tristate
rlabel metal2 s 227902 163200 227958 164400 6 la_output[67]
port 544 nsew signal tristate
rlabel metal2 s 231306 163200 231362 164400 6 la_output[68]
port 545 nsew signal tristate
rlabel metal2 s 234618 163200 234674 164400 6 la_output[69]
port 546 nsew signal tristate
rlabel metal2 s 23018 163200 23074 164400 6 la_output[6]
port 547 nsew signal tristate
rlabel metal2 s 238022 163200 238078 164400 6 la_output[70]
port 548 nsew signal tristate
rlabel metal2 s 241334 163200 241390 164400 6 la_output[71]
port 549 nsew signal tristate
rlabel metal2 s 244738 163200 244794 164400 6 la_output[72]
port 550 nsew signal tristate
rlabel metal2 s 248050 163200 248106 164400 6 la_output[73]
port 551 nsew signal tristate
rlabel metal2 s 251454 163200 251510 164400 6 la_output[74]
port 552 nsew signal tristate
rlabel metal2 s 254766 163200 254822 164400 6 la_output[75]
port 553 nsew signal tristate
rlabel metal2 s 258170 163200 258226 164400 6 la_output[76]
port 554 nsew signal tristate
rlabel metal2 s 261482 163200 261538 164400 6 la_output[77]
port 555 nsew signal tristate
rlabel metal2 s 264886 163200 264942 164400 6 la_output[78]
port 556 nsew signal tristate
rlabel metal2 s 268198 163200 268254 164400 6 la_output[79]
port 557 nsew signal tristate
rlabel metal2 s 26330 163200 26386 164400 6 la_output[7]
port 558 nsew signal tristate
rlabel metal2 s 271602 163200 271658 164400 6 la_output[80]
port 559 nsew signal tristate
rlabel metal2 s 274914 163200 274970 164400 6 la_output[81]
port 560 nsew signal tristate
rlabel metal2 s 278318 163200 278374 164400 6 la_output[82]
port 561 nsew signal tristate
rlabel metal2 s 281630 163200 281686 164400 6 la_output[83]
port 562 nsew signal tristate
rlabel metal2 s 285034 163200 285090 164400 6 la_output[84]
port 563 nsew signal tristate
rlabel metal2 s 288346 163200 288402 164400 6 la_output[85]
port 564 nsew signal tristate
rlabel metal2 s 291750 163200 291806 164400 6 la_output[86]
port 565 nsew signal tristate
rlabel metal2 s 295154 163200 295210 164400 6 la_output[87]
port 566 nsew signal tristate
rlabel metal2 s 298466 163200 298522 164400 6 la_output[88]
port 567 nsew signal tristate
rlabel metal2 s 301870 163200 301926 164400 6 la_output[89]
port 568 nsew signal tristate
rlabel metal2 s 29734 163200 29790 164400 6 la_output[8]
port 569 nsew signal tristate
rlabel metal2 s 305182 163200 305238 164400 6 la_output[90]
port 570 nsew signal tristate
rlabel metal2 s 308586 163200 308642 164400 6 la_output[91]
port 571 nsew signal tristate
rlabel metal2 s 311898 163200 311954 164400 6 la_output[92]
port 572 nsew signal tristate
rlabel metal2 s 315302 163200 315358 164400 6 la_output[93]
port 573 nsew signal tristate
rlabel metal2 s 318614 163200 318670 164400 6 la_output[94]
port 574 nsew signal tristate
rlabel metal2 s 322018 163200 322074 164400 6 la_output[95]
port 575 nsew signal tristate
rlabel metal2 s 325330 163200 325386 164400 6 la_output[96]
port 576 nsew signal tristate
rlabel metal2 s 328734 163200 328790 164400 6 la_output[97]
port 577 nsew signal tristate
rlabel metal2 s 332046 163200 332102 164400 6 la_output[98]
port 578 nsew signal tristate
rlabel metal2 s 335450 163200 335506 164400 6 la_output[99]
port 579 nsew signal tristate
rlabel metal2 s 33138 163200 33194 164400 6 la_output[9]
port 580 nsew signal tristate
rlabel metal2 s 430302 163200 430358 164400 6 mprj_ack_i
port 581 nsew signal input
rlabel metal2 s 434534 163200 434590 164400 6 mprj_adr_o[0]
port 582 nsew signal tristate
rlabel metal2 s 463054 163200 463110 164400 6 mprj_adr_o[10]
port 583 nsew signal tristate
rlabel metal2 s 465630 163200 465686 164400 6 mprj_adr_o[11]
port 584 nsew signal tristate
rlabel metal2 s 468114 163200 468170 164400 6 mprj_adr_o[12]
port 585 nsew signal tristate
rlabel metal2 s 470598 163200 470654 164400 6 mprj_adr_o[13]
port 586 nsew signal tristate
rlabel metal2 s 473174 163200 473230 164400 6 mprj_adr_o[14]
port 587 nsew signal tristate
rlabel metal2 s 475658 163200 475714 164400 6 mprj_adr_o[15]
port 588 nsew signal tristate
rlabel metal2 s 478142 163200 478198 164400 6 mprj_adr_o[16]
port 589 nsew signal tristate
rlabel metal2 s 480718 163200 480774 164400 6 mprj_adr_o[17]
port 590 nsew signal tristate
rlabel metal2 s 483202 163200 483258 164400 6 mprj_adr_o[18]
port 591 nsew signal tristate
rlabel metal2 s 485778 163200 485834 164400 6 mprj_adr_o[19]
port 592 nsew signal tristate
rlabel metal2 s 437846 163200 437902 164400 6 mprj_adr_o[1]
port 593 nsew signal tristate
rlabel metal2 s 488262 163200 488318 164400 6 mprj_adr_o[20]
port 594 nsew signal tristate
rlabel metal2 s 490746 163200 490802 164400 6 mprj_adr_o[21]
port 595 nsew signal tristate
rlabel metal2 s 493322 163200 493378 164400 6 mprj_adr_o[22]
port 596 nsew signal tristate
rlabel metal2 s 495806 163200 495862 164400 6 mprj_adr_o[23]
port 597 nsew signal tristate
rlabel metal2 s 498382 163200 498438 164400 6 mprj_adr_o[24]
port 598 nsew signal tristate
rlabel metal2 s 500866 163200 500922 164400 6 mprj_adr_o[25]
port 599 nsew signal tristate
rlabel metal2 s 503350 163200 503406 164400 6 mprj_adr_o[26]
port 600 nsew signal tristate
rlabel metal2 s 505926 163200 505982 164400 6 mprj_adr_o[27]
port 601 nsew signal tristate
rlabel metal2 s 508410 163200 508466 164400 6 mprj_adr_o[28]
port 602 nsew signal tristate
rlabel metal2 s 510894 163200 510950 164400 6 mprj_adr_o[29]
port 603 nsew signal tristate
rlabel metal2 s 441250 163200 441306 164400 6 mprj_adr_o[2]
port 604 nsew signal tristate
rlabel metal2 s 513470 163200 513526 164400 6 mprj_adr_o[30]
port 605 nsew signal tristate
rlabel metal2 s 515954 163200 516010 164400 6 mprj_adr_o[31]
port 606 nsew signal tristate
rlabel metal2 s 444562 163200 444618 164400 6 mprj_adr_o[3]
port 607 nsew signal tristate
rlabel metal2 s 447966 163200 448022 164400 6 mprj_adr_o[4]
port 608 nsew signal tristate
rlabel metal2 s 450450 163200 450506 164400 6 mprj_adr_o[5]
port 609 nsew signal tristate
rlabel metal2 s 453026 163200 453082 164400 6 mprj_adr_o[6]
port 610 nsew signal tristate
rlabel metal2 s 455510 163200 455566 164400 6 mprj_adr_o[7]
port 611 nsew signal tristate
rlabel metal2 s 457994 163200 458050 164400 6 mprj_adr_o[8]
port 612 nsew signal tristate
rlabel metal2 s 460570 163200 460626 164400 6 mprj_adr_o[9]
port 613 nsew signal tristate
rlabel metal2 s 431130 163200 431186 164400 6 mprj_cyc_o
port 614 nsew signal tristate
rlabel metal2 s 435362 163200 435418 164400 6 mprj_dat_i[0]
port 615 nsew signal input
rlabel metal2 s 463882 163200 463938 164400 6 mprj_dat_i[10]
port 616 nsew signal input
rlabel metal2 s 466458 163200 466514 164400 6 mprj_dat_i[11]
port 617 nsew signal input
rlabel metal2 s 468942 163200 468998 164400 6 mprj_dat_i[12]
port 618 nsew signal input
rlabel metal2 s 471426 163200 471482 164400 6 mprj_dat_i[13]
port 619 nsew signal input
rlabel metal2 s 474002 163200 474058 164400 6 mprj_dat_i[14]
port 620 nsew signal input
rlabel metal2 s 476486 163200 476542 164400 6 mprj_dat_i[15]
port 621 nsew signal input
rlabel metal2 s 479062 163200 479118 164400 6 mprj_dat_i[16]
port 622 nsew signal input
rlabel metal2 s 481546 163200 481602 164400 6 mprj_dat_i[17]
port 623 nsew signal input
rlabel metal2 s 484030 163200 484086 164400 6 mprj_dat_i[18]
port 624 nsew signal input
rlabel metal2 s 486606 163200 486662 164400 6 mprj_dat_i[19]
port 625 nsew signal input
rlabel metal2 s 438674 163200 438730 164400 6 mprj_dat_i[1]
port 626 nsew signal input
rlabel metal2 s 489090 163200 489146 164400 6 mprj_dat_i[20]
port 627 nsew signal input
rlabel metal2 s 491666 163200 491722 164400 6 mprj_dat_i[21]
port 628 nsew signal input
rlabel metal2 s 494150 163200 494206 164400 6 mprj_dat_i[22]
port 629 nsew signal input
rlabel metal2 s 496634 163200 496690 164400 6 mprj_dat_i[23]
port 630 nsew signal input
rlabel metal2 s 499210 163200 499266 164400 6 mprj_dat_i[24]
port 631 nsew signal input
rlabel metal2 s 501694 163200 501750 164400 6 mprj_dat_i[25]
port 632 nsew signal input
rlabel metal2 s 504178 163200 504234 164400 6 mprj_dat_i[26]
port 633 nsew signal input
rlabel metal2 s 506754 163200 506810 164400 6 mprj_dat_i[27]
port 634 nsew signal input
rlabel metal2 s 509238 163200 509294 164400 6 mprj_dat_i[28]
port 635 nsew signal input
rlabel metal2 s 511814 163200 511870 164400 6 mprj_dat_i[29]
port 636 nsew signal input
rlabel metal2 s 442078 163200 442134 164400 6 mprj_dat_i[2]
port 637 nsew signal input
rlabel metal2 s 514298 163200 514354 164400 6 mprj_dat_i[30]
port 638 nsew signal input
rlabel metal2 s 516782 163200 516838 164400 6 mprj_dat_i[31]
port 639 nsew signal input
rlabel metal2 s 445390 163200 445446 164400 6 mprj_dat_i[3]
port 640 nsew signal input
rlabel metal2 s 448794 163200 448850 164400 6 mprj_dat_i[4]
port 641 nsew signal input
rlabel metal2 s 451278 163200 451334 164400 6 mprj_dat_i[5]
port 642 nsew signal input
rlabel metal2 s 453854 163200 453910 164400 6 mprj_dat_i[6]
port 643 nsew signal input
rlabel metal2 s 456338 163200 456394 164400 6 mprj_dat_i[7]
port 644 nsew signal input
rlabel metal2 s 458914 163200 458970 164400 6 mprj_dat_i[8]
port 645 nsew signal input
rlabel metal2 s 461398 163200 461454 164400 6 mprj_dat_i[9]
port 646 nsew signal input
rlabel metal2 s 436190 163200 436246 164400 6 mprj_dat_o[0]
port 647 nsew signal tristate
rlabel metal2 s 464710 163200 464766 164400 6 mprj_dat_o[10]
port 648 nsew signal tristate
rlabel metal2 s 467286 163200 467342 164400 6 mprj_dat_o[11]
port 649 nsew signal tristate
rlabel metal2 s 469770 163200 469826 164400 6 mprj_dat_o[12]
port 650 nsew signal tristate
rlabel metal2 s 472346 163200 472402 164400 6 mprj_dat_o[13]
port 651 nsew signal tristate
rlabel metal2 s 474830 163200 474886 164400 6 mprj_dat_o[14]
port 652 nsew signal tristate
rlabel metal2 s 477314 163200 477370 164400 6 mprj_dat_o[15]
port 653 nsew signal tristate
rlabel metal2 s 479890 163200 479946 164400 6 mprj_dat_o[16]
port 654 nsew signal tristate
rlabel metal2 s 482374 163200 482430 164400 6 mprj_dat_o[17]
port 655 nsew signal tristate
rlabel metal2 s 484858 163200 484914 164400 6 mprj_dat_o[18]
port 656 nsew signal tristate
rlabel metal2 s 487434 163200 487490 164400 6 mprj_dat_o[19]
port 657 nsew signal tristate
rlabel metal2 s 439594 163200 439650 164400 6 mprj_dat_o[1]
port 658 nsew signal tristate
rlabel metal2 s 489918 163200 489974 164400 6 mprj_dat_o[20]
port 659 nsew signal tristate
rlabel metal2 s 492494 163200 492550 164400 6 mprj_dat_o[21]
port 660 nsew signal tristate
rlabel metal2 s 494978 163200 495034 164400 6 mprj_dat_o[22]
port 661 nsew signal tristate
rlabel metal2 s 497462 163200 497518 164400 6 mprj_dat_o[23]
port 662 nsew signal tristate
rlabel metal2 s 500038 163200 500094 164400 6 mprj_dat_o[24]
port 663 nsew signal tristate
rlabel metal2 s 502522 163200 502578 164400 6 mprj_dat_o[25]
port 664 nsew signal tristate
rlabel metal2 s 505098 163200 505154 164400 6 mprj_dat_o[26]
port 665 nsew signal tristate
rlabel metal2 s 507582 163200 507638 164400 6 mprj_dat_o[27]
port 666 nsew signal tristate
rlabel metal2 s 510066 163200 510122 164400 6 mprj_dat_o[28]
port 667 nsew signal tristate
rlabel metal2 s 512642 163200 512698 164400 6 mprj_dat_o[29]
port 668 nsew signal tristate
rlabel metal2 s 442906 163200 442962 164400 6 mprj_dat_o[2]
port 669 nsew signal tristate
rlabel metal2 s 515126 163200 515182 164400 6 mprj_dat_o[30]
port 670 nsew signal tristate
rlabel metal2 s 517610 163200 517666 164400 6 mprj_dat_o[31]
port 671 nsew signal tristate
rlabel metal2 s 446310 163200 446366 164400 6 mprj_dat_o[3]
port 672 nsew signal tristate
rlabel metal2 s 449622 163200 449678 164400 6 mprj_dat_o[4]
port 673 nsew signal tristate
rlabel metal2 s 452106 163200 452162 164400 6 mprj_dat_o[5]
port 674 nsew signal tristate
rlabel metal2 s 454682 163200 454738 164400 6 mprj_dat_o[6]
port 675 nsew signal tristate
rlabel metal2 s 457166 163200 457222 164400 6 mprj_dat_o[7]
port 676 nsew signal tristate
rlabel metal2 s 459742 163200 459798 164400 6 mprj_dat_o[8]
port 677 nsew signal tristate
rlabel metal2 s 462226 163200 462282 164400 6 mprj_dat_o[9]
port 678 nsew signal tristate
rlabel metal2 s 437018 163200 437074 164400 6 mprj_sel_o[0]
port 679 nsew signal tristate
rlabel metal2 s 440422 163200 440478 164400 6 mprj_sel_o[1]
port 680 nsew signal tristate
rlabel metal2 s 443734 163200 443790 164400 6 mprj_sel_o[2]
port 681 nsew signal tristate
rlabel metal2 s 447138 163200 447194 164400 6 mprj_sel_o[3]
port 682 nsew signal tristate
rlabel metal2 s 431958 163200 432014 164400 6 mprj_stb_o
port 683 nsew signal tristate
rlabel metal2 s 432878 163200 432934 164400 6 mprj_wb_iena
port 684 nsew signal tristate
rlabel metal2 s 433706 163200 433762 164400 6 mprj_we_o
port 685 nsew signal tristate
rlabel metal3 s 523200 90176 524400 90296 6 qspi_enabled
port 686 nsew signal tristate
rlabel metal3 s 523200 84192 524400 84312 6 ser_rx
port 687 nsew signal input
rlabel metal3 s 523200 85688 524400 85808 6 ser_tx
port 688 nsew signal tristate
rlabel metal3 s 523200 81064 524400 81184 6 spi_csb
port 689 nsew signal tristate
rlabel metal3 s 523200 87184 524400 87304 6 spi_enabled
port 690 nsew signal tristate
rlabel metal3 s 523200 79568 524400 79688 6 spi_sck
port 691 nsew signal tristate
rlabel metal3 s 523200 82696 524400 82816 6 spi_sdi
port 692 nsew signal input
rlabel metal3 s 523200 78072 524400 78192 6 spi_sdo
port 693 nsew signal tristate
rlabel metal3 s 523200 76576 524400 76696 6 spi_sdoenb
port 694 nsew signal tristate
rlabel metal3 s 523200 2184 524400 2304 6 sram_ro_addr[0]
port 695 nsew signal input
rlabel metal3 s 523200 3680 524400 3800 6 sram_ro_addr[1]
port 696 nsew signal input
rlabel metal3 s 523200 5176 524400 5296 6 sram_ro_addr[2]
port 697 nsew signal input
rlabel metal3 s 523200 6672 524400 6792 6 sram_ro_addr[3]
port 698 nsew signal input
rlabel metal3 s 523200 8168 524400 8288 6 sram_ro_addr[4]
port 699 nsew signal input
rlabel metal3 s 523200 9800 524400 9920 6 sram_ro_addr[5]
port 700 nsew signal input
rlabel metal3 s 523200 11296 524400 11416 6 sram_ro_addr[6]
port 701 nsew signal input
rlabel metal3 s 523200 12792 524400 12912 6 sram_ro_addr[7]
port 702 nsew signal input
rlabel metal3 s 523200 14288 524400 14408 6 sram_ro_clk
port 703 nsew signal input
rlabel metal3 s 523200 688 524400 808 6 sram_ro_csb
port 704 nsew signal input
rlabel metal3 s 523200 15784 524400 15904 6 sram_ro_data[0]
port 705 nsew signal tristate
rlabel metal3 s 523200 31016 524400 31136 6 sram_ro_data[10]
port 706 nsew signal tristate
rlabel metal3 s 523200 32512 524400 32632 6 sram_ro_data[11]
port 707 nsew signal tristate
rlabel metal3 s 523200 34008 524400 34128 6 sram_ro_data[12]
port 708 nsew signal tristate
rlabel metal3 s 523200 35504 524400 35624 6 sram_ro_data[13]
port 709 nsew signal tristate
rlabel metal3 s 523200 37136 524400 37256 6 sram_ro_data[14]
port 710 nsew signal tristate
rlabel metal3 s 523200 38632 524400 38752 6 sram_ro_data[15]
port 711 nsew signal tristate
rlabel metal3 s 523200 40128 524400 40248 6 sram_ro_data[16]
port 712 nsew signal tristate
rlabel metal3 s 523200 41624 524400 41744 6 sram_ro_data[17]
port 713 nsew signal tristate
rlabel metal3 s 523200 43120 524400 43240 6 sram_ro_data[18]
port 714 nsew signal tristate
rlabel metal3 s 523200 44616 524400 44736 6 sram_ro_data[19]
port 715 nsew signal tristate
rlabel metal3 s 523200 17280 524400 17400 6 sram_ro_data[1]
port 716 nsew signal tristate
rlabel metal3 s 523200 46248 524400 46368 6 sram_ro_data[20]
port 717 nsew signal tristate
rlabel metal3 s 523200 47744 524400 47864 6 sram_ro_data[21]
port 718 nsew signal tristate
rlabel metal3 s 523200 49240 524400 49360 6 sram_ro_data[22]
port 719 nsew signal tristate
rlabel metal3 s 523200 50736 524400 50856 6 sram_ro_data[23]
port 720 nsew signal tristate
rlabel metal3 s 523200 52232 524400 52352 6 sram_ro_data[24]
port 721 nsew signal tristate
rlabel metal3 s 523200 53728 524400 53848 6 sram_ro_data[25]
port 722 nsew signal tristate
rlabel metal3 s 523200 55360 524400 55480 6 sram_ro_data[26]
port 723 nsew signal tristate
rlabel metal3 s 523200 56856 524400 56976 6 sram_ro_data[27]
port 724 nsew signal tristate
rlabel metal3 s 523200 58352 524400 58472 6 sram_ro_data[28]
port 725 nsew signal tristate
rlabel metal3 s 523200 59848 524400 59968 6 sram_ro_data[29]
port 726 nsew signal tristate
rlabel metal3 s 523200 18912 524400 19032 6 sram_ro_data[2]
port 727 nsew signal tristate
rlabel metal3 s 523200 61344 524400 61464 6 sram_ro_data[30]
port 728 nsew signal tristate
rlabel metal3 s 523200 62840 524400 62960 6 sram_ro_data[31]
port 729 nsew signal tristate
rlabel metal3 s 523200 20408 524400 20528 6 sram_ro_data[3]
port 730 nsew signal tristate
rlabel metal3 s 523200 21904 524400 22024 6 sram_ro_data[4]
port 731 nsew signal tristate
rlabel metal3 s 523200 23400 524400 23520 6 sram_ro_data[5]
port 732 nsew signal tristate
rlabel metal3 s 523200 24896 524400 25016 6 sram_ro_data[6]
port 733 nsew signal tristate
rlabel metal3 s 523200 26392 524400 26512 6 sram_ro_data[7]
port 734 nsew signal tristate
rlabel metal3 s 523200 28024 524400 28144 6 sram_ro_data[8]
port 735 nsew signal tristate
rlabel metal3 s 523200 29520 524400 29640 6 sram_ro_data[9]
port 736 nsew signal tristate
rlabel metal3 s 523200 70456 524400 70576 6 trap
port 737 nsew signal tristate
rlabel metal3 s 523200 88680 524400 88800 6 uart_enabled
port 738 nsew signal tristate
rlabel metal2 s 518530 163200 518586 164400 6 user_irq_ena[0]
port 739 nsew signal tristate
rlabel metal2 s 519358 163200 519414 164400 6 user_irq_ena[1]
port 740 nsew signal tristate
rlabel metal2 s 520186 163200 520242 164400 6 user_irq_ena[2]
port 741 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 524000 164000
<< end >>
