VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM128
  CLASS BLOCK ;
  FOREIGN RAM128 ;
  ORIGIN 0.000 0.000 ;
  SIZE 402.040 BY 394.400 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.040 180.240 402.040 180.840 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.040 212.880 402.040 213.480 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.040 245.520 402.040 246.120 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.040 278.160 402.040 278.760 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.040 310.800 402.040 311.400 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.040 343.440 402.040 344.040 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.040 376.080 402.040 376.680 ;
    END
  END A0[6]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 2.000 197.160 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 0.000 294.310 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 0.000 381.250 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 2.000 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 2.000 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 2.000 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 2.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 392.400 8.650 394.400 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 392.400 132.850 394.400 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 392.400 145.270 394.400 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 392.400 157.690 394.400 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 392.400 170.110 394.400 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 392.400 182.530 394.400 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 392.400 194.950 394.400 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 392.400 207.370 394.400 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 392.400 219.790 394.400 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 392.400 232.210 394.400 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 392.400 244.630 394.400 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 392.400 21.070 394.400 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 392.400 257.050 394.400 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 392.400 269.470 394.400 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 392.400 281.890 394.400 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 392.400 294.310 394.400 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 392.400 306.730 394.400 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 392.400 319.150 394.400 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 392.400 331.570 394.400 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 392.400 343.990 394.400 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 392.400 356.410 394.400 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 392.400 368.830 394.400 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 392.400 33.490 394.400 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 392.400 381.250 394.400 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 392.400 393.670 394.400 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 392.400 45.910 394.400 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 392.400 58.330 394.400 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 392.400 70.750 394.400 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 392.400 83.170 394.400 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 392.400 95.590 394.400 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 392.400 108.010 394.400 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 392.400 120.430 394.400 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.040 17.040 402.040 17.640 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 391.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.680 2.480 250.280 391.920 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 391.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 391.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 391.920 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.040 49.680 402.040 50.280 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.040 82.320 402.040 82.920 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.040 114.960 402.040 115.560 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.040 147.600 402.040 148.200 ;
    END
  END WE0[3]
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 399.280 391.765 ;
      LAYER met1 ;
        RECT 2.760 0.040 401.970 394.360 ;
      LAYER met2 ;
        RECT 3.310 392.120 8.090 394.390 ;
        RECT 8.930 392.120 20.510 394.390 ;
        RECT 21.350 392.120 32.930 394.390 ;
        RECT 33.770 392.120 45.350 394.390 ;
        RECT 46.190 392.120 57.770 394.390 ;
        RECT 58.610 392.120 70.190 394.390 ;
        RECT 71.030 392.120 82.610 394.390 ;
        RECT 83.450 392.120 95.030 394.390 ;
        RECT 95.870 392.120 107.450 394.390 ;
        RECT 108.290 392.120 119.870 394.390 ;
        RECT 120.710 392.120 132.290 394.390 ;
        RECT 133.130 392.120 144.710 394.390 ;
        RECT 145.550 392.120 157.130 394.390 ;
        RECT 157.970 392.120 169.550 394.390 ;
        RECT 170.390 392.120 181.970 394.390 ;
        RECT 182.810 392.120 194.390 394.390 ;
        RECT 195.230 392.120 206.810 394.390 ;
        RECT 207.650 392.120 219.230 394.390 ;
        RECT 220.070 392.120 231.650 394.390 ;
        RECT 232.490 392.120 244.070 394.390 ;
        RECT 244.910 392.120 256.490 394.390 ;
        RECT 257.330 392.120 268.910 394.390 ;
        RECT 269.750 392.120 281.330 394.390 ;
        RECT 282.170 392.120 293.750 394.390 ;
        RECT 294.590 392.120 306.170 394.390 ;
        RECT 307.010 392.120 318.590 394.390 ;
        RECT 319.430 392.120 331.010 394.390 ;
        RECT 331.850 392.120 343.430 394.390 ;
        RECT 344.270 392.120 355.850 394.390 ;
        RECT 356.690 392.120 368.270 394.390 ;
        RECT 369.110 392.120 380.690 394.390 ;
        RECT 381.530 392.120 393.110 394.390 ;
        RECT 393.950 392.120 401.940 394.390 ;
        RECT 3.310 2.280 401.940 392.120 ;
        RECT 3.310 0.010 8.090 2.280 ;
        RECT 8.930 0.010 20.510 2.280 ;
        RECT 21.350 0.010 32.930 2.280 ;
        RECT 33.770 0.010 45.350 2.280 ;
        RECT 46.190 0.010 57.770 2.280 ;
        RECT 58.610 0.010 70.190 2.280 ;
        RECT 71.030 0.010 82.610 2.280 ;
        RECT 83.450 0.010 95.030 2.280 ;
        RECT 95.870 0.010 107.450 2.280 ;
        RECT 108.290 0.010 119.870 2.280 ;
        RECT 120.710 0.010 132.290 2.280 ;
        RECT 133.130 0.010 144.710 2.280 ;
        RECT 145.550 0.010 157.130 2.280 ;
        RECT 157.970 0.010 169.550 2.280 ;
        RECT 170.390 0.010 181.970 2.280 ;
        RECT 182.810 0.010 194.390 2.280 ;
        RECT 195.230 0.010 206.810 2.280 ;
        RECT 207.650 0.010 219.230 2.280 ;
        RECT 220.070 0.010 231.650 2.280 ;
        RECT 232.490 0.010 244.070 2.280 ;
        RECT 244.910 0.010 256.490 2.280 ;
        RECT 257.330 0.010 268.910 2.280 ;
        RECT 269.750 0.010 281.330 2.280 ;
        RECT 282.170 0.010 293.750 2.280 ;
        RECT 294.590 0.010 306.170 2.280 ;
        RECT 307.010 0.010 318.590 2.280 ;
        RECT 319.430 0.010 331.010 2.280 ;
        RECT 331.850 0.010 343.430 2.280 ;
        RECT 344.270 0.010 355.850 2.280 ;
        RECT 356.690 0.010 368.270 2.280 ;
        RECT 369.110 0.010 380.690 2.280 ;
        RECT 381.530 0.010 393.110 2.280 ;
        RECT 393.950 0.010 401.940 2.280 ;
      LAYER met3 ;
        RECT 2.000 377.080 401.515 394.225 ;
        RECT 2.000 375.680 399.640 377.080 ;
        RECT 2.000 344.440 401.515 375.680 ;
        RECT 2.000 343.040 399.640 344.440 ;
        RECT 2.000 311.800 401.515 343.040 ;
        RECT 2.000 310.400 399.640 311.800 ;
        RECT 2.000 279.160 401.515 310.400 ;
        RECT 2.000 277.760 399.640 279.160 ;
        RECT 2.000 246.520 401.515 277.760 ;
        RECT 2.000 245.120 399.640 246.520 ;
        RECT 2.000 213.880 401.515 245.120 ;
        RECT 2.000 212.480 399.640 213.880 ;
        RECT 2.000 197.560 401.515 212.480 ;
        RECT 2.400 196.160 401.515 197.560 ;
        RECT 2.000 181.240 401.515 196.160 ;
        RECT 2.000 179.840 399.640 181.240 ;
        RECT 2.000 148.600 401.515 179.840 ;
        RECT 2.000 147.200 399.640 148.600 ;
        RECT 2.000 115.960 401.515 147.200 ;
        RECT 2.000 114.560 399.640 115.960 ;
        RECT 2.000 83.320 401.515 114.560 ;
        RECT 2.000 81.920 399.640 83.320 ;
        RECT 2.000 50.680 401.515 81.920 ;
        RECT 2.000 49.280 399.640 50.680 ;
        RECT 2.000 18.040 401.515 49.280 ;
        RECT 2.000 16.640 399.640 18.040 ;
        RECT 2.000 0.855 401.515 16.640 ;
      LAYER met4 ;
        RECT 44.455 392.320 392.545 394.225 ;
        RECT 44.455 18.535 94.680 392.320 ;
        RECT 97.080 18.535 171.480 392.320 ;
        RECT 173.880 18.535 248.280 392.320 ;
        RECT 250.680 18.535 325.080 392.320 ;
        RECT 327.480 18.535 392.545 392.320 ;
  END
END RAM128
END LIBRARY

