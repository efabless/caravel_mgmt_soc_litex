VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DFFRAM
  CLASS BLOCK ;
  FOREIGN DFFRAM ;
  ORIGIN 0.000 0.000 ;
  SIZE 550.000 BY 740.000 ;
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 27.920 550.000 28.520 ;
    END
  END A[0]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 84.360 550.000 84.960 ;
    END
  END A[1]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 141.480 550.000 142.080 ;
    END
  END A[2]
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 198.600 550.000 199.200 ;
    END
  END A[3]
  PIN A[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 255.040 550.000 255.640 ;
    END
  END A[4]
  PIN A[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 312.160 550.000 312.760 ;
    END
  END A[5]
  PIN A[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 369.280 550.000 369.880 ;
    END
  END A[6]
  PIN A[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 425.720 550.000 426.320 ;
    END
  END A[7]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END CLK
  PIN Di[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END Di[0]
  PIN Di[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END Di[10]
  PIN Di[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END Di[11]
  PIN Di[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END Di[12]
  PIN Di[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END Di[13]
  PIN Di[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END Di[14]
  PIN Di[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 0.000 258.430 4.000 ;
    END
  END Di[15]
  PIN Di[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 0.000 292.010 4.000 ;
    END
  END Di[16]
  PIN Di[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END Di[17]
  PIN Di[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.850 0.000 325.130 4.000 ;
    END
  END Di[18]
  PIN Di[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 0.000 341.690 4.000 ;
    END
  END Di[19]
  PIN Di[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END Di[1]
  PIN Di[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.430 0.000 358.710 4.000 ;
    END
  END Di[20]
  PIN Di[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END Di[21]
  PIN Di[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 0.000 391.830 4.000 ;
    END
  END Di[22]
  PIN Di[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END Di[23]
  PIN Di[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 0.000 425.410 4.000 ;
    END
  END Di[24]
  PIN Di[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.690 0.000 441.970 4.000 ;
    END
  END Di[25]
  PIN Di[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.250 0.000 458.530 4.000 ;
    END
  END Di[26]
  PIN Di[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.810 0.000 475.090 4.000 ;
    END
  END Di[27]
  PIN Di[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 0.000 492.110 4.000 ;
    END
  END Di[28]
  PIN Di[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 0.000 508.670 4.000 ;
    END
  END Di[29]
  PIN Di[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END Di[2]
  PIN Di[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END Di[30]
  PIN Di[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 0.000 541.790 4.000 ;
    END
  END Di[31]
  PIN Di[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END Di[3]
  PIN Di[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END Di[4]
  PIN Di[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 0.000 91.910 4.000 ;
    END
  END Di[5]
  PIN Di[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END Di[6]
  PIN Di[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END Di[7]
  PIN Di[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 0.000 141.590 4.000 ;
    END
  END Di[8]
  PIN Di[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END Di[9]
  PIN Do[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 736.000 8.650 740.000 ;
    END
  END Do[0]
  PIN Do[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 736.000 180.230 740.000 ;
    END
  END Do[10]
  PIN Do[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 736.000 197.710 740.000 ;
    END
  END Do[11]
  PIN Do[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 736.000 214.730 740.000 ;
    END
  END Do[12]
  PIN Do[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.470 736.000 231.750 740.000 ;
    END
  END Do[13]
  PIN Do[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 736.000 249.230 740.000 ;
    END
  END Do[14]
  PIN Do[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.970 736.000 266.250 740.000 ;
    END
  END Do[15]
  PIN Do[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 736.000 283.730 740.000 ;
    END
  END Do[16]
  PIN Do[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 736.000 300.750 740.000 ;
    END
  END Do[17]
  PIN Do[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 736.000 317.770 740.000 ;
    END
  END Do[18]
  PIN Do[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 736.000 335.250 740.000 ;
    END
  END Do[19]
  PIN Do[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.390 736.000 25.670 740.000 ;
    END
  END Do[1]
  PIN Do[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 736.000 352.270 740.000 ;
    END
  END Do[20]
  PIN Do[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 736.000 369.290 740.000 ;
    END
  END Do[21]
  PIN Do[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 736.000 386.770 740.000 ;
    END
  END Do[22]
  PIN Do[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 736.000 403.790 740.000 ;
    END
  END Do[23]
  PIN Do[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 736.000 421.270 740.000 ;
    END
  END Do[24]
  PIN Do[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 736.000 438.290 740.000 ;
    END
  END Do[25]
  PIN Do[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 736.000 455.310 740.000 ;
    END
  END Do[26]
  PIN Do[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.510 736.000 472.790 740.000 ;
    END
  END Do[27]
  PIN Do[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 736.000 489.810 740.000 ;
    END
  END Do[28]
  PIN Do[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 736.000 506.830 740.000 ;
    END
  END Do[29]
  PIN Do[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.410 736.000 42.690 740.000 ;
    END
  END Do[2]
  PIN Do[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 736.000 524.310 740.000 ;
    END
  END Do[30]
  PIN Do[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 736.000 541.330 740.000 ;
    END
  END Do[31]
  PIN Do[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 736.000 60.170 740.000 ;
    END
  END Do[3]
  PIN Do[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.910 736.000 77.190 740.000 ;
    END
  END Do[4]
  PIN Do[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.930 736.000 94.210 740.000 ;
    END
  END Do[5]
  PIN Do[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.410 736.000 111.690 740.000 ;
    END
  END Do[6]
  PIN Do[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 736.000 128.710 740.000 ;
    END
  END Do[7]
  PIN Do[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 736.000 146.190 740.000 ;
    END
  END Do[8]
  PIN Do[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 736.000 163.210 740.000 ;
    END
  END Do[9]
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 710.640 550.000 711.240 ;
    END
  END EN
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.020 0.780 549.680 2.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 91.490 549.680 93.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 221.490 549.680 223.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 351.490 549.680 353.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 481.490 549.680 483.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 611.490 549.680 613.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 737.460 549.680 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.020 0.780 1.620 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 102.440 0.780 104.040 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 256.040 0.780 257.640 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 409.640 0.780 411.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.080 0.780 549.680 739.060 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 3.320 4.080 546.380 5.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 26.490 549.680 28.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 156.490 549.680 158.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 286.490 549.680 288.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 416.490 549.680 418.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 546.490 549.680 548.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 676.490 549.680 678.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 3.320 734.160 546.380 735.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 3.320 4.080 4.920 735.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 544.780 4.080 546.380 735.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 25.640 0.780 27.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 179.240 0.780 180.840 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 332.840 0.780 334.440 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 486.440 0.780 488.040 739.060 ;
    END
  END VPWR
  PIN WE[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 482.840 550.000 483.440 ;
    END
  END WE[0]
  PIN WE[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 539.960 550.000 540.560 ;
    END
  END WE[1]
  PIN WE[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 596.400 550.000 597.000 ;
    END
  END WE[2]
  PIN WE[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 653.520 550.000 654.120 ;
    END
  END WE[3]
  OBS
      LAYER li1 ;
        RECT 9.345 10.795 539.580 729.045 ;
      LAYER met1 ;
        RECT 8.350 9.900 541.350 730.960 ;
      LAYER met2 ;
        RECT 8.930 735.720 25.110 736.170 ;
        RECT 25.950 735.720 42.130 736.170 ;
        RECT 42.970 735.720 59.610 736.170 ;
        RECT 60.450 735.720 76.630 736.170 ;
        RECT 77.470 735.720 93.650 736.170 ;
        RECT 94.490 735.720 111.130 736.170 ;
        RECT 111.970 735.720 128.150 736.170 ;
        RECT 128.990 735.720 145.630 736.170 ;
        RECT 146.470 735.720 162.650 736.170 ;
        RECT 163.490 735.720 179.670 736.170 ;
        RECT 180.510 735.720 197.150 736.170 ;
        RECT 197.990 735.720 214.170 736.170 ;
        RECT 215.010 735.720 231.190 736.170 ;
        RECT 232.030 735.720 248.670 736.170 ;
        RECT 249.510 735.720 265.690 736.170 ;
        RECT 266.530 735.720 283.170 736.170 ;
        RECT 284.010 735.720 300.190 736.170 ;
        RECT 301.030 735.720 317.210 736.170 ;
        RECT 318.050 735.720 334.690 736.170 ;
        RECT 335.530 735.720 351.710 736.170 ;
        RECT 352.550 735.720 368.730 736.170 ;
        RECT 369.570 735.720 386.210 736.170 ;
        RECT 387.050 735.720 403.230 736.170 ;
        RECT 404.070 735.720 420.710 736.170 ;
        RECT 421.550 735.720 437.730 736.170 ;
        RECT 438.570 735.720 454.750 736.170 ;
        RECT 455.590 735.720 472.230 736.170 ;
        RECT 473.070 735.720 489.250 736.170 ;
        RECT 490.090 735.720 506.270 736.170 ;
        RECT 507.110 735.720 523.750 736.170 ;
        RECT 524.590 735.720 540.770 736.170 ;
        RECT 541.610 735.720 541.720 736.170 ;
        RECT 8.370 4.280 541.720 735.720 ;
        RECT 8.930 3.670 24.650 4.280 ;
        RECT 25.490 3.670 41.210 4.280 ;
        RECT 42.050 3.670 57.770 4.280 ;
        RECT 58.610 3.670 74.330 4.280 ;
        RECT 75.170 3.670 91.350 4.280 ;
        RECT 92.190 3.670 107.910 4.280 ;
        RECT 108.750 3.670 124.470 4.280 ;
        RECT 125.310 3.670 141.030 4.280 ;
        RECT 141.870 3.670 158.050 4.280 ;
        RECT 158.890 3.670 174.610 4.280 ;
        RECT 175.450 3.670 191.170 4.280 ;
        RECT 192.010 3.670 207.730 4.280 ;
        RECT 208.570 3.670 224.750 4.280 ;
        RECT 225.590 3.670 241.310 4.280 ;
        RECT 242.150 3.670 257.870 4.280 ;
        RECT 258.710 3.670 274.430 4.280 ;
        RECT 275.270 3.670 291.450 4.280 ;
        RECT 292.290 3.670 308.010 4.280 ;
        RECT 308.850 3.670 324.570 4.280 ;
        RECT 325.410 3.670 341.130 4.280 ;
        RECT 341.970 3.670 358.150 4.280 ;
        RECT 358.990 3.670 374.710 4.280 ;
        RECT 375.550 3.670 391.270 4.280 ;
        RECT 392.110 3.670 407.830 4.280 ;
        RECT 408.670 3.670 424.850 4.280 ;
        RECT 425.690 3.670 441.410 4.280 ;
        RECT 442.250 3.670 457.970 4.280 ;
        RECT 458.810 3.670 474.530 4.280 ;
        RECT 475.370 3.670 491.550 4.280 ;
        RECT 492.390 3.670 508.110 4.280 ;
        RECT 508.950 3.670 524.670 4.280 ;
        RECT 525.510 3.670 541.230 4.280 ;
      LAYER met3 ;
        RECT 8.345 711.640 546.000 729.125 ;
        RECT 8.345 710.240 545.600 711.640 ;
        RECT 8.345 654.520 546.000 710.240 ;
        RECT 8.345 653.120 545.600 654.520 ;
        RECT 8.345 597.400 546.000 653.120 ;
        RECT 8.345 596.000 545.600 597.400 ;
        RECT 8.345 540.960 546.000 596.000 ;
        RECT 8.345 539.560 545.600 540.960 ;
        RECT 8.345 483.840 546.000 539.560 ;
        RECT 8.345 482.440 545.600 483.840 ;
        RECT 8.345 426.720 546.000 482.440 ;
        RECT 8.345 425.320 545.600 426.720 ;
        RECT 8.345 370.280 546.000 425.320 ;
        RECT 8.345 368.880 545.600 370.280 ;
        RECT 8.345 313.160 546.000 368.880 ;
        RECT 8.345 311.760 545.600 313.160 ;
        RECT 8.345 256.040 546.000 311.760 ;
        RECT 8.345 254.640 545.600 256.040 ;
        RECT 8.345 199.600 546.000 254.640 ;
        RECT 8.345 198.200 545.600 199.600 ;
        RECT 8.345 142.480 546.000 198.200 ;
        RECT 8.345 141.080 545.600 142.480 ;
        RECT 8.345 85.360 546.000 141.080 ;
        RECT 8.345 83.960 545.600 85.360 ;
        RECT 8.345 28.920 546.000 83.960 ;
        RECT 8.345 27.520 545.600 28.920 ;
        RECT 8.345 10.715 546.000 27.520 ;
      LAYER met4 ;
        RECT 22.375 14.455 25.240 727.425 ;
        RECT 27.640 14.455 102.040 727.425 ;
        RECT 104.440 14.455 178.840 727.425 ;
        RECT 181.240 14.455 255.640 727.425 ;
        RECT 258.040 14.455 332.440 727.425 ;
        RECT 334.840 14.455 409.240 727.425 ;
        RECT 411.640 14.455 486.040 727.425 ;
        RECT 488.440 14.455 500.185 727.425 ;
  END
END DFFRAM
END LIBRARY

