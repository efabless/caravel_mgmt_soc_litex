magic
tech sky130A
magscale 1 2
timestamp 1638166645
<< obsli1 >>
rect 2024 2159 397900 145809
<< obsm1 >>
rect 290 1300 399634 146532
<< metal2 >>
rect 294 147200 350 148000
rect 938 147200 994 148000
rect 1582 147200 1638 148000
rect 2226 147200 2282 148000
rect 2870 147200 2926 148000
rect 3514 147200 3570 148000
rect 4158 147200 4214 148000
rect 4802 147200 4858 148000
rect 5446 147200 5502 148000
rect 6090 147200 6146 148000
rect 6734 147200 6790 148000
rect 7378 147200 7434 148000
rect 8022 147200 8078 148000
rect 8666 147200 8722 148000
rect 9310 147200 9366 148000
rect 10046 147200 10102 148000
rect 10690 147200 10746 148000
rect 11334 147200 11390 148000
rect 11978 147200 12034 148000
rect 12622 147200 12678 148000
rect 13266 147200 13322 148000
rect 13910 147200 13966 148000
rect 14554 147200 14610 148000
rect 15198 147200 15254 148000
rect 15842 147200 15898 148000
rect 16486 147200 16542 148000
rect 17130 147200 17186 148000
rect 17774 147200 17830 148000
rect 18418 147200 18474 148000
rect 19154 147200 19210 148000
rect 19798 147200 19854 148000
rect 20442 147200 20498 148000
rect 21086 147200 21142 148000
rect 21730 147200 21786 148000
rect 22374 147200 22430 148000
rect 23018 147200 23074 148000
rect 23662 147200 23718 148000
rect 24306 147200 24362 148000
rect 24950 147200 25006 148000
rect 25594 147200 25650 148000
rect 26238 147200 26294 148000
rect 26882 147200 26938 148000
rect 27526 147200 27582 148000
rect 28262 147200 28318 148000
rect 28906 147200 28962 148000
rect 29550 147200 29606 148000
rect 30194 147200 30250 148000
rect 30838 147200 30894 148000
rect 31482 147200 31538 148000
rect 32126 147200 32182 148000
rect 32770 147200 32826 148000
rect 33414 147200 33470 148000
rect 34058 147200 34114 148000
rect 34702 147200 34758 148000
rect 35346 147200 35402 148000
rect 35990 147200 36046 148000
rect 36634 147200 36690 148000
rect 37278 147200 37334 148000
rect 38014 147200 38070 148000
rect 38658 147200 38714 148000
rect 39302 147200 39358 148000
rect 39946 147200 40002 148000
rect 40590 147200 40646 148000
rect 41234 147200 41290 148000
rect 41878 147200 41934 148000
rect 42522 147200 42578 148000
rect 43166 147200 43222 148000
rect 43810 147200 43866 148000
rect 44454 147200 44510 148000
rect 45098 147200 45154 148000
rect 45742 147200 45798 148000
rect 46386 147200 46442 148000
rect 47122 147200 47178 148000
rect 47766 147200 47822 148000
rect 48410 147200 48466 148000
rect 49054 147200 49110 148000
rect 49698 147200 49754 148000
rect 50342 147200 50398 148000
rect 50986 147200 51042 148000
rect 51630 147200 51686 148000
rect 52274 147200 52330 148000
rect 52918 147200 52974 148000
rect 53562 147200 53618 148000
rect 54206 147200 54262 148000
rect 54850 147200 54906 148000
rect 55494 147200 55550 148000
rect 56230 147200 56286 148000
rect 56874 147200 56930 148000
rect 57518 147200 57574 148000
rect 58162 147200 58218 148000
rect 58806 147200 58862 148000
rect 59450 147200 59506 148000
rect 60094 147200 60150 148000
rect 60738 147200 60794 148000
rect 61382 147200 61438 148000
rect 62026 147200 62082 148000
rect 62670 147200 62726 148000
rect 63314 147200 63370 148000
rect 63958 147200 64014 148000
rect 64602 147200 64658 148000
rect 65246 147200 65302 148000
rect 65982 147200 66038 148000
rect 66626 147200 66682 148000
rect 67270 147200 67326 148000
rect 67914 147200 67970 148000
rect 68558 147200 68614 148000
rect 69202 147200 69258 148000
rect 69846 147200 69902 148000
rect 70490 147200 70546 148000
rect 71134 147200 71190 148000
rect 71778 147200 71834 148000
rect 72422 147200 72478 148000
rect 73066 147200 73122 148000
rect 73710 147200 73766 148000
rect 74354 147200 74410 148000
rect 75090 147200 75146 148000
rect 75734 147200 75790 148000
rect 76378 147200 76434 148000
rect 77022 147200 77078 148000
rect 77666 147200 77722 148000
rect 78310 147200 78366 148000
rect 78954 147200 79010 148000
rect 79598 147200 79654 148000
rect 80242 147200 80298 148000
rect 80886 147200 80942 148000
rect 81530 147200 81586 148000
rect 82174 147200 82230 148000
rect 82818 147200 82874 148000
rect 83462 147200 83518 148000
rect 84198 147200 84254 148000
rect 84842 147200 84898 148000
rect 85486 147200 85542 148000
rect 86130 147200 86186 148000
rect 86774 147200 86830 148000
rect 87418 147200 87474 148000
rect 88062 147200 88118 148000
rect 88706 147200 88762 148000
rect 89350 147200 89406 148000
rect 89994 147200 90050 148000
rect 90638 147200 90694 148000
rect 91282 147200 91338 148000
rect 91926 147200 91982 148000
rect 92570 147200 92626 148000
rect 93214 147200 93270 148000
rect 93950 147200 94006 148000
rect 94594 147200 94650 148000
rect 95238 147200 95294 148000
rect 95882 147200 95938 148000
rect 96526 147200 96582 148000
rect 97170 147200 97226 148000
rect 97814 147200 97870 148000
rect 98458 147200 98514 148000
rect 99102 147200 99158 148000
rect 99746 147200 99802 148000
rect 100390 147200 100446 148000
rect 101034 147200 101090 148000
rect 101678 147200 101734 148000
rect 102322 147200 102378 148000
rect 103058 147200 103114 148000
rect 103702 147200 103758 148000
rect 104346 147200 104402 148000
rect 104990 147200 105046 148000
rect 105634 147200 105690 148000
rect 106278 147200 106334 148000
rect 106922 147200 106978 148000
rect 107566 147200 107622 148000
rect 108210 147200 108266 148000
rect 108854 147200 108910 148000
rect 109498 147200 109554 148000
rect 110142 147200 110198 148000
rect 110786 147200 110842 148000
rect 111430 147200 111486 148000
rect 112166 147200 112222 148000
rect 112810 147200 112866 148000
rect 113454 147200 113510 148000
rect 114098 147200 114154 148000
rect 114742 147200 114798 148000
rect 115386 147200 115442 148000
rect 116030 147200 116086 148000
rect 116674 147200 116730 148000
rect 117318 147200 117374 148000
rect 117962 147200 118018 148000
rect 118606 147200 118662 148000
rect 119250 147200 119306 148000
rect 119894 147200 119950 148000
rect 120538 147200 120594 148000
rect 121274 147200 121330 148000
rect 121918 147200 121974 148000
rect 122562 147200 122618 148000
rect 123206 147200 123262 148000
rect 123850 147200 123906 148000
rect 124494 147200 124550 148000
rect 125138 147200 125194 148000
rect 125782 147200 125838 148000
rect 126426 147200 126482 148000
rect 127070 147200 127126 148000
rect 127714 147200 127770 148000
rect 128358 147200 128414 148000
rect 129002 147200 129058 148000
rect 129646 147200 129702 148000
rect 130290 147200 130346 148000
rect 131026 147200 131082 148000
rect 131670 147200 131726 148000
rect 132314 147200 132370 148000
rect 132958 147200 133014 148000
rect 133602 147200 133658 148000
rect 134246 147200 134302 148000
rect 134890 147200 134946 148000
rect 135534 147200 135590 148000
rect 136178 147200 136234 148000
rect 136822 147200 136878 148000
rect 137466 147200 137522 148000
rect 138110 147200 138166 148000
rect 138754 147200 138810 148000
rect 139398 147200 139454 148000
rect 140134 147200 140190 148000
rect 140778 147200 140834 148000
rect 141422 147200 141478 148000
rect 142066 147200 142122 148000
rect 142710 147200 142766 148000
rect 143354 147200 143410 148000
rect 143998 147200 144054 148000
rect 144642 147200 144698 148000
rect 145286 147200 145342 148000
rect 145930 147200 145986 148000
rect 146574 147200 146630 148000
rect 147218 147200 147274 148000
rect 147862 147200 147918 148000
rect 148506 147200 148562 148000
rect 149242 147200 149298 148000
rect 149886 147200 149942 148000
rect 150530 147200 150586 148000
rect 151174 147200 151230 148000
rect 151818 147200 151874 148000
rect 152462 147200 152518 148000
rect 153106 147200 153162 148000
rect 153750 147200 153806 148000
rect 154394 147200 154450 148000
rect 155038 147200 155094 148000
rect 155682 147200 155738 148000
rect 156326 147200 156382 148000
rect 156970 147200 157026 148000
rect 157614 147200 157670 148000
rect 158258 147200 158314 148000
rect 158994 147200 159050 148000
rect 159638 147200 159694 148000
rect 160282 147200 160338 148000
rect 160926 147200 160982 148000
rect 161570 147200 161626 148000
rect 162214 147200 162270 148000
rect 162858 147200 162914 148000
rect 163502 147200 163558 148000
rect 164146 147200 164202 148000
rect 164790 147200 164846 148000
rect 165434 147200 165490 148000
rect 166078 147200 166134 148000
rect 166722 147200 166778 148000
rect 167366 147200 167422 148000
rect 168102 147200 168158 148000
rect 168746 147200 168802 148000
rect 169390 147200 169446 148000
rect 170034 147200 170090 148000
rect 170678 147200 170734 148000
rect 171322 147200 171378 148000
rect 171966 147200 172022 148000
rect 172610 147200 172666 148000
rect 173254 147200 173310 148000
rect 173898 147200 173954 148000
rect 174542 147200 174598 148000
rect 175186 147200 175242 148000
rect 175830 147200 175886 148000
rect 176474 147200 176530 148000
rect 177210 147200 177266 148000
rect 177854 147200 177910 148000
rect 178498 147200 178554 148000
rect 179142 147200 179198 148000
rect 179786 147200 179842 148000
rect 180430 147200 180486 148000
rect 181074 147200 181130 148000
rect 181718 147200 181774 148000
rect 182362 147200 182418 148000
rect 183006 147200 183062 148000
rect 183650 147200 183706 148000
rect 184294 147200 184350 148000
rect 184938 147200 184994 148000
rect 185582 147200 185638 148000
rect 186226 147200 186282 148000
rect 186962 147200 187018 148000
rect 187606 147200 187662 148000
rect 188250 147200 188306 148000
rect 188894 147200 188950 148000
rect 189538 147200 189594 148000
rect 190182 147200 190238 148000
rect 190826 147200 190882 148000
rect 191470 147200 191526 148000
rect 192114 147200 192170 148000
rect 192758 147200 192814 148000
rect 193402 147200 193458 148000
rect 194046 147200 194102 148000
rect 194690 147200 194746 148000
rect 195334 147200 195390 148000
rect 196070 147200 196126 148000
rect 196714 147200 196770 148000
rect 197358 147200 197414 148000
rect 198002 147200 198058 148000
rect 198646 147200 198702 148000
rect 199290 147200 199346 148000
rect 199934 147200 199990 148000
rect 200578 147200 200634 148000
rect 201222 147200 201278 148000
rect 201866 147200 201922 148000
rect 202510 147200 202566 148000
rect 203154 147200 203210 148000
rect 203798 147200 203854 148000
rect 204442 147200 204498 148000
rect 205178 147200 205234 148000
rect 205822 147200 205878 148000
rect 206466 147200 206522 148000
rect 207110 147200 207166 148000
rect 207754 147200 207810 148000
rect 208398 147200 208454 148000
rect 209042 147200 209098 148000
rect 209686 147200 209742 148000
rect 210330 147200 210386 148000
rect 210974 147200 211030 148000
rect 211618 147200 211674 148000
rect 212262 147200 212318 148000
rect 212906 147200 212962 148000
rect 213550 147200 213606 148000
rect 214286 147200 214342 148000
rect 214930 147200 214986 148000
rect 215574 147200 215630 148000
rect 216218 147200 216274 148000
rect 216862 147200 216918 148000
rect 217506 147200 217562 148000
rect 218150 147200 218206 148000
rect 218794 147200 218850 148000
rect 219438 147200 219494 148000
rect 220082 147200 220138 148000
rect 220726 147200 220782 148000
rect 221370 147200 221426 148000
rect 222014 147200 222070 148000
rect 222658 147200 222714 148000
rect 223302 147200 223358 148000
rect 224038 147200 224094 148000
rect 224682 147200 224738 148000
rect 225326 147200 225382 148000
rect 225970 147200 226026 148000
rect 226614 147200 226670 148000
rect 227258 147200 227314 148000
rect 227902 147200 227958 148000
rect 228546 147200 228602 148000
rect 229190 147200 229246 148000
rect 229834 147200 229890 148000
rect 230478 147200 230534 148000
rect 231122 147200 231178 148000
rect 231766 147200 231822 148000
rect 232410 147200 232466 148000
rect 233146 147200 233202 148000
rect 233790 147200 233846 148000
rect 234434 147200 234490 148000
rect 235078 147200 235134 148000
rect 235722 147200 235778 148000
rect 236366 147200 236422 148000
rect 237010 147200 237066 148000
rect 237654 147200 237710 148000
rect 238298 147200 238354 148000
rect 238942 147200 238998 148000
rect 239586 147200 239642 148000
rect 240230 147200 240286 148000
rect 240874 147200 240930 148000
rect 241518 147200 241574 148000
rect 242254 147200 242310 148000
rect 242898 147200 242954 148000
rect 243542 147200 243598 148000
rect 244186 147200 244242 148000
rect 244830 147200 244886 148000
rect 245474 147200 245530 148000
rect 246118 147200 246174 148000
rect 246762 147200 246818 148000
rect 247406 147200 247462 148000
rect 248050 147200 248106 148000
rect 248694 147200 248750 148000
rect 249338 147200 249394 148000
rect 249982 147200 250038 148000
rect 250626 147200 250682 148000
rect 251270 147200 251326 148000
rect 252006 147200 252062 148000
rect 252650 147200 252706 148000
rect 253294 147200 253350 148000
rect 253938 147200 253994 148000
rect 254582 147200 254638 148000
rect 255226 147200 255282 148000
rect 255870 147200 255926 148000
rect 256514 147200 256570 148000
rect 257158 147200 257214 148000
rect 257802 147200 257858 148000
rect 258446 147200 258502 148000
rect 259090 147200 259146 148000
rect 259734 147200 259790 148000
rect 260378 147200 260434 148000
rect 261114 147200 261170 148000
rect 261758 147200 261814 148000
rect 262402 147200 262458 148000
rect 263046 147200 263102 148000
rect 263690 147200 263746 148000
rect 264334 147200 264390 148000
rect 264978 147200 265034 148000
rect 265622 147200 265678 148000
rect 266266 147200 266322 148000
rect 266910 147200 266966 148000
rect 267554 147200 267610 148000
rect 268198 147200 268254 148000
rect 268842 147200 268898 148000
rect 269486 147200 269542 148000
rect 270222 147200 270278 148000
rect 270866 147200 270922 148000
rect 271510 147200 271566 148000
rect 272154 147200 272210 148000
rect 272798 147200 272854 148000
rect 273442 147200 273498 148000
rect 274086 147200 274142 148000
rect 274730 147200 274786 148000
rect 275374 147200 275430 148000
rect 276018 147200 276074 148000
rect 276662 147200 276718 148000
rect 277306 147200 277362 148000
rect 277950 147200 278006 148000
rect 278594 147200 278650 148000
rect 279238 147200 279294 148000
rect 279974 147200 280030 148000
rect 280618 147200 280674 148000
rect 281262 147200 281318 148000
rect 281906 147200 281962 148000
rect 282550 147200 282606 148000
rect 283194 147200 283250 148000
rect 283838 147200 283894 148000
rect 284482 147200 284538 148000
rect 285126 147200 285182 148000
rect 285770 147200 285826 148000
rect 286414 147200 286470 148000
rect 287058 147200 287114 148000
rect 287702 147200 287758 148000
rect 288346 147200 288402 148000
rect 289082 147200 289138 148000
rect 289726 147200 289782 148000
rect 290370 147200 290426 148000
rect 291014 147200 291070 148000
rect 291658 147200 291714 148000
rect 292302 147200 292358 148000
rect 292946 147200 293002 148000
rect 293590 147200 293646 148000
rect 294234 147200 294290 148000
rect 294878 147200 294934 148000
rect 295522 147200 295578 148000
rect 296166 147200 296222 148000
rect 296810 147200 296866 148000
rect 297454 147200 297510 148000
rect 298190 147200 298246 148000
rect 298834 147200 298890 148000
rect 299478 147200 299534 148000
rect 300122 147200 300178 148000
rect 300766 147200 300822 148000
rect 301410 147200 301466 148000
rect 302054 147200 302110 148000
rect 302698 147200 302754 148000
rect 303342 147200 303398 148000
rect 303986 147200 304042 148000
rect 304630 147200 304686 148000
rect 305274 147200 305330 148000
rect 305918 147200 305974 148000
rect 306562 147200 306618 148000
rect 307298 147200 307354 148000
rect 307942 147200 307998 148000
rect 308586 147200 308642 148000
rect 309230 147200 309286 148000
rect 309874 147200 309930 148000
rect 310518 147200 310574 148000
rect 311162 147200 311218 148000
rect 311806 147200 311862 148000
rect 312450 147200 312506 148000
rect 313094 147200 313150 148000
rect 313738 147200 313794 148000
rect 314382 147200 314438 148000
rect 315026 147200 315082 148000
rect 315670 147200 315726 148000
rect 316314 147200 316370 148000
rect 317050 147200 317106 148000
rect 317694 147200 317750 148000
rect 318338 147200 318394 148000
rect 318982 147200 319038 148000
rect 319626 147200 319682 148000
rect 320270 147200 320326 148000
rect 320914 147200 320970 148000
rect 321558 147200 321614 148000
rect 322202 147200 322258 148000
rect 322846 147200 322902 148000
rect 323490 147200 323546 148000
rect 324134 147200 324190 148000
rect 324778 147200 324834 148000
rect 325422 147200 325478 148000
rect 326158 147200 326214 148000
rect 326802 147200 326858 148000
rect 327446 147200 327502 148000
rect 328090 147200 328146 148000
rect 328734 147200 328790 148000
rect 329378 147200 329434 148000
rect 330022 147200 330078 148000
rect 330666 147200 330722 148000
rect 331310 147200 331366 148000
rect 331954 147200 332010 148000
rect 332598 147200 332654 148000
rect 333242 147200 333298 148000
rect 333886 147200 333942 148000
rect 334530 147200 334586 148000
rect 335266 147200 335322 148000
rect 335910 147200 335966 148000
rect 336554 147200 336610 148000
rect 337198 147200 337254 148000
rect 337842 147200 337898 148000
rect 338486 147200 338542 148000
rect 339130 147200 339186 148000
rect 339774 147200 339830 148000
rect 340418 147200 340474 148000
rect 341062 147200 341118 148000
rect 341706 147200 341762 148000
rect 342350 147200 342406 148000
rect 342994 147200 343050 148000
rect 343638 147200 343694 148000
rect 344282 147200 344338 148000
rect 345018 147200 345074 148000
rect 345662 147200 345718 148000
rect 346306 147200 346362 148000
rect 346950 147200 347006 148000
rect 347594 147200 347650 148000
rect 348238 147200 348294 148000
rect 348882 147200 348938 148000
rect 349526 147200 349582 148000
rect 350170 147200 350226 148000
rect 350814 147200 350870 148000
rect 351458 147200 351514 148000
rect 352102 147200 352158 148000
rect 352746 147200 352802 148000
rect 353390 147200 353446 148000
rect 354126 147200 354182 148000
rect 354770 147200 354826 148000
rect 355414 147200 355470 148000
rect 356058 147200 356114 148000
rect 356702 147200 356758 148000
rect 357346 147200 357402 148000
rect 357990 147200 358046 148000
rect 358634 147200 358690 148000
rect 359278 147200 359334 148000
rect 359922 147200 359978 148000
rect 360566 147200 360622 148000
rect 361210 147200 361266 148000
rect 361854 147200 361910 148000
rect 362498 147200 362554 148000
rect 363234 147200 363290 148000
rect 363878 147200 363934 148000
rect 364522 147200 364578 148000
rect 365166 147200 365222 148000
rect 365810 147200 365866 148000
rect 366454 147200 366510 148000
rect 367098 147200 367154 148000
rect 367742 147200 367798 148000
rect 368386 147200 368442 148000
rect 369030 147200 369086 148000
rect 369674 147200 369730 148000
rect 370318 147200 370374 148000
rect 370962 147200 371018 148000
rect 371606 147200 371662 148000
rect 372250 147200 372306 148000
rect 372986 147200 373042 148000
rect 373630 147200 373686 148000
rect 374274 147200 374330 148000
rect 374918 147200 374974 148000
rect 375562 147200 375618 148000
rect 376206 147200 376262 148000
rect 376850 147200 376906 148000
rect 377494 147200 377550 148000
rect 378138 147200 378194 148000
rect 378782 147200 378838 148000
rect 379426 147200 379482 148000
rect 380070 147200 380126 148000
rect 380714 147200 380770 148000
rect 381358 147200 381414 148000
rect 382094 147200 382150 148000
rect 382738 147200 382794 148000
rect 383382 147200 383438 148000
rect 384026 147200 384082 148000
rect 384670 147200 384726 148000
rect 385314 147200 385370 148000
rect 385958 147200 386014 148000
rect 386602 147200 386658 148000
rect 387246 147200 387302 148000
rect 387890 147200 387946 148000
rect 388534 147200 388590 148000
rect 389178 147200 389234 148000
rect 389822 147200 389878 148000
rect 390466 147200 390522 148000
rect 391202 147200 391258 148000
rect 391846 147200 391902 148000
rect 392490 147200 392546 148000
rect 393134 147200 393190 148000
rect 393778 147200 393834 148000
rect 394422 147200 394478 148000
rect 395066 147200 395122 148000
rect 395710 147200 395766 148000
rect 396354 147200 396410 148000
rect 396998 147200 397054 148000
rect 397642 147200 397698 148000
rect 398286 147200 398342 148000
rect 398930 147200 398986 148000
rect 399574 147200 399630 148000
rect 1674 0 1730 800
rect 4986 0 5042 800
rect 8390 0 8446 800
rect 11702 0 11758 800
rect 15106 0 15162 800
rect 18418 0 18474 800
rect 21822 0 21878 800
rect 25134 0 25190 800
rect 28538 0 28594 800
rect 31850 0 31906 800
rect 35254 0 35310 800
rect 38566 0 38622 800
rect 41970 0 42026 800
rect 45282 0 45338 800
rect 48686 0 48742 800
rect 52090 0 52146 800
rect 55402 0 55458 800
rect 58806 0 58862 800
rect 62118 0 62174 800
rect 65522 0 65578 800
rect 68834 0 68890 800
rect 72238 0 72294 800
rect 75550 0 75606 800
rect 78954 0 79010 800
rect 82266 0 82322 800
rect 85670 0 85726 800
rect 88982 0 89038 800
rect 92386 0 92442 800
rect 95790 0 95846 800
rect 99102 0 99158 800
rect 102506 0 102562 800
rect 105818 0 105874 800
rect 109222 0 109278 800
rect 112534 0 112590 800
rect 115938 0 115994 800
rect 119250 0 119306 800
rect 122654 0 122710 800
rect 125966 0 126022 800
rect 129370 0 129426 800
rect 132682 0 132738 800
rect 136086 0 136142 800
rect 139490 0 139546 800
rect 142802 0 142858 800
rect 146206 0 146262 800
rect 149518 0 149574 800
rect 152922 0 152978 800
rect 156234 0 156290 800
rect 159638 0 159694 800
rect 162950 0 163006 800
rect 166354 0 166410 800
rect 169666 0 169722 800
rect 173070 0 173126 800
rect 176382 0 176438 800
rect 179786 0 179842 800
rect 183190 0 183246 800
rect 186502 0 186558 800
rect 189906 0 189962 800
rect 193218 0 193274 800
rect 196622 0 196678 800
rect 199934 0 199990 800
rect 203338 0 203394 800
rect 206650 0 206706 800
rect 210054 0 210110 800
rect 213366 0 213422 800
rect 216770 0 216826 800
rect 220082 0 220138 800
rect 223486 0 223542 800
rect 226890 0 226946 800
rect 230202 0 230258 800
rect 233606 0 233662 800
rect 236918 0 236974 800
rect 240322 0 240378 800
rect 243634 0 243690 800
rect 247038 0 247094 800
rect 250350 0 250406 800
rect 253754 0 253810 800
rect 257066 0 257122 800
rect 260470 0 260526 800
rect 263782 0 263838 800
rect 267186 0 267242 800
rect 270590 0 270646 800
rect 273902 0 273958 800
rect 277306 0 277362 800
rect 280618 0 280674 800
rect 284022 0 284078 800
rect 287334 0 287390 800
rect 290738 0 290794 800
rect 294050 0 294106 800
rect 297454 0 297510 800
rect 300766 0 300822 800
rect 304170 0 304226 800
rect 307482 0 307538 800
rect 310886 0 310942 800
rect 314290 0 314346 800
rect 317602 0 317658 800
rect 321006 0 321062 800
rect 324318 0 324374 800
rect 327722 0 327778 800
rect 331034 0 331090 800
rect 334438 0 334494 800
rect 337750 0 337806 800
rect 341154 0 341210 800
rect 344466 0 344522 800
rect 347870 0 347926 800
rect 351182 0 351238 800
rect 354586 0 354642 800
rect 357990 0 358046 800
rect 361302 0 361358 800
rect 364706 0 364762 800
rect 368018 0 368074 800
rect 371422 0 371478 800
rect 374734 0 374790 800
rect 378138 0 378194 800
rect 381450 0 381506 800
rect 384854 0 384910 800
rect 388166 0 388222 800
rect 391570 0 391626 800
rect 394882 0 394938 800
rect 398286 0 398342 800
<< obsm2 >>
rect 406 147144 882 147234
rect 1050 147144 1526 147234
rect 1694 147144 2170 147234
rect 2338 147144 2814 147234
rect 2982 147144 3458 147234
rect 3626 147144 4102 147234
rect 4270 147144 4746 147234
rect 4914 147144 5390 147234
rect 5558 147144 6034 147234
rect 6202 147144 6678 147234
rect 6846 147144 7322 147234
rect 7490 147144 7966 147234
rect 8134 147144 8610 147234
rect 8778 147144 9254 147234
rect 9422 147144 9990 147234
rect 10158 147144 10634 147234
rect 10802 147144 11278 147234
rect 11446 147144 11922 147234
rect 12090 147144 12566 147234
rect 12734 147144 13210 147234
rect 13378 147144 13854 147234
rect 14022 147144 14498 147234
rect 14666 147144 15142 147234
rect 15310 147144 15786 147234
rect 15954 147144 16430 147234
rect 16598 147144 17074 147234
rect 17242 147144 17718 147234
rect 17886 147144 18362 147234
rect 18530 147144 19098 147234
rect 19266 147144 19742 147234
rect 19910 147144 20386 147234
rect 20554 147144 21030 147234
rect 21198 147144 21674 147234
rect 21842 147144 22318 147234
rect 22486 147144 22962 147234
rect 23130 147144 23606 147234
rect 23774 147144 24250 147234
rect 24418 147144 24894 147234
rect 25062 147144 25538 147234
rect 25706 147144 26182 147234
rect 26350 147144 26826 147234
rect 26994 147144 27470 147234
rect 27638 147144 28206 147234
rect 28374 147144 28850 147234
rect 29018 147144 29494 147234
rect 29662 147144 30138 147234
rect 30306 147144 30782 147234
rect 30950 147144 31426 147234
rect 31594 147144 32070 147234
rect 32238 147144 32714 147234
rect 32882 147144 33358 147234
rect 33526 147144 34002 147234
rect 34170 147144 34646 147234
rect 34814 147144 35290 147234
rect 35458 147144 35934 147234
rect 36102 147144 36578 147234
rect 36746 147144 37222 147234
rect 37390 147144 37958 147234
rect 38126 147144 38602 147234
rect 38770 147144 39246 147234
rect 39414 147144 39890 147234
rect 40058 147144 40534 147234
rect 40702 147144 41178 147234
rect 41346 147144 41822 147234
rect 41990 147144 42466 147234
rect 42634 147144 43110 147234
rect 43278 147144 43754 147234
rect 43922 147144 44398 147234
rect 44566 147144 45042 147234
rect 45210 147144 45686 147234
rect 45854 147144 46330 147234
rect 46498 147144 47066 147234
rect 47234 147144 47710 147234
rect 47878 147144 48354 147234
rect 48522 147144 48998 147234
rect 49166 147144 49642 147234
rect 49810 147144 50286 147234
rect 50454 147144 50930 147234
rect 51098 147144 51574 147234
rect 51742 147144 52218 147234
rect 52386 147144 52862 147234
rect 53030 147144 53506 147234
rect 53674 147144 54150 147234
rect 54318 147144 54794 147234
rect 54962 147144 55438 147234
rect 55606 147144 56174 147234
rect 56342 147144 56818 147234
rect 56986 147144 57462 147234
rect 57630 147144 58106 147234
rect 58274 147144 58750 147234
rect 58918 147144 59394 147234
rect 59562 147144 60038 147234
rect 60206 147144 60682 147234
rect 60850 147144 61326 147234
rect 61494 147144 61970 147234
rect 62138 147144 62614 147234
rect 62782 147144 63258 147234
rect 63426 147144 63902 147234
rect 64070 147144 64546 147234
rect 64714 147144 65190 147234
rect 65358 147144 65926 147234
rect 66094 147144 66570 147234
rect 66738 147144 67214 147234
rect 67382 147144 67858 147234
rect 68026 147144 68502 147234
rect 68670 147144 69146 147234
rect 69314 147144 69790 147234
rect 69958 147144 70434 147234
rect 70602 147144 71078 147234
rect 71246 147144 71722 147234
rect 71890 147144 72366 147234
rect 72534 147144 73010 147234
rect 73178 147144 73654 147234
rect 73822 147144 74298 147234
rect 74466 147144 75034 147234
rect 75202 147144 75678 147234
rect 75846 147144 76322 147234
rect 76490 147144 76966 147234
rect 77134 147144 77610 147234
rect 77778 147144 78254 147234
rect 78422 147144 78898 147234
rect 79066 147144 79542 147234
rect 79710 147144 80186 147234
rect 80354 147144 80830 147234
rect 80998 147144 81474 147234
rect 81642 147144 82118 147234
rect 82286 147144 82762 147234
rect 82930 147144 83406 147234
rect 83574 147144 84142 147234
rect 84310 147144 84786 147234
rect 84954 147144 85430 147234
rect 85598 147144 86074 147234
rect 86242 147144 86718 147234
rect 86886 147144 87362 147234
rect 87530 147144 88006 147234
rect 88174 147144 88650 147234
rect 88818 147144 89294 147234
rect 89462 147144 89938 147234
rect 90106 147144 90582 147234
rect 90750 147144 91226 147234
rect 91394 147144 91870 147234
rect 92038 147144 92514 147234
rect 92682 147144 93158 147234
rect 93326 147144 93894 147234
rect 94062 147144 94538 147234
rect 94706 147144 95182 147234
rect 95350 147144 95826 147234
rect 95994 147144 96470 147234
rect 96638 147144 97114 147234
rect 97282 147144 97758 147234
rect 97926 147144 98402 147234
rect 98570 147144 99046 147234
rect 99214 147144 99690 147234
rect 99858 147144 100334 147234
rect 100502 147144 100978 147234
rect 101146 147144 101622 147234
rect 101790 147144 102266 147234
rect 102434 147144 103002 147234
rect 103170 147144 103646 147234
rect 103814 147144 104290 147234
rect 104458 147144 104934 147234
rect 105102 147144 105578 147234
rect 105746 147144 106222 147234
rect 106390 147144 106866 147234
rect 107034 147144 107510 147234
rect 107678 147144 108154 147234
rect 108322 147144 108798 147234
rect 108966 147144 109442 147234
rect 109610 147144 110086 147234
rect 110254 147144 110730 147234
rect 110898 147144 111374 147234
rect 111542 147144 112110 147234
rect 112278 147144 112754 147234
rect 112922 147144 113398 147234
rect 113566 147144 114042 147234
rect 114210 147144 114686 147234
rect 114854 147144 115330 147234
rect 115498 147144 115974 147234
rect 116142 147144 116618 147234
rect 116786 147144 117262 147234
rect 117430 147144 117906 147234
rect 118074 147144 118550 147234
rect 118718 147144 119194 147234
rect 119362 147144 119838 147234
rect 120006 147144 120482 147234
rect 120650 147144 121218 147234
rect 121386 147144 121862 147234
rect 122030 147144 122506 147234
rect 122674 147144 123150 147234
rect 123318 147144 123794 147234
rect 123962 147144 124438 147234
rect 124606 147144 125082 147234
rect 125250 147144 125726 147234
rect 125894 147144 126370 147234
rect 126538 147144 127014 147234
rect 127182 147144 127658 147234
rect 127826 147144 128302 147234
rect 128470 147144 128946 147234
rect 129114 147144 129590 147234
rect 129758 147144 130234 147234
rect 130402 147144 130970 147234
rect 131138 147144 131614 147234
rect 131782 147144 132258 147234
rect 132426 147144 132902 147234
rect 133070 147144 133546 147234
rect 133714 147144 134190 147234
rect 134358 147144 134834 147234
rect 135002 147144 135478 147234
rect 135646 147144 136122 147234
rect 136290 147144 136766 147234
rect 136934 147144 137410 147234
rect 137578 147144 138054 147234
rect 138222 147144 138698 147234
rect 138866 147144 139342 147234
rect 139510 147144 140078 147234
rect 140246 147144 140722 147234
rect 140890 147144 141366 147234
rect 141534 147144 142010 147234
rect 142178 147144 142654 147234
rect 142822 147144 143298 147234
rect 143466 147144 143942 147234
rect 144110 147144 144586 147234
rect 144754 147144 145230 147234
rect 145398 147144 145874 147234
rect 146042 147144 146518 147234
rect 146686 147144 147162 147234
rect 147330 147144 147806 147234
rect 147974 147144 148450 147234
rect 148618 147144 149186 147234
rect 149354 147144 149830 147234
rect 149998 147144 150474 147234
rect 150642 147144 151118 147234
rect 151286 147144 151762 147234
rect 151930 147144 152406 147234
rect 152574 147144 153050 147234
rect 153218 147144 153694 147234
rect 153862 147144 154338 147234
rect 154506 147144 154982 147234
rect 155150 147144 155626 147234
rect 155794 147144 156270 147234
rect 156438 147144 156914 147234
rect 157082 147144 157558 147234
rect 157726 147144 158202 147234
rect 158370 147144 158938 147234
rect 159106 147144 159582 147234
rect 159750 147144 160226 147234
rect 160394 147144 160870 147234
rect 161038 147144 161514 147234
rect 161682 147144 162158 147234
rect 162326 147144 162802 147234
rect 162970 147144 163446 147234
rect 163614 147144 164090 147234
rect 164258 147144 164734 147234
rect 164902 147144 165378 147234
rect 165546 147144 166022 147234
rect 166190 147144 166666 147234
rect 166834 147144 167310 147234
rect 167478 147144 168046 147234
rect 168214 147144 168690 147234
rect 168858 147144 169334 147234
rect 169502 147144 169978 147234
rect 170146 147144 170622 147234
rect 170790 147144 171266 147234
rect 171434 147144 171910 147234
rect 172078 147144 172554 147234
rect 172722 147144 173198 147234
rect 173366 147144 173842 147234
rect 174010 147144 174486 147234
rect 174654 147144 175130 147234
rect 175298 147144 175774 147234
rect 175942 147144 176418 147234
rect 176586 147144 177154 147234
rect 177322 147144 177798 147234
rect 177966 147144 178442 147234
rect 178610 147144 179086 147234
rect 179254 147144 179730 147234
rect 179898 147144 180374 147234
rect 180542 147144 181018 147234
rect 181186 147144 181662 147234
rect 181830 147144 182306 147234
rect 182474 147144 182950 147234
rect 183118 147144 183594 147234
rect 183762 147144 184238 147234
rect 184406 147144 184882 147234
rect 185050 147144 185526 147234
rect 185694 147144 186170 147234
rect 186338 147144 186906 147234
rect 187074 147144 187550 147234
rect 187718 147144 188194 147234
rect 188362 147144 188838 147234
rect 189006 147144 189482 147234
rect 189650 147144 190126 147234
rect 190294 147144 190770 147234
rect 190938 147144 191414 147234
rect 191582 147144 192058 147234
rect 192226 147144 192702 147234
rect 192870 147144 193346 147234
rect 193514 147144 193990 147234
rect 194158 147144 194634 147234
rect 194802 147144 195278 147234
rect 195446 147144 196014 147234
rect 196182 147144 196658 147234
rect 196826 147144 197302 147234
rect 197470 147144 197946 147234
rect 198114 147144 198590 147234
rect 198758 147144 199234 147234
rect 199402 147144 199878 147234
rect 200046 147144 200522 147234
rect 200690 147144 201166 147234
rect 201334 147144 201810 147234
rect 201978 147144 202454 147234
rect 202622 147144 203098 147234
rect 203266 147144 203742 147234
rect 203910 147144 204386 147234
rect 204554 147144 205122 147234
rect 205290 147144 205766 147234
rect 205934 147144 206410 147234
rect 206578 147144 207054 147234
rect 207222 147144 207698 147234
rect 207866 147144 208342 147234
rect 208510 147144 208986 147234
rect 209154 147144 209630 147234
rect 209798 147144 210274 147234
rect 210442 147144 210918 147234
rect 211086 147144 211562 147234
rect 211730 147144 212206 147234
rect 212374 147144 212850 147234
rect 213018 147144 213494 147234
rect 213662 147144 214230 147234
rect 214398 147144 214874 147234
rect 215042 147144 215518 147234
rect 215686 147144 216162 147234
rect 216330 147144 216806 147234
rect 216974 147144 217450 147234
rect 217618 147144 218094 147234
rect 218262 147144 218738 147234
rect 218906 147144 219382 147234
rect 219550 147144 220026 147234
rect 220194 147144 220670 147234
rect 220838 147144 221314 147234
rect 221482 147144 221958 147234
rect 222126 147144 222602 147234
rect 222770 147144 223246 147234
rect 223414 147144 223982 147234
rect 224150 147144 224626 147234
rect 224794 147144 225270 147234
rect 225438 147144 225914 147234
rect 226082 147144 226558 147234
rect 226726 147144 227202 147234
rect 227370 147144 227846 147234
rect 228014 147144 228490 147234
rect 228658 147144 229134 147234
rect 229302 147144 229778 147234
rect 229946 147144 230422 147234
rect 230590 147144 231066 147234
rect 231234 147144 231710 147234
rect 231878 147144 232354 147234
rect 232522 147144 233090 147234
rect 233258 147144 233734 147234
rect 233902 147144 234378 147234
rect 234546 147144 235022 147234
rect 235190 147144 235666 147234
rect 235834 147144 236310 147234
rect 236478 147144 236954 147234
rect 237122 147144 237598 147234
rect 237766 147144 238242 147234
rect 238410 147144 238886 147234
rect 239054 147144 239530 147234
rect 239698 147144 240174 147234
rect 240342 147144 240818 147234
rect 240986 147144 241462 147234
rect 241630 147144 242198 147234
rect 242366 147144 242842 147234
rect 243010 147144 243486 147234
rect 243654 147144 244130 147234
rect 244298 147144 244774 147234
rect 244942 147144 245418 147234
rect 245586 147144 246062 147234
rect 246230 147144 246706 147234
rect 246874 147144 247350 147234
rect 247518 147144 247994 147234
rect 248162 147144 248638 147234
rect 248806 147144 249282 147234
rect 249450 147144 249926 147234
rect 250094 147144 250570 147234
rect 250738 147144 251214 147234
rect 251382 147144 251950 147234
rect 252118 147144 252594 147234
rect 252762 147144 253238 147234
rect 253406 147144 253882 147234
rect 254050 147144 254526 147234
rect 254694 147144 255170 147234
rect 255338 147144 255814 147234
rect 255982 147144 256458 147234
rect 256626 147144 257102 147234
rect 257270 147144 257746 147234
rect 257914 147144 258390 147234
rect 258558 147144 259034 147234
rect 259202 147144 259678 147234
rect 259846 147144 260322 147234
rect 260490 147144 261058 147234
rect 261226 147144 261702 147234
rect 261870 147144 262346 147234
rect 262514 147144 262990 147234
rect 263158 147144 263634 147234
rect 263802 147144 264278 147234
rect 264446 147144 264922 147234
rect 265090 147144 265566 147234
rect 265734 147144 266210 147234
rect 266378 147144 266854 147234
rect 267022 147144 267498 147234
rect 267666 147144 268142 147234
rect 268310 147144 268786 147234
rect 268954 147144 269430 147234
rect 269598 147144 270166 147234
rect 270334 147144 270810 147234
rect 270978 147144 271454 147234
rect 271622 147144 272098 147234
rect 272266 147144 272742 147234
rect 272910 147144 273386 147234
rect 273554 147144 274030 147234
rect 274198 147144 274674 147234
rect 274842 147144 275318 147234
rect 275486 147144 275962 147234
rect 276130 147144 276606 147234
rect 276774 147144 277250 147234
rect 277418 147144 277894 147234
rect 278062 147144 278538 147234
rect 278706 147144 279182 147234
rect 279350 147144 279918 147234
rect 280086 147144 280562 147234
rect 280730 147144 281206 147234
rect 281374 147144 281850 147234
rect 282018 147144 282494 147234
rect 282662 147144 283138 147234
rect 283306 147144 283782 147234
rect 283950 147144 284426 147234
rect 284594 147144 285070 147234
rect 285238 147144 285714 147234
rect 285882 147144 286358 147234
rect 286526 147144 287002 147234
rect 287170 147144 287646 147234
rect 287814 147144 288290 147234
rect 288458 147144 289026 147234
rect 289194 147144 289670 147234
rect 289838 147144 290314 147234
rect 290482 147144 290958 147234
rect 291126 147144 291602 147234
rect 291770 147144 292246 147234
rect 292414 147144 292890 147234
rect 293058 147144 293534 147234
rect 293702 147144 294178 147234
rect 294346 147144 294822 147234
rect 294990 147144 295466 147234
rect 295634 147144 296110 147234
rect 296278 147144 296754 147234
rect 296922 147144 297398 147234
rect 297566 147144 298134 147234
rect 298302 147144 298778 147234
rect 298946 147144 299422 147234
rect 299590 147144 300066 147234
rect 300234 147144 300710 147234
rect 300878 147144 301354 147234
rect 301522 147144 301998 147234
rect 302166 147144 302642 147234
rect 302810 147144 303286 147234
rect 303454 147144 303930 147234
rect 304098 147144 304574 147234
rect 304742 147144 305218 147234
rect 305386 147144 305862 147234
rect 306030 147144 306506 147234
rect 306674 147144 307242 147234
rect 307410 147144 307886 147234
rect 308054 147144 308530 147234
rect 308698 147144 309174 147234
rect 309342 147144 309818 147234
rect 309986 147144 310462 147234
rect 310630 147144 311106 147234
rect 311274 147144 311750 147234
rect 311918 147144 312394 147234
rect 312562 147144 313038 147234
rect 313206 147144 313682 147234
rect 313850 147144 314326 147234
rect 314494 147144 314970 147234
rect 315138 147144 315614 147234
rect 315782 147144 316258 147234
rect 316426 147144 316994 147234
rect 317162 147144 317638 147234
rect 317806 147144 318282 147234
rect 318450 147144 318926 147234
rect 319094 147144 319570 147234
rect 319738 147144 320214 147234
rect 320382 147144 320858 147234
rect 321026 147144 321502 147234
rect 321670 147144 322146 147234
rect 322314 147144 322790 147234
rect 322958 147144 323434 147234
rect 323602 147144 324078 147234
rect 324246 147144 324722 147234
rect 324890 147144 325366 147234
rect 325534 147144 326102 147234
rect 326270 147144 326746 147234
rect 326914 147144 327390 147234
rect 327558 147144 328034 147234
rect 328202 147144 328678 147234
rect 328846 147144 329322 147234
rect 329490 147144 329966 147234
rect 330134 147144 330610 147234
rect 330778 147144 331254 147234
rect 331422 147144 331898 147234
rect 332066 147144 332542 147234
rect 332710 147144 333186 147234
rect 333354 147144 333830 147234
rect 333998 147144 334474 147234
rect 334642 147144 335210 147234
rect 335378 147144 335854 147234
rect 336022 147144 336498 147234
rect 336666 147144 337142 147234
rect 337310 147144 337786 147234
rect 337954 147144 338430 147234
rect 338598 147144 339074 147234
rect 339242 147144 339718 147234
rect 339886 147144 340362 147234
rect 340530 147144 341006 147234
rect 341174 147144 341650 147234
rect 341818 147144 342294 147234
rect 342462 147144 342938 147234
rect 343106 147144 343582 147234
rect 343750 147144 344226 147234
rect 344394 147144 344962 147234
rect 345130 147144 345606 147234
rect 345774 147144 346250 147234
rect 346418 147144 346894 147234
rect 347062 147144 347538 147234
rect 347706 147144 348182 147234
rect 348350 147144 348826 147234
rect 348994 147144 349470 147234
rect 349638 147144 350114 147234
rect 350282 147144 350758 147234
rect 350926 147144 351402 147234
rect 351570 147144 352046 147234
rect 352214 147144 352690 147234
rect 352858 147144 353334 147234
rect 353502 147144 354070 147234
rect 354238 147144 354714 147234
rect 354882 147144 355358 147234
rect 355526 147144 356002 147234
rect 356170 147144 356646 147234
rect 356814 147144 357290 147234
rect 357458 147144 357934 147234
rect 358102 147144 358578 147234
rect 358746 147144 359222 147234
rect 359390 147144 359866 147234
rect 360034 147144 360510 147234
rect 360678 147144 361154 147234
rect 361322 147144 361798 147234
rect 361966 147144 362442 147234
rect 362610 147144 363178 147234
rect 363346 147144 363822 147234
rect 363990 147144 364466 147234
rect 364634 147144 365110 147234
rect 365278 147144 365754 147234
rect 365922 147144 366398 147234
rect 366566 147144 367042 147234
rect 367210 147144 367686 147234
rect 367854 147144 368330 147234
rect 368498 147144 368974 147234
rect 369142 147144 369618 147234
rect 369786 147144 370262 147234
rect 370430 147144 370906 147234
rect 371074 147144 371550 147234
rect 371718 147144 372194 147234
rect 372362 147144 372930 147234
rect 373098 147144 373574 147234
rect 373742 147144 374218 147234
rect 374386 147144 374862 147234
rect 375030 147144 375506 147234
rect 375674 147144 376150 147234
rect 376318 147144 376794 147234
rect 376962 147144 377438 147234
rect 377606 147144 378082 147234
rect 378250 147144 378726 147234
rect 378894 147144 379370 147234
rect 379538 147144 380014 147234
rect 380182 147144 380658 147234
rect 380826 147144 381302 147234
rect 381470 147144 382038 147234
rect 382206 147144 382682 147234
rect 382850 147144 383326 147234
rect 383494 147144 383970 147234
rect 384138 147144 384614 147234
rect 384782 147144 385258 147234
rect 385426 147144 385902 147234
rect 386070 147144 386546 147234
rect 386714 147144 387190 147234
rect 387358 147144 387834 147234
rect 388002 147144 388478 147234
rect 388646 147144 389122 147234
rect 389290 147144 389766 147234
rect 389934 147144 390410 147234
rect 390578 147144 391146 147234
rect 391314 147144 391790 147234
rect 391958 147144 392434 147234
rect 392602 147144 393078 147234
rect 393246 147144 393722 147234
rect 393890 147144 394366 147234
rect 394534 147144 395010 147234
rect 395178 147144 395654 147234
rect 395822 147144 396298 147234
rect 396466 147144 396942 147234
rect 397110 147144 397586 147234
rect 397754 147144 398230 147234
rect 398398 147144 398874 147234
rect 399042 147144 399518 147234
rect 296 856 399628 147144
rect 296 734 1618 856
rect 1786 734 4930 856
rect 5098 734 8334 856
rect 8502 734 11646 856
rect 11814 734 15050 856
rect 15218 734 18362 856
rect 18530 734 21766 856
rect 21934 734 25078 856
rect 25246 734 28482 856
rect 28650 734 31794 856
rect 31962 734 35198 856
rect 35366 734 38510 856
rect 38678 734 41914 856
rect 42082 734 45226 856
rect 45394 734 48630 856
rect 48798 734 52034 856
rect 52202 734 55346 856
rect 55514 734 58750 856
rect 58918 734 62062 856
rect 62230 734 65466 856
rect 65634 734 68778 856
rect 68946 734 72182 856
rect 72350 734 75494 856
rect 75662 734 78898 856
rect 79066 734 82210 856
rect 82378 734 85614 856
rect 85782 734 88926 856
rect 89094 734 92330 856
rect 92498 734 95734 856
rect 95902 734 99046 856
rect 99214 734 102450 856
rect 102618 734 105762 856
rect 105930 734 109166 856
rect 109334 734 112478 856
rect 112646 734 115882 856
rect 116050 734 119194 856
rect 119362 734 122598 856
rect 122766 734 125910 856
rect 126078 734 129314 856
rect 129482 734 132626 856
rect 132794 734 136030 856
rect 136198 734 139434 856
rect 139602 734 142746 856
rect 142914 734 146150 856
rect 146318 734 149462 856
rect 149630 734 152866 856
rect 153034 734 156178 856
rect 156346 734 159582 856
rect 159750 734 162894 856
rect 163062 734 166298 856
rect 166466 734 169610 856
rect 169778 734 173014 856
rect 173182 734 176326 856
rect 176494 734 179730 856
rect 179898 734 183134 856
rect 183302 734 186446 856
rect 186614 734 189850 856
rect 190018 734 193162 856
rect 193330 734 196566 856
rect 196734 734 199878 856
rect 200046 734 203282 856
rect 203450 734 206594 856
rect 206762 734 209998 856
rect 210166 734 213310 856
rect 213478 734 216714 856
rect 216882 734 220026 856
rect 220194 734 223430 856
rect 223598 734 226834 856
rect 227002 734 230146 856
rect 230314 734 233550 856
rect 233718 734 236862 856
rect 237030 734 240266 856
rect 240434 734 243578 856
rect 243746 734 246982 856
rect 247150 734 250294 856
rect 250462 734 253698 856
rect 253866 734 257010 856
rect 257178 734 260414 856
rect 260582 734 263726 856
rect 263894 734 267130 856
rect 267298 734 270534 856
rect 270702 734 273846 856
rect 274014 734 277250 856
rect 277418 734 280562 856
rect 280730 734 283966 856
rect 284134 734 287278 856
rect 287446 734 290682 856
rect 290850 734 293994 856
rect 294162 734 297398 856
rect 297566 734 300710 856
rect 300878 734 304114 856
rect 304282 734 307426 856
rect 307594 734 310830 856
rect 310998 734 314234 856
rect 314402 734 317546 856
rect 317714 734 320950 856
rect 321118 734 324262 856
rect 324430 734 327666 856
rect 327834 734 330978 856
rect 331146 734 334382 856
rect 334550 734 337694 856
rect 337862 734 341098 856
rect 341266 734 344410 856
rect 344578 734 347814 856
rect 347982 734 351126 856
rect 351294 734 354530 856
rect 354698 734 357934 856
rect 358102 734 361246 856
rect 361414 734 364650 856
rect 364818 734 367962 856
rect 368130 734 371366 856
rect 371534 734 374678 856
rect 374846 734 378082 856
rect 378250 734 381394 856
rect 381562 734 384798 856
rect 384966 734 388110 856
rect 388278 734 391514 856
rect 391682 734 394826 856
rect 394994 734 398230 856
rect 398398 734 399628 856
<< metal3 >>
rect 0 146616 800 146736
rect 399200 144440 400000 144560
rect 0 144168 800 144288
rect 0 141720 800 141840
rect 0 139272 800 139392
rect 399200 137776 400000 137896
rect 0 136824 800 136944
rect 0 134376 800 134496
rect 0 132064 800 132184
rect 399200 130976 400000 131096
rect 0 129616 800 129736
rect 0 127168 800 127288
rect 0 124720 800 124840
rect 399200 124312 400000 124432
rect 0 122272 800 122392
rect 0 119824 800 119944
rect 0 117512 800 117632
rect 399200 117512 400000 117632
rect 0 115064 800 115184
rect 0 112616 800 112736
rect 399200 110848 400000 110968
rect 0 110168 800 110288
rect 0 107720 800 107840
rect 0 105272 800 105392
rect 399200 104048 400000 104168
rect 0 102960 800 103080
rect 0 100512 800 100632
rect 0 98064 800 98184
rect 399200 97384 400000 97504
rect 0 95616 800 95736
rect 0 93168 800 93288
rect 0 90720 800 90840
rect 399200 90584 400000 90704
rect 0 88408 800 88528
rect 0 85960 800 86080
rect 399200 83920 400000 84040
rect 0 83512 800 83632
rect 0 81064 800 81184
rect 0 78616 800 78736
rect 399200 77256 400000 77376
rect 0 76168 800 76288
rect 0 73856 800 73976
rect 0 71408 800 71528
rect 399200 70456 400000 70576
rect 0 68960 800 69080
rect 0 66512 800 66632
rect 0 64064 800 64184
rect 399200 63792 400000 63912
rect 0 61616 800 61736
rect 0 59304 800 59424
rect 0 56856 800 56976
rect 399200 56992 400000 57112
rect 0 54408 800 54528
rect 0 51960 800 52080
rect 399200 50328 400000 50448
rect 0 49512 800 49632
rect 0 47064 800 47184
rect 0 44752 800 44872
rect 399200 43528 400000 43648
rect 0 42304 800 42424
rect 0 39856 800 39976
rect 0 37408 800 37528
rect 399200 36864 400000 36984
rect 0 34960 800 35080
rect 0 32512 800 32632
rect 0 30200 800 30320
rect 399200 30064 400000 30184
rect 0 27752 800 27872
rect 0 25304 800 25424
rect 399200 23400 400000 23520
rect 0 22856 800 22976
rect 0 20408 800 20528
rect 0 17960 800 18080
rect 399200 16600 400000 16720
rect 0 15648 800 15768
rect 0 13200 800 13320
rect 0 10752 800 10872
rect 399200 9936 400000 10056
rect 0 8304 800 8424
rect 0 5856 800 5976
rect 0 3408 800 3528
rect 399200 3272 400000 3392
rect 0 1096 800 1216
<< obsm3 >>
rect 880 146536 399200 146709
rect 800 144640 399200 146536
rect 800 144368 399120 144640
rect 880 144360 399120 144368
rect 880 144088 399200 144360
rect 800 141920 399200 144088
rect 880 141640 399200 141920
rect 800 139472 399200 141640
rect 880 139192 399200 139472
rect 800 137976 399200 139192
rect 800 137696 399120 137976
rect 800 137024 399200 137696
rect 880 136744 399200 137024
rect 800 134576 399200 136744
rect 880 134296 399200 134576
rect 800 132264 399200 134296
rect 880 131984 399200 132264
rect 800 131176 399200 131984
rect 800 130896 399120 131176
rect 800 129816 399200 130896
rect 880 129536 399200 129816
rect 800 127368 399200 129536
rect 880 127088 399200 127368
rect 800 124920 399200 127088
rect 880 124640 399200 124920
rect 800 124512 399200 124640
rect 800 124232 399120 124512
rect 800 122472 399200 124232
rect 880 122192 399200 122472
rect 800 120024 399200 122192
rect 880 119744 399200 120024
rect 800 117712 399200 119744
rect 880 117432 399120 117712
rect 800 115264 399200 117432
rect 880 114984 399200 115264
rect 800 112816 399200 114984
rect 880 112536 399200 112816
rect 800 111048 399200 112536
rect 800 110768 399120 111048
rect 800 110368 399200 110768
rect 880 110088 399200 110368
rect 800 107920 399200 110088
rect 880 107640 399200 107920
rect 800 105472 399200 107640
rect 880 105192 399200 105472
rect 800 104248 399200 105192
rect 800 103968 399120 104248
rect 800 103160 399200 103968
rect 880 102880 399200 103160
rect 800 100712 399200 102880
rect 880 100432 399200 100712
rect 800 98264 399200 100432
rect 880 97984 399200 98264
rect 800 97584 399200 97984
rect 800 97304 399120 97584
rect 800 95816 399200 97304
rect 880 95536 399200 95816
rect 800 93368 399200 95536
rect 880 93088 399200 93368
rect 800 90920 399200 93088
rect 880 90784 399200 90920
rect 880 90640 399120 90784
rect 800 90504 399120 90640
rect 800 88608 399200 90504
rect 880 88328 399200 88608
rect 800 86160 399200 88328
rect 880 85880 399200 86160
rect 800 84120 399200 85880
rect 800 83840 399120 84120
rect 800 83712 399200 83840
rect 880 83432 399200 83712
rect 800 81264 399200 83432
rect 880 80984 399200 81264
rect 800 78816 399200 80984
rect 880 78536 399200 78816
rect 800 77456 399200 78536
rect 800 77176 399120 77456
rect 800 76368 399200 77176
rect 880 76088 399200 76368
rect 800 74056 399200 76088
rect 880 73776 399200 74056
rect 800 71608 399200 73776
rect 880 71328 399200 71608
rect 800 70656 399200 71328
rect 800 70376 399120 70656
rect 800 69160 399200 70376
rect 880 68880 399200 69160
rect 800 66712 399200 68880
rect 880 66432 399200 66712
rect 800 64264 399200 66432
rect 880 63992 399200 64264
rect 880 63984 399120 63992
rect 800 63712 399120 63984
rect 800 61816 399200 63712
rect 880 61536 399200 61816
rect 800 59504 399200 61536
rect 880 59224 399200 59504
rect 800 57192 399200 59224
rect 800 57056 399120 57192
rect 880 56912 399120 57056
rect 880 56776 399200 56912
rect 800 54608 399200 56776
rect 880 54328 399200 54608
rect 800 52160 399200 54328
rect 880 51880 399200 52160
rect 800 50528 399200 51880
rect 800 50248 399120 50528
rect 800 49712 399200 50248
rect 880 49432 399200 49712
rect 800 47264 399200 49432
rect 880 46984 399200 47264
rect 800 44952 399200 46984
rect 880 44672 399200 44952
rect 800 43728 399200 44672
rect 800 43448 399120 43728
rect 800 42504 399200 43448
rect 880 42224 399200 42504
rect 800 40056 399200 42224
rect 880 39776 399200 40056
rect 800 37608 399200 39776
rect 880 37328 399200 37608
rect 800 37064 399200 37328
rect 800 36784 399120 37064
rect 800 35160 399200 36784
rect 880 34880 399200 35160
rect 800 32712 399200 34880
rect 880 32432 399200 32712
rect 800 30400 399200 32432
rect 880 30264 399200 30400
rect 880 30120 399120 30264
rect 800 29984 399120 30120
rect 800 27952 399200 29984
rect 880 27672 399200 27952
rect 800 25504 399200 27672
rect 880 25224 399200 25504
rect 800 23600 399200 25224
rect 800 23320 399120 23600
rect 800 23056 399200 23320
rect 880 22776 399200 23056
rect 800 20608 399200 22776
rect 880 20328 399200 20608
rect 800 18160 399200 20328
rect 880 17880 399200 18160
rect 800 16800 399200 17880
rect 800 16520 399120 16800
rect 800 15848 399200 16520
rect 880 15568 399200 15848
rect 800 13400 399200 15568
rect 880 13120 399200 13400
rect 800 10952 399200 13120
rect 880 10672 399200 10952
rect 800 10136 399200 10672
rect 800 9856 399120 10136
rect 800 8504 399200 9856
rect 880 8224 399200 8504
rect 800 6056 399200 8224
rect 880 5776 399200 6056
rect 800 3608 399200 5776
rect 880 3472 399200 3608
rect 880 3328 399120 3472
rect 800 3192 399120 3328
rect 800 1296 399200 3192
rect 880 1123 399200 1296
<< metal4 >>
rect 4 156 324 147812
rect 664 816 984 147152
rect 5128 156 5448 147812
rect 10128 156 10448 147812
rect 15128 156 15448 147812
rect 20128 107460 20448 147812
rect 25128 107460 25448 147812
rect 30128 107460 30448 147812
rect 35128 107460 35448 147812
rect 40128 107460 40448 147812
rect 45128 107460 45448 147812
rect 50128 107460 50448 147812
rect 55128 107460 55448 147812
rect 60128 107460 60448 147812
rect 65128 107460 65448 147812
rect 70128 107460 70448 147812
rect 75128 107460 75448 147812
rect 80128 107460 80448 147812
rect 85128 107460 85448 147812
rect 90128 107460 90448 147812
rect 95128 107460 95448 147812
rect 100128 107460 100448 147812
rect 105128 107460 105448 147812
rect 110128 107460 110448 147812
rect 115128 107460 115448 147812
rect 120128 107460 120448 147812
rect 125128 107460 125448 147812
rect 130128 107460 130448 147812
rect 135128 107460 135448 147812
rect 140128 107460 140448 147812
rect 145128 107460 145448 147812
rect 150128 107460 150448 147812
rect 155128 107460 155448 147812
rect 20128 156 20448 20248
rect 25128 156 25448 20248
rect 30128 156 30448 20248
rect 35128 156 35448 20248
rect 40128 156 40448 20248
rect 45128 156 45448 20248
rect 50128 156 50448 20248
rect 55128 156 55448 20248
rect 60128 156 60448 20248
rect 65128 156 65448 20248
rect 70128 156 70448 20248
rect 75128 156 75448 20248
rect 80128 156 80448 20248
rect 85128 156 85448 20248
rect 90128 156 90448 20248
rect 95128 156 95448 20248
rect 100128 156 100448 20248
rect 105128 156 105448 20248
rect 110128 156 110448 20248
rect 115128 156 115448 20248
rect 120128 156 120448 20248
rect 125128 156 125448 20248
rect 130128 156 130448 20248
rect 135128 156 135448 20248
rect 140128 156 140448 20248
rect 145128 156 145448 20248
rect 150128 156 150448 20248
rect 155128 156 155448 20248
rect 160128 156 160448 147812
rect 165128 156 165448 147812
rect 170128 156 170448 147812
rect 175128 156 175448 147812
rect 180128 156 180448 147812
rect 185128 156 185448 147812
rect 190128 156 190448 147812
rect 195128 156 195448 147812
rect 200128 156 200448 147812
rect 205128 156 205448 147812
rect 210128 156 210448 147812
rect 215128 156 215448 147812
rect 220128 156 220448 147812
rect 225128 156 225448 147812
rect 230128 156 230448 147812
rect 235128 156 235448 147812
rect 240128 156 240448 147812
rect 245128 156 245448 147812
rect 250128 156 250448 147812
rect 255128 156 255448 147812
rect 260128 156 260448 147812
rect 265128 156 265448 147812
rect 270128 156 270448 147812
rect 275128 156 275448 147812
rect 280128 156 280448 147812
rect 285128 156 285448 147812
rect 290128 156 290448 147812
rect 295128 156 295448 147812
rect 300128 156 300448 147812
rect 305128 156 305448 147812
rect 310128 156 310448 147812
rect 315128 156 315448 147812
rect 320128 156 320448 147812
rect 325128 156 325448 147812
rect 330128 156 330448 147812
rect 335128 156 335448 147812
rect 340128 156 340448 147812
rect 345128 156 345448 147812
rect 350128 156 350448 147812
rect 355128 156 355448 147812
rect 360128 156 360448 147812
rect 365128 156 365448 147812
rect 370128 156 370448 147812
rect 375128 156 375448 147812
rect 380128 156 380448 147812
rect 385128 156 385448 147812
rect 390128 156 390448 147812
rect 395128 156 395448 147812
rect 398940 816 399260 147152
rect 399600 156 399920 147812
<< obsm4 >>
rect 3654 2347 5048 144669
rect 5528 2347 10048 144669
rect 10528 2347 15048 144669
rect 15528 107380 20048 144669
rect 20528 107380 25048 144669
rect 25528 107380 30048 144669
rect 30528 107380 35048 144669
rect 35528 107380 40048 144669
rect 40528 107380 45048 144669
rect 45528 107380 50048 144669
rect 50528 107380 55048 144669
rect 55528 107380 60048 144669
rect 60528 107380 65048 144669
rect 65528 107380 70048 144669
rect 70528 107380 75048 144669
rect 75528 107380 80048 144669
rect 80528 107380 85048 144669
rect 85528 107380 90048 144669
rect 90528 107380 95048 144669
rect 95528 107380 100048 144669
rect 100528 107380 105048 144669
rect 105528 107380 110048 144669
rect 110528 107380 115048 144669
rect 115528 107380 120048 144669
rect 120528 107380 125048 144669
rect 125528 107380 130048 144669
rect 130528 107380 135048 144669
rect 135528 107380 140048 144669
rect 140528 107380 145048 144669
rect 145528 107380 150048 144669
rect 150528 107380 155048 144669
rect 155528 107380 160048 144669
rect 15528 20328 160048 107380
rect 15528 2347 20048 20328
rect 20528 2347 25048 20328
rect 25528 2347 30048 20328
rect 30528 2347 35048 20328
rect 35528 2347 40048 20328
rect 40528 2347 45048 20328
rect 45528 2347 50048 20328
rect 50528 2347 55048 20328
rect 55528 2347 60048 20328
rect 60528 2347 65048 20328
rect 65528 2347 70048 20328
rect 70528 2347 75048 20328
rect 75528 2347 80048 20328
rect 80528 2347 85048 20328
rect 85528 2347 90048 20328
rect 90528 2347 95048 20328
rect 95528 2347 100048 20328
rect 100528 2347 105048 20328
rect 105528 2347 110048 20328
rect 110528 2347 115048 20328
rect 115528 2347 120048 20328
rect 120528 2347 125048 20328
rect 125528 2347 130048 20328
rect 130528 2347 135048 20328
rect 135528 2347 140048 20328
rect 140528 2347 145048 20328
rect 145528 2347 150048 20328
rect 150528 2347 155048 20328
rect 155528 2347 160048 20328
rect 160528 2347 165048 144669
rect 165528 2347 170048 144669
rect 170528 2347 175048 144669
rect 175528 2347 180048 144669
rect 180528 2347 185048 144669
rect 185528 2347 190048 144669
rect 190528 2347 195048 144669
rect 195528 2347 200048 144669
rect 200528 2347 205048 144669
rect 205528 2347 210048 144669
rect 210528 2347 215048 144669
rect 215528 2347 220048 144669
rect 220528 2347 225048 144669
rect 225528 2347 230048 144669
rect 230528 2347 235048 144669
rect 235528 2347 240048 144669
rect 240528 2347 245048 144669
rect 245528 2347 250048 144669
rect 250528 2347 255048 144669
rect 255528 2347 260048 144669
rect 260528 2347 265048 144669
rect 265528 2347 270048 144669
rect 270528 2347 275048 144669
rect 275528 2347 280048 144669
rect 280528 2347 285048 144669
rect 285528 2347 290048 144669
rect 290528 2347 295048 144669
rect 295528 2347 300048 144669
rect 300528 2347 305048 144669
rect 305528 2347 310048 144669
rect 310528 2347 315048 144669
rect 315528 2347 320048 144669
rect 320528 2347 325048 144669
rect 325528 2347 330048 144669
rect 330528 2347 335048 144669
rect 335528 2347 340048 144669
rect 340528 2347 345048 144669
rect 345528 2347 350048 144669
rect 350528 2347 355048 144669
rect 355528 2347 356165 144669
<< metal5 >>
rect 4 147492 399920 147812
rect 664 146832 399260 147152
rect 4 135298 399920 135618
rect 4 122298 399920 122618
rect 4 109298 399920 109618
rect 4 96298 399920 96618
rect 4 83298 399920 83618
rect 4 70298 399920 70618
rect 4 57298 399920 57618
rect 4 44298 399920 44618
rect 4 31298 399920 31618
rect 4 18298 399920 18618
rect 4 5298 399920 5618
rect 664 816 399260 1136
rect 4 156 399920 476
<< obsm5 >>
rect 3612 135938 272572 143300
rect 3612 122938 272572 134978
rect 3612 109938 272572 121978
rect 3612 96938 272572 108978
rect 3612 83938 272572 95978
rect 3612 70938 272572 82978
rect 3612 57938 272572 69978
rect 3612 44938 272572 56978
rect 3612 31938 272572 43978
rect 3612 21940 272572 30978
<< labels >>
rlabel metal5 s 4 156 399920 476 6 VGND
port 1 nsew ground input
rlabel metal5 s 4 18298 399920 18618 6 VGND
port 1 nsew ground input
rlabel metal5 s 4 44298 399920 44618 6 VGND
port 1 nsew ground input
rlabel metal5 s 4 70298 399920 70618 6 VGND
port 1 nsew ground input
rlabel metal5 s 4 96298 399920 96618 6 VGND
port 1 nsew ground input
rlabel metal5 s 4 122298 399920 122618 6 VGND
port 1 nsew ground input
rlabel metal5 s 4 147492 399920 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 20128 156 20448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 30128 156 30448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 40128 156 40448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 50128 156 50448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 60128 156 60448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 70128 156 70448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 80128 156 80448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 90128 156 90448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 100128 156 100448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 110128 156 110448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 120128 156 120448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 130128 156 130448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 140128 156 140448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 150128 156 150448 20248 6 VGND
port 1 nsew ground input
rlabel metal4 s 4 156 324 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 10128 156 10448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 20128 107460 20448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 30128 107460 30448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 40128 107460 40448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 50128 107460 50448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 60128 107460 60448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 70128 107460 70448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 80128 107460 80448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 90128 107460 90448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 100128 107460 100448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 110128 107460 110448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 120128 107460 120448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 130128 107460 130448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 140128 107460 140448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 150128 107460 150448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 160128 156 160448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 170128 156 170448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 180128 156 180448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 190128 156 190448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 200128 156 200448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 210128 156 210448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 220128 156 220448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 230128 156 230448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 240128 156 240448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 250128 156 250448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 260128 156 260448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 270128 156 270448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 280128 156 280448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 290128 156 290448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 300128 156 300448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 310128 156 310448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 320128 156 320448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 330128 156 330448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 340128 156 340448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 350128 156 350448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 360128 156 360448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 370128 156 370448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 380128 156 380448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 390128 156 390448 147812 6 VGND
port 1 nsew ground input
rlabel metal4 s 399600 156 399920 147812 6 VGND
port 1 nsew ground input
rlabel metal5 s 664 816 399260 1136 6 VPWR
port 2 nsew power input
rlabel metal5 s 4 5298 399920 5618 6 VPWR
port 2 nsew power input
rlabel metal5 s 4 31298 399920 31618 6 VPWR
port 2 nsew power input
rlabel metal5 s 4 57298 399920 57618 6 VPWR
port 2 nsew power input
rlabel metal5 s 4 83298 399920 83618 6 VPWR
port 2 nsew power input
rlabel metal5 s 4 109298 399920 109618 6 VPWR
port 2 nsew power input
rlabel metal5 s 4 135298 399920 135618 6 VPWR
port 2 nsew power input
rlabel metal5 s 664 146832 399260 147152 6 VPWR
port 2 nsew power input
rlabel metal4 s 25128 156 25448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 35128 156 35448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 45128 156 45448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 55128 156 55448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 65128 156 65448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 75128 156 75448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 85128 156 85448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 95128 156 95448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 105128 156 105448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 115128 156 115448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 125128 156 125448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 135128 156 135448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 145128 156 145448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 155128 156 155448 20248 6 VPWR
port 2 nsew power input
rlabel metal4 s 664 816 984 147152 6 VPWR
port 2 nsew power input
rlabel metal4 s 398940 816 399260 147152 6 VPWR
port 2 nsew power input
rlabel metal4 s 5128 156 5448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 15128 156 15448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 25128 107460 25448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 35128 107460 35448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 45128 107460 45448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 55128 107460 55448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 65128 107460 65448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 75128 107460 75448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 85128 107460 85448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 95128 107460 95448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 105128 107460 105448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 115128 107460 115448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 125128 107460 125448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 135128 107460 135448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 145128 107460 145448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 155128 107460 155448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 165128 156 165448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 175128 156 175448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 185128 156 185448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 195128 156 195448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 205128 156 205448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 215128 156 215448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 225128 156 225448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 235128 156 235448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 245128 156 245448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 255128 156 255448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 265128 156 265448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 275128 156 275448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 285128 156 285448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 295128 156 295448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 305128 156 305448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 315128 156 315448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 325128 156 325448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 335128 156 335448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 345128 156 345448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 355128 156 355448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 365128 156 365448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 375128 156 375448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 385128 156 385448 147812 6 VPWR
port 2 nsew power input
rlabel metal4 s 395128 156 395448 147812 6 VPWR
port 2 nsew power input
rlabel metal2 s 294 147200 350 148000 6 core_clk
port 3 nsew signal input
rlabel metal2 s 938 147200 994 148000 6 core_rstn
port 4 nsew signal input
rlabel metal2 s 317602 0 317658 800 6 debug_mode
port 5 nsew signal output
rlabel metal2 s 321006 0 321062 800 6 debug_oeb
port 6 nsew signal output
rlabel metal2 s 383382 147200 383438 148000 6 debug_rx
port 7 nsew signal input
rlabel metal3 s 0 85960 800 86080 6 debug_tx
port 8 nsew signal output
rlabel metal2 s 21822 0 21878 800 6 flash_clk
port 9 nsew signal output
rlabel metal2 s 337750 0 337806 800 6 flash_cs_n
port 10 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 flash_io0_di
port 11 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 flash_io0_do
port 12 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 flash_io0_oeb
port 13 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 flash_io1_di
port 14 nsew signal input
rlabel metal2 s 38566 0 38622 800 6 flash_io1_do
port 15 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 flash_io1_oeb
port 16 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 flash_io2_di
port 17 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 flash_io2_do
port 18 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 flash_io2_oeb
port 19 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 flash_io3_di
port 20 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 flash_io3_do
port 21 nsew signal output
rlabel metal3 s 0 1096 800 1216 6 flash_io3_oeb
port 22 nsew signal output
rlabel metal2 s 1674 0 1730 800 6 gpio_in_pad
port 23 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 gpio_inenb_pad
port 24 nsew signal output
rlabel metal2 s 8390 0 8446 800 6 gpio_mode0_pad
port 25 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 gpio_mode1_pad
port 26 nsew signal output
rlabel metal2 s 15106 0 15162 800 6 gpio_out_pad
port 27 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 gpio_outenb_pad
port 28 nsew signal output
rlabel metal2 s 62118 0 62174 800 6 hk_ack_i
port 29 nsew signal input
rlabel metal2 s 384026 147200 384082 148000 6 hk_cyc_o
port 30 nsew signal output
rlabel metal2 s 68834 0 68890 800 6 hk_dat_i[0]
port 31 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 hk_dat_i[10]
port 32 nsew signal input
rlabel metal2 s 105818 0 105874 800 6 hk_dat_i[11]
port 33 nsew signal input
rlabel metal2 s 109222 0 109278 800 6 hk_dat_i[12]
port 34 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 hk_dat_i[13]
port 35 nsew signal input
rlabel metal2 s 115938 0 115994 800 6 hk_dat_i[14]
port 36 nsew signal input
rlabel metal2 s 119250 0 119306 800 6 hk_dat_i[15]
port 37 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 hk_dat_i[16]
port 38 nsew signal input
rlabel metal2 s 125966 0 126022 800 6 hk_dat_i[17]
port 39 nsew signal input
rlabel metal2 s 129370 0 129426 800 6 hk_dat_i[18]
port 40 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 hk_dat_i[19]
port 41 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 hk_dat_i[1]
port 42 nsew signal input
rlabel metal2 s 136086 0 136142 800 6 hk_dat_i[20]
port 43 nsew signal input
rlabel metal2 s 139490 0 139546 800 6 hk_dat_i[21]
port 44 nsew signal input
rlabel metal2 s 142802 0 142858 800 6 hk_dat_i[22]
port 45 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 hk_dat_i[23]
port 46 nsew signal input
rlabel metal2 s 149518 0 149574 800 6 hk_dat_i[24]
port 47 nsew signal input
rlabel metal2 s 152922 0 152978 800 6 hk_dat_i[25]
port 48 nsew signal input
rlabel metal2 s 156234 0 156290 800 6 hk_dat_i[26]
port 49 nsew signal input
rlabel metal2 s 159638 0 159694 800 6 hk_dat_i[27]
port 50 nsew signal input
rlabel metal2 s 162950 0 163006 800 6 hk_dat_i[28]
port 51 nsew signal input
rlabel metal2 s 166354 0 166410 800 6 hk_dat_i[29]
port 52 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 hk_dat_i[2]
port 53 nsew signal input
rlabel metal2 s 169666 0 169722 800 6 hk_dat_i[30]
port 54 nsew signal input
rlabel metal2 s 173070 0 173126 800 6 hk_dat_i[31]
port 55 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 hk_dat_i[3]
port 56 nsew signal input
rlabel metal2 s 82266 0 82322 800 6 hk_dat_i[4]
port 57 nsew signal input
rlabel metal2 s 85670 0 85726 800 6 hk_dat_i[5]
port 58 nsew signal input
rlabel metal2 s 88982 0 89038 800 6 hk_dat_i[6]
port 59 nsew signal input
rlabel metal2 s 92386 0 92442 800 6 hk_dat_i[7]
port 60 nsew signal input
rlabel metal2 s 95790 0 95846 800 6 hk_dat_i[8]
port 61 nsew signal input
rlabel metal2 s 99102 0 99158 800 6 hk_dat_i[9]
port 62 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 hk_stb_o
port 63 nsew signal output
rlabel metal2 s 1582 147200 1638 148000 6 la_iena[0]
port 64 nsew signal output
rlabel metal2 s 261758 147200 261814 148000 6 la_iena[100]
port 65 nsew signal output
rlabel metal2 s 264334 147200 264390 148000 6 la_iena[101]
port 66 nsew signal output
rlabel metal2 s 266910 147200 266966 148000 6 la_iena[102]
port 67 nsew signal output
rlabel metal2 s 269486 147200 269542 148000 6 la_iena[103]
port 68 nsew signal output
rlabel metal2 s 272154 147200 272210 148000 6 la_iena[104]
port 69 nsew signal output
rlabel metal2 s 274730 147200 274786 148000 6 la_iena[105]
port 70 nsew signal output
rlabel metal2 s 277306 147200 277362 148000 6 la_iena[106]
port 71 nsew signal output
rlabel metal2 s 279974 147200 280030 148000 6 la_iena[107]
port 72 nsew signal output
rlabel metal2 s 282550 147200 282606 148000 6 la_iena[108]
port 73 nsew signal output
rlabel metal2 s 285126 147200 285182 148000 6 la_iena[109]
port 74 nsew signal output
rlabel metal2 s 27526 147200 27582 148000 6 la_iena[10]
port 75 nsew signal output
rlabel metal2 s 287702 147200 287758 148000 6 la_iena[110]
port 76 nsew signal output
rlabel metal2 s 290370 147200 290426 148000 6 la_iena[111]
port 77 nsew signal output
rlabel metal2 s 292946 147200 293002 148000 6 la_iena[112]
port 78 nsew signal output
rlabel metal2 s 295522 147200 295578 148000 6 la_iena[113]
port 79 nsew signal output
rlabel metal2 s 298190 147200 298246 148000 6 la_iena[114]
port 80 nsew signal output
rlabel metal2 s 300766 147200 300822 148000 6 la_iena[115]
port 81 nsew signal output
rlabel metal2 s 303342 147200 303398 148000 6 la_iena[116]
port 82 nsew signal output
rlabel metal2 s 305918 147200 305974 148000 6 la_iena[117]
port 83 nsew signal output
rlabel metal2 s 308586 147200 308642 148000 6 la_iena[118]
port 84 nsew signal output
rlabel metal2 s 311162 147200 311218 148000 6 la_iena[119]
port 85 nsew signal output
rlabel metal2 s 30194 147200 30250 148000 6 la_iena[11]
port 86 nsew signal output
rlabel metal2 s 313738 147200 313794 148000 6 la_iena[120]
port 87 nsew signal output
rlabel metal2 s 316314 147200 316370 148000 6 la_iena[121]
port 88 nsew signal output
rlabel metal2 s 318982 147200 319038 148000 6 la_iena[122]
port 89 nsew signal output
rlabel metal2 s 321558 147200 321614 148000 6 la_iena[123]
port 90 nsew signal output
rlabel metal2 s 324134 147200 324190 148000 6 la_iena[124]
port 91 nsew signal output
rlabel metal2 s 326802 147200 326858 148000 6 la_iena[125]
port 92 nsew signal output
rlabel metal2 s 329378 147200 329434 148000 6 la_iena[126]
port 93 nsew signal output
rlabel metal2 s 331954 147200 332010 148000 6 la_iena[127]
port 94 nsew signal output
rlabel metal2 s 32770 147200 32826 148000 6 la_iena[12]
port 95 nsew signal output
rlabel metal2 s 35346 147200 35402 148000 6 la_iena[13]
port 96 nsew signal output
rlabel metal2 s 38014 147200 38070 148000 6 la_iena[14]
port 97 nsew signal output
rlabel metal2 s 40590 147200 40646 148000 6 la_iena[15]
port 98 nsew signal output
rlabel metal2 s 43166 147200 43222 148000 6 la_iena[16]
port 99 nsew signal output
rlabel metal2 s 45742 147200 45798 148000 6 la_iena[17]
port 100 nsew signal output
rlabel metal2 s 48410 147200 48466 148000 6 la_iena[18]
port 101 nsew signal output
rlabel metal2 s 50986 147200 51042 148000 6 la_iena[19]
port 102 nsew signal output
rlabel metal2 s 4158 147200 4214 148000 6 la_iena[1]
port 103 nsew signal output
rlabel metal2 s 53562 147200 53618 148000 6 la_iena[20]
port 104 nsew signal output
rlabel metal2 s 56230 147200 56286 148000 6 la_iena[21]
port 105 nsew signal output
rlabel metal2 s 58806 147200 58862 148000 6 la_iena[22]
port 106 nsew signal output
rlabel metal2 s 61382 147200 61438 148000 6 la_iena[23]
port 107 nsew signal output
rlabel metal2 s 63958 147200 64014 148000 6 la_iena[24]
port 108 nsew signal output
rlabel metal2 s 66626 147200 66682 148000 6 la_iena[25]
port 109 nsew signal output
rlabel metal2 s 69202 147200 69258 148000 6 la_iena[26]
port 110 nsew signal output
rlabel metal2 s 71778 147200 71834 148000 6 la_iena[27]
port 111 nsew signal output
rlabel metal2 s 74354 147200 74410 148000 6 la_iena[28]
port 112 nsew signal output
rlabel metal2 s 77022 147200 77078 148000 6 la_iena[29]
port 113 nsew signal output
rlabel metal2 s 6734 147200 6790 148000 6 la_iena[2]
port 114 nsew signal output
rlabel metal2 s 79598 147200 79654 148000 6 la_iena[30]
port 115 nsew signal output
rlabel metal2 s 82174 147200 82230 148000 6 la_iena[31]
port 116 nsew signal output
rlabel metal2 s 84842 147200 84898 148000 6 la_iena[32]
port 117 nsew signal output
rlabel metal2 s 87418 147200 87474 148000 6 la_iena[33]
port 118 nsew signal output
rlabel metal2 s 89994 147200 90050 148000 6 la_iena[34]
port 119 nsew signal output
rlabel metal2 s 92570 147200 92626 148000 6 la_iena[35]
port 120 nsew signal output
rlabel metal2 s 95238 147200 95294 148000 6 la_iena[36]
port 121 nsew signal output
rlabel metal2 s 97814 147200 97870 148000 6 la_iena[37]
port 122 nsew signal output
rlabel metal2 s 100390 147200 100446 148000 6 la_iena[38]
port 123 nsew signal output
rlabel metal2 s 103058 147200 103114 148000 6 la_iena[39]
port 124 nsew signal output
rlabel metal2 s 9310 147200 9366 148000 6 la_iena[3]
port 125 nsew signal output
rlabel metal2 s 105634 147200 105690 148000 6 la_iena[40]
port 126 nsew signal output
rlabel metal2 s 108210 147200 108266 148000 6 la_iena[41]
port 127 nsew signal output
rlabel metal2 s 110786 147200 110842 148000 6 la_iena[42]
port 128 nsew signal output
rlabel metal2 s 113454 147200 113510 148000 6 la_iena[43]
port 129 nsew signal output
rlabel metal2 s 116030 147200 116086 148000 6 la_iena[44]
port 130 nsew signal output
rlabel metal2 s 118606 147200 118662 148000 6 la_iena[45]
port 131 nsew signal output
rlabel metal2 s 121274 147200 121330 148000 6 la_iena[46]
port 132 nsew signal output
rlabel metal2 s 123850 147200 123906 148000 6 la_iena[47]
port 133 nsew signal output
rlabel metal2 s 126426 147200 126482 148000 6 la_iena[48]
port 134 nsew signal output
rlabel metal2 s 129002 147200 129058 148000 6 la_iena[49]
port 135 nsew signal output
rlabel metal2 s 11978 147200 12034 148000 6 la_iena[4]
port 136 nsew signal output
rlabel metal2 s 131670 147200 131726 148000 6 la_iena[50]
port 137 nsew signal output
rlabel metal2 s 134246 147200 134302 148000 6 la_iena[51]
port 138 nsew signal output
rlabel metal2 s 136822 147200 136878 148000 6 la_iena[52]
port 139 nsew signal output
rlabel metal2 s 139398 147200 139454 148000 6 la_iena[53]
port 140 nsew signal output
rlabel metal2 s 142066 147200 142122 148000 6 la_iena[54]
port 141 nsew signal output
rlabel metal2 s 144642 147200 144698 148000 6 la_iena[55]
port 142 nsew signal output
rlabel metal2 s 147218 147200 147274 148000 6 la_iena[56]
port 143 nsew signal output
rlabel metal2 s 149886 147200 149942 148000 6 la_iena[57]
port 144 nsew signal output
rlabel metal2 s 152462 147200 152518 148000 6 la_iena[58]
port 145 nsew signal output
rlabel metal2 s 155038 147200 155094 148000 6 la_iena[59]
port 146 nsew signal output
rlabel metal2 s 14554 147200 14610 148000 6 la_iena[5]
port 147 nsew signal output
rlabel metal2 s 157614 147200 157670 148000 6 la_iena[60]
port 148 nsew signal output
rlabel metal2 s 160282 147200 160338 148000 6 la_iena[61]
port 149 nsew signal output
rlabel metal2 s 162858 147200 162914 148000 6 la_iena[62]
port 150 nsew signal output
rlabel metal2 s 165434 147200 165490 148000 6 la_iena[63]
port 151 nsew signal output
rlabel metal2 s 168102 147200 168158 148000 6 la_iena[64]
port 152 nsew signal output
rlabel metal2 s 170678 147200 170734 148000 6 la_iena[65]
port 153 nsew signal output
rlabel metal2 s 173254 147200 173310 148000 6 la_iena[66]
port 154 nsew signal output
rlabel metal2 s 175830 147200 175886 148000 6 la_iena[67]
port 155 nsew signal output
rlabel metal2 s 178498 147200 178554 148000 6 la_iena[68]
port 156 nsew signal output
rlabel metal2 s 181074 147200 181130 148000 6 la_iena[69]
port 157 nsew signal output
rlabel metal2 s 17130 147200 17186 148000 6 la_iena[6]
port 158 nsew signal output
rlabel metal2 s 183650 147200 183706 148000 6 la_iena[70]
port 159 nsew signal output
rlabel metal2 s 186226 147200 186282 148000 6 la_iena[71]
port 160 nsew signal output
rlabel metal2 s 188894 147200 188950 148000 6 la_iena[72]
port 161 nsew signal output
rlabel metal2 s 191470 147200 191526 148000 6 la_iena[73]
port 162 nsew signal output
rlabel metal2 s 194046 147200 194102 148000 6 la_iena[74]
port 163 nsew signal output
rlabel metal2 s 196714 147200 196770 148000 6 la_iena[75]
port 164 nsew signal output
rlabel metal2 s 199290 147200 199346 148000 6 la_iena[76]
port 165 nsew signal output
rlabel metal2 s 201866 147200 201922 148000 6 la_iena[77]
port 166 nsew signal output
rlabel metal2 s 204442 147200 204498 148000 6 la_iena[78]
port 167 nsew signal output
rlabel metal2 s 207110 147200 207166 148000 6 la_iena[79]
port 168 nsew signal output
rlabel metal2 s 19798 147200 19854 148000 6 la_iena[7]
port 169 nsew signal output
rlabel metal2 s 209686 147200 209742 148000 6 la_iena[80]
port 170 nsew signal output
rlabel metal2 s 212262 147200 212318 148000 6 la_iena[81]
port 171 nsew signal output
rlabel metal2 s 214930 147200 214986 148000 6 la_iena[82]
port 172 nsew signal output
rlabel metal2 s 217506 147200 217562 148000 6 la_iena[83]
port 173 nsew signal output
rlabel metal2 s 220082 147200 220138 148000 6 la_iena[84]
port 174 nsew signal output
rlabel metal2 s 222658 147200 222714 148000 6 la_iena[85]
port 175 nsew signal output
rlabel metal2 s 225326 147200 225382 148000 6 la_iena[86]
port 176 nsew signal output
rlabel metal2 s 227902 147200 227958 148000 6 la_iena[87]
port 177 nsew signal output
rlabel metal2 s 230478 147200 230534 148000 6 la_iena[88]
port 178 nsew signal output
rlabel metal2 s 233146 147200 233202 148000 6 la_iena[89]
port 179 nsew signal output
rlabel metal2 s 22374 147200 22430 148000 6 la_iena[8]
port 180 nsew signal output
rlabel metal2 s 235722 147200 235778 148000 6 la_iena[90]
port 181 nsew signal output
rlabel metal2 s 238298 147200 238354 148000 6 la_iena[91]
port 182 nsew signal output
rlabel metal2 s 240874 147200 240930 148000 6 la_iena[92]
port 183 nsew signal output
rlabel metal2 s 243542 147200 243598 148000 6 la_iena[93]
port 184 nsew signal output
rlabel metal2 s 246118 147200 246174 148000 6 la_iena[94]
port 185 nsew signal output
rlabel metal2 s 248694 147200 248750 148000 6 la_iena[95]
port 186 nsew signal output
rlabel metal2 s 251270 147200 251326 148000 6 la_iena[96]
port 187 nsew signal output
rlabel metal2 s 253938 147200 253994 148000 6 la_iena[97]
port 188 nsew signal output
rlabel metal2 s 256514 147200 256570 148000 6 la_iena[98]
port 189 nsew signal output
rlabel metal2 s 259090 147200 259146 148000 6 la_iena[99]
port 190 nsew signal output
rlabel metal2 s 24950 147200 25006 148000 6 la_iena[9]
port 191 nsew signal output
rlabel metal2 s 2226 147200 2282 148000 6 la_input[0]
port 192 nsew signal input
rlabel metal2 s 262402 147200 262458 148000 6 la_input[100]
port 193 nsew signal input
rlabel metal2 s 264978 147200 265034 148000 6 la_input[101]
port 194 nsew signal input
rlabel metal2 s 267554 147200 267610 148000 6 la_input[102]
port 195 nsew signal input
rlabel metal2 s 270222 147200 270278 148000 6 la_input[103]
port 196 nsew signal input
rlabel metal2 s 272798 147200 272854 148000 6 la_input[104]
port 197 nsew signal input
rlabel metal2 s 275374 147200 275430 148000 6 la_input[105]
port 198 nsew signal input
rlabel metal2 s 277950 147200 278006 148000 6 la_input[106]
port 199 nsew signal input
rlabel metal2 s 280618 147200 280674 148000 6 la_input[107]
port 200 nsew signal input
rlabel metal2 s 283194 147200 283250 148000 6 la_input[108]
port 201 nsew signal input
rlabel metal2 s 285770 147200 285826 148000 6 la_input[109]
port 202 nsew signal input
rlabel metal2 s 28262 147200 28318 148000 6 la_input[10]
port 203 nsew signal input
rlabel metal2 s 288346 147200 288402 148000 6 la_input[110]
port 204 nsew signal input
rlabel metal2 s 291014 147200 291070 148000 6 la_input[111]
port 205 nsew signal input
rlabel metal2 s 293590 147200 293646 148000 6 la_input[112]
port 206 nsew signal input
rlabel metal2 s 296166 147200 296222 148000 6 la_input[113]
port 207 nsew signal input
rlabel metal2 s 298834 147200 298890 148000 6 la_input[114]
port 208 nsew signal input
rlabel metal2 s 301410 147200 301466 148000 6 la_input[115]
port 209 nsew signal input
rlabel metal2 s 303986 147200 304042 148000 6 la_input[116]
port 210 nsew signal input
rlabel metal2 s 306562 147200 306618 148000 6 la_input[117]
port 211 nsew signal input
rlabel metal2 s 309230 147200 309286 148000 6 la_input[118]
port 212 nsew signal input
rlabel metal2 s 311806 147200 311862 148000 6 la_input[119]
port 213 nsew signal input
rlabel metal2 s 30838 147200 30894 148000 6 la_input[11]
port 214 nsew signal input
rlabel metal2 s 314382 147200 314438 148000 6 la_input[120]
port 215 nsew signal input
rlabel metal2 s 317050 147200 317106 148000 6 la_input[121]
port 216 nsew signal input
rlabel metal2 s 319626 147200 319682 148000 6 la_input[122]
port 217 nsew signal input
rlabel metal2 s 322202 147200 322258 148000 6 la_input[123]
port 218 nsew signal input
rlabel metal2 s 324778 147200 324834 148000 6 la_input[124]
port 219 nsew signal input
rlabel metal2 s 327446 147200 327502 148000 6 la_input[125]
port 220 nsew signal input
rlabel metal2 s 330022 147200 330078 148000 6 la_input[126]
port 221 nsew signal input
rlabel metal2 s 332598 147200 332654 148000 6 la_input[127]
port 222 nsew signal input
rlabel metal2 s 33414 147200 33470 148000 6 la_input[12]
port 223 nsew signal input
rlabel metal2 s 35990 147200 36046 148000 6 la_input[13]
port 224 nsew signal input
rlabel metal2 s 38658 147200 38714 148000 6 la_input[14]
port 225 nsew signal input
rlabel metal2 s 41234 147200 41290 148000 6 la_input[15]
port 226 nsew signal input
rlabel metal2 s 43810 147200 43866 148000 6 la_input[16]
port 227 nsew signal input
rlabel metal2 s 46386 147200 46442 148000 6 la_input[17]
port 228 nsew signal input
rlabel metal2 s 49054 147200 49110 148000 6 la_input[18]
port 229 nsew signal input
rlabel metal2 s 51630 147200 51686 148000 6 la_input[19]
port 230 nsew signal input
rlabel metal2 s 4802 147200 4858 148000 6 la_input[1]
port 231 nsew signal input
rlabel metal2 s 54206 147200 54262 148000 6 la_input[20]
port 232 nsew signal input
rlabel metal2 s 56874 147200 56930 148000 6 la_input[21]
port 233 nsew signal input
rlabel metal2 s 59450 147200 59506 148000 6 la_input[22]
port 234 nsew signal input
rlabel metal2 s 62026 147200 62082 148000 6 la_input[23]
port 235 nsew signal input
rlabel metal2 s 64602 147200 64658 148000 6 la_input[24]
port 236 nsew signal input
rlabel metal2 s 67270 147200 67326 148000 6 la_input[25]
port 237 nsew signal input
rlabel metal2 s 69846 147200 69902 148000 6 la_input[26]
port 238 nsew signal input
rlabel metal2 s 72422 147200 72478 148000 6 la_input[27]
port 239 nsew signal input
rlabel metal2 s 75090 147200 75146 148000 6 la_input[28]
port 240 nsew signal input
rlabel metal2 s 77666 147200 77722 148000 6 la_input[29]
port 241 nsew signal input
rlabel metal2 s 7378 147200 7434 148000 6 la_input[2]
port 242 nsew signal input
rlabel metal2 s 80242 147200 80298 148000 6 la_input[30]
port 243 nsew signal input
rlabel metal2 s 82818 147200 82874 148000 6 la_input[31]
port 244 nsew signal input
rlabel metal2 s 85486 147200 85542 148000 6 la_input[32]
port 245 nsew signal input
rlabel metal2 s 88062 147200 88118 148000 6 la_input[33]
port 246 nsew signal input
rlabel metal2 s 90638 147200 90694 148000 6 la_input[34]
port 247 nsew signal input
rlabel metal2 s 93214 147200 93270 148000 6 la_input[35]
port 248 nsew signal input
rlabel metal2 s 95882 147200 95938 148000 6 la_input[36]
port 249 nsew signal input
rlabel metal2 s 98458 147200 98514 148000 6 la_input[37]
port 250 nsew signal input
rlabel metal2 s 101034 147200 101090 148000 6 la_input[38]
port 251 nsew signal input
rlabel metal2 s 103702 147200 103758 148000 6 la_input[39]
port 252 nsew signal input
rlabel metal2 s 10046 147200 10102 148000 6 la_input[3]
port 253 nsew signal input
rlabel metal2 s 106278 147200 106334 148000 6 la_input[40]
port 254 nsew signal input
rlabel metal2 s 108854 147200 108910 148000 6 la_input[41]
port 255 nsew signal input
rlabel metal2 s 111430 147200 111486 148000 6 la_input[42]
port 256 nsew signal input
rlabel metal2 s 114098 147200 114154 148000 6 la_input[43]
port 257 nsew signal input
rlabel metal2 s 116674 147200 116730 148000 6 la_input[44]
port 258 nsew signal input
rlabel metal2 s 119250 147200 119306 148000 6 la_input[45]
port 259 nsew signal input
rlabel metal2 s 121918 147200 121974 148000 6 la_input[46]
port 260 nsew signal input
rlabel metal2 s 124494 147200 124550 148000 6 la_input[47]
port 261 nsew signal input
rlabel metal2 s 127070 147200 127126 148000 6 la_input[48]
port 262 nsew signal input
rlabel metal2 s 129646 147200 129702 148000 6 la_input[49]
port 263 nsew signal input
rlabel metal2 s 12622 147200 12678 148000 6 la_input[4]
port 264 nsew signal input
rlabel metal2 s 132314 147200 132370 148000 6 la_input[50]
port 265 nsew signal input
rlabel metal2 s 134890 147200 134946 148000 6 la_input[51]
port 266 nsew signal input
rlabel metal2 s 137466 147200 137522 148000 6 la_input[52]
port 267 nsew signal input
rlabel metal2 s 140134 147200 140190 148000 6 la_input[53]
port 268 nsew signal input
rlabel metal2 s 142710 147200 142766 148000 6 la_input[54]
port 269 nsew signal input
rlabel metal2 s 145286 147200 145342 148000 6 la_input[55]
port 270 nsew signal input
rlabel metal2 s 147862 147200 147918 148000 6 la_input[56]
port 271 nsew signal input
rlabel metal2 s 150530 147200 150586 148000 6 la_input[57]
port 272 nsew signal input
rlabel metal2 s 153106 147200 153162 148000 6 la_input[58]
port 273 nsew signal input
rlabel metal2 s 155682 147200 155738 148000 6 la_input[59]
port 274 nsew signal input
rlabel metal2 s 15198 147200 15254 148000 6 la_input[5]
port 275 nsew signal input
rlabel metal2 s 158258 147200 158314 148000 6 la_input[60]
port 276 nsew signal input
rlabel metal2 s 160926 147200 160982 148000 6 la_input[61]
port 277 nsew signal input
rlabel metal2 s 163502 147200 163558 148000 6 la_input[62]
port 278 nsew signal input
rlabel metal2 s 166078 147200 166134 148000 6 la_input[63]
port 279 nsew signal input
rlabel metal2 s 168746 147200 168802 148000 6 la_input[64]
port 280 nsew signal input
rlabel metal2 s 171322 147200 171378 148000 6 la_input[65]
port 281 nsew signal input
rlabel metal2 s 173898 147200 173954 148000 6 la_input[66]
port 282 nsew signal input
rlabel metal2 s 176474 147200 176530 148000 6 la_input[67]
port 283 nsew signal input
rlabel metal2 s 179142 147200 179198 148000 6 la_input[68]
port 284 nsew signal input
rlabel metal2 s 181718 147200 181774 148000 6 la_input[69]
port 285 nsew signal input
rlabel metal2 s 17774 147200 17830 148000 6 la_input[6]
port 286 nsew signal input
rlabel metal2 s 184294 147200 184350 148000 6 la_input[70]
port 287 nsew signal input
rlabel metal2 s 186962 147200 187018 148000 6 la_input[71]
port 288 nsew signal input
rlabel metal2 s 189538 147200 189594 148000 6 la_input[72]
port 289 nsew signal input
rlabel metal2 s 192114 147200 192170 148000 6 la_input[73]
port 290 nsew signal input
rlabel metal2 s 194690 147200 194746 148000 6 la_input[74]
port 291 nsew signal input
rlabel metal2 s 197358 147200 197414 148000 6 la_input[75]
port 292 nsew signal input
rlabel metal2 s 199934 147200 199990 148000 6 la_input[76]
port 293 nsew signal input
rlabel metal2 s 202510 147200 202566 148000 6 la_input[77]
port 294 nsew signal input
rlabel metal2 s 205178 147200 205234 148000 6 la_input[78]
port 295 nsew signal input
rlabel metal2 s 207754 147200 207810 148000 6 la_input[79]
port 296 nsew signal input
rlabel metal2 s 20442 147200 20498 148000 6 la_input[7]
port 297 nsew signal input
rlabel metal2 s 210330 147200 210386 148000 6 la_input[80]
port 298 nsew signal input
rlabel metal2 s 212906 147200 212962 148000 6 la_input[81]
port 299 nsew signal input
rlabel metal2 s 215574 147200 215630 148000 6 la_input[82]
port 300 nsew signal input
rlabel metal2 s 218150 147200 218206 148000 6 la_input[83]
port 301 nsew signal input
rlabel metal2 s 220726 147200 220782 148000 6 la_input[84]
port 302 nsew signal input
rlabel metal2 s 223302 147200 223358 148000 6 la_input[85]
port 303 nsew signal input
rlabel metal2 s 225970 147200 226026 148000 6 la_input[86]
port 304 nsew signal input
rlabel metal2 s 228546 147200 228602 148000 6 la_input[87]
port 305 nsew signal input
rlabel metal2 s 231122 147200 231178 148000 6 la_input[88]
port 306 nsew signal input
rlabel metal2 s 233790 147200 233846 148000 6 la_input[89]
port 307 nsew signal input
rlabel metal2 s 23018 147200 23074 148000 6 la_input[8]
port 308 nsew signal input
rlabel metal2 s 236366 147200 236422 148000 6 la_input[90]
port 309 nsew signal input
rlabel metal2 s 238942 147200 238998 148000 6 la_input[91]
port 310 nsew signal input
rlabel metal2 s 241518 147200 241574 148000 6 la_input[92]
port 311 nsew signal input
rlabel metal2 s 244186 147200 244242 148000 6 la_input[93]
port 312 nsew signal input
rlabel metal2 s 246762 147200 246818 148000 6 la_input[94]
port 313 nsew signal input
rlabel metal2 s 249338 147200 249394 148000 6 la_input[95]
port 314 nsew signal input
rlabel metal2 s 252006 147200 252062 148000 6 la_input[96]
port 315 nsew signal input
rlabel metal2 s 254582 147200 254638 148000 6 la_input[97]
port 316 nsew signal input
rlabel metal2 s 257158 147200 257214 148000 6 la_input[98]
port 317 nsew signal input
rlabel metal2 s 259734 147200 259790 148000 6 la_input[99]
port 318 nsew signal input
rlabel metal2 s 25594 147200 25650 148000 6 la_input[9]
port 319 nsew signal input
rlabel metal2 s 2870 147200 2926 148000 6 la_oenb[0]
port 320 nsew signal output
rlabel metal2 s 263046 147200 263102 148000 6 la_oenb[100]
port 321 nsew signal output
rlabel metal2 s 265622 147200 265678 148000 6 la_oenb[101]
port 322 nsew signal output
rlabel metal2 s 268198 147200 268254 148000 6 la_oenb[102]
port 323 nsew signal output
rlabel metal2 s 270866 147200 270922 148000 6 la_oenb[103]
port 324 nsew signal output
rlabel metal2 s 273442 147200 273498 148000 6 la_oenb[104]
port 325 nsew signal output
rlabel metal2 s 276018 147200 276074 148000 6 la_oenb[105]
port 326 nsew signal output
rlabel metal2 s 278594 147200 278650 148000 6 la_oenb[106]
port 327 nsew signal output
rlabel metal2 s 281262 147200 281318 148000 6 la_oenb[107]
port 328 nsew signal output
rlabel metal2 s 283838 147200 283894 148000 6 la_oenb[108]
port 329 nsew signal output
rlabel metal2 s 286414 147200 286470 148000 6 la_oenb[109]
port 330 nsew signal output
rlabel metal2 s 28906 147200 28962 148000 6 la_oenb[10]
port 331 nsew signal output
rlabel metal2 s 289082 147200 289138 148000 6 la_oenb[110]
port 332 nsew signal output
rlabel metal2 s 291658 147200 291714 148000 6 la_oenb[111]
port 333 nsew signal output
rlabel metal2 s 294234 147200 294290 148000 6 la_oenb[112]
port 334 nsew signal output
rlabel metal2 s 296810 147200 296866 148000 6 la_oenb[113]
port 335 nsew signal output
rlabel metal2 s 299478 147200 299534 148000 6 la_oenb[114]
port 336 nsew signal output
rlabel metal2 s 302054 147200 302110 148000 6 la_oenb[115]
port 337 nsew signal output
rlabel metal2 s 304630 147200 304686 148000 6 la_oenb[116]
port 338 nsew signal output
rlabel metal2 s 307298 147200 307354 148000 6 la_oenb[117]
port 339 nsew signal output
rlabel metal2 s 309874 147200 309930 148000 6 la_oenb[118]
port 340 nsew signal output
rlabel metal2 s 312450 147200 312506 148000 6 la_oenb[119]
port 341 nsew signal output
rlabel metal2 s 31482 147200 31538 148000 6 la_oenb[11]
port 342 nsew signal output
rlabel metal2 s 315026 147200 315082 148000 6 la_oenb[120]
port 343 nsew signal output
rlabel metal2 s 317694 147200 317750 148000 6 la_oenb[121]
port 344 nsew signal output
rlabel metal2 s 320270 147200 320326 148000 6 la_oenb[122]
port 345 nsew signal output
rlabel metal2 s 322846 147200 322902 148000 6 la_oenb[123]
port 346 nsew signal output
rlabel metal2 s 325422 147200 325478 148000 6 la_oenb[124]
port 347 nsew signal output
rlabel metal2 s 328090 147200 328146 148000 6 la_oenb[125]
port 348 nsew signal output
rlabel metal2 s 330666 147200 330722 148000 6 la_oenb[126]
port 349 nsew signal output
rlabel metal2 s 333242 147200 333298 148000 6 la_oenb[127]
port 350 nsew signal output
rlabel metal2 s 34058 147200 34114 148000 6 la_oenb[12]
port 351 nsew signal output
rlabel metal2 s 36634 147200 36690 148000 6 la_oenb[13]
port 352 nsew signal output
rlabel metal2 s 39302 147200 39358 148000 6 la_oenb[14]
port 353 nsew signal output
rlabel metal2 s 41878 147200 41934 148000 6 la_oenb[15]
port 354 nsew signal output
rlabel metal2 s 44454 147200 44510 148000 6 la_oenb[16]
port 355 nsew signal output
rlabel metal2 s 47122 147200 47178 148000 6 la_oenb[17]
port 356 nsew signal output
rlabel metal2 s 49698 147200 49754 148000 6 la_oenb[18]
port 357 nsew signal output
rlabel metal2 s 52274 147200 52330 148000 6 la_oenb[19]
port 358 nsew signal output
rlabel metal2 s 5446 147200 5502 148000 6 la_oenb[1]
port 359 nsew signal output
rlabel metal2 s 54850 147200 54906 148000 6 la_oenb[20]
port 360 nsew signal output
rlabel metal2 s 57518 147200 57574 148000 6 la_oenb[21]
port 361 nsew signal output
rlabel metal2 s 60094 147200 60150 148000 6 la_oenb[22]
port 362 nsew signal output
rlabel metal2 s 62670 147200 62726 148000 6 la_oenb[23]
port 363 nsew signal output
rlabel metal2 s 65246 147200 65302 148000 6 la_oenb[24]
port 364 nsew signal output
rlabel metal2 s 67914 147200 67970 148000 6 la_oenb[25]
port 365 nsew signal output
rlabel metal2 s 70490 147200 70546 148000 6 la_oenb[26]
port 366 nsew signal output
rlabel metal2 s 73066 147200 73122 148000 6 la_oenb[27]
port 367 nsew signal output
rlabel metal2 s 75734 147200 75790 148000 6 la_oenb[28]
port 368 nsew signal output
rlabel metal2 s 78310 147200 78366 148000 6 la_oenb[29]
port 369 nsew signal output
rlabel metal2 s 8022 147200 8078 148000 6 la_oenb[2]
port 370 nsew signal output
rlabel metal2 s 80886 147200 80942 148000 6 la_oenb[30]
port 371 nsew signal output
rlabel metal2 s 83462 147200 83518 148000 6 la_oenb[31]
port 372 nsew signal output
rlabel metal2 s 86130 147200 86186 148000 6 la_oenb[32]
port 373 nsew signal output
rlabel metal2 s 88706 147200 88762 148000 6 la_oenb[33]
port 374 nsew signal output
rlabel metal2 s 91282 147200 91338 148000 6 la_oenb[34]
port 375 nsew signal output
rlabel metal2 s 93950 147200 94006 148000 6 la_oenb[35]
port 376 nsew signal output
rlabel metal2 s 96526 147200 96582 148000 6 la_oenb[36]
port 377 nsew signal output
rlabel metal2 s 99102 147200 99158 148000 6 la_oenb[37]
port 378 nsew signal output
rlabel metal2 s 101678 147200 101734 148000 6 la_oenb[38]
port 379 nsew signal output
rlabel metal2 s 104346 147200 104402 148000 6 la_oenb[39]
port 380 nsew signal output
rlabel metal2 s 10690 147200 10746 148000 6 la_oenb[3]
port 381 nsew signal output
rlabel metal2 s 106922 147200 106978 148000 6 la_oenb[40]
port 382 nsew signal output
rlabel metal2 s 109498 147200 109554 148000 6 la_oenb[41]
port 383 nsew signal output
rlabel metal2 s 112166 147200 112222 148000 6 la_oenb[42]
port 384 nsew signal output
rlabel metal2 s 114742 147200 114798 148000 6 la_oenb[43]
port 385 nsew signal output
rlabel metal2 s 117318 147200 117374 148000 6 la_oenb[44]
port 386 nsew signal output
rlabel metal2 s 119894 147200 119950 148000 6 la_oenb[45]
port 387 nsew signal output
rlabel metal2 s 122562 147200 122618 148000 6 la_oenb[46]
port 388 nsew signal output
rlabel metal2 s 125138 147200 125194 148000 6 la_oenb[47]
port 389 nsew signal output
rlabel metal2 s 127714 147200 127770 148000 6 la_oenb[48]
port 390 nsew signal output
rlabel metal2 s 130290 147200 130346 148000 6 la_oenb[49]
port 391 nsew signal output
rlabel metal2 s 13266 147200 13322 148000 6 la_oenb[4]
port 392 nsew signal output
rlabel metal2 s 132958 147200 133014 148000 6 la_oenb[50]
port 393 nsew signal output
rlabel metal2 s 135534 147200 135590 148000 6 la_oenb[51]
port 394 nsew signal output
rlabel metal2 s 138110 147200 138166 148000 6 la_oenb[52]
port 395 nsew signal output
rlabel metal2 s 140778 147200 140834 148000 6 la_oenb[53]
port 396 nsew signal output
rlabel metal2 s 143354 147200 143410 148000 6 la_oenb[54]
port 397 nsew signal output
rlabel metal2 s 145930 147200 145986 148000 6 la_oenb[55]
port 398 nsew signal output
rlabel metal2 s 148506 147200 148562 148000 6 la_oenb[56]
port 399 nsew signal output
rlabel metal2 s 151174 147200 151230 148000 6 la_oenb[57]
port 400 nsew signal output
rlabel metal2 s 153750 147200 153806 148000 6 la_oenb[58]
port 401 nsew signal output
rlabel metal2 s 156326 147200 156382 148000 6 la_oenb[59]
port 402 nsew signal output
rlabel metal2 s 15842 147200 15898 148000 6 la_oenb[5]
port 403 nsew signal output
rlabel metal2 s 158994 147200 159050 148000 6 la_oenb[60]
port 404 nsew signal output
rlabel metal2 s 161570 147200 161626 148000 6 la_oenb[61]
port 405 nsew signal output
rlabel metal2 s 164146 147200 164202 148000 6 la_oenb[62]
port 406 nsew signal output
rlabel metal2 s 166722 147200 166778 148000 6 la_oenb[63]
port 407 nsew signal output
rlabel metal2 s 169390 147200 169446 148000 6 la_oenb[64]
port 408 nsew signal output
rlabel metal2 s 171966 147200 172022 148000 6 la_oenb[65]
port 409 nsew signal output
rlabel metal2 s 174542 147200 174598 148000 6 la_oenb[66]
port 410 nsew signal output
rlabel metal2 s 177210 147200 177266 148000 6 la_oenb[67]
port 411 nsew signal output
rlabel metal2 s 179786 147200 179842 148000 6 la_oenb[68]
port 412 nsew signal output
rlabel metal2 s 182362 147200 182418 148000 6 la_oenb[69]
port 413 nsew signal output
rlabel metal2 s 18418 147200 18474 148000 6 la_oenb[6]
port 414 nsew signal output
rlabel metal2 s 184938 147200 184994 148000 6 la_oenb[70]
port 415 nsew signal output
rlabel metal2 s 187606 147200 187662 148000 6 la_oenb[71]
port 416 nsew signal output
rlabel metal2 s 190182 147200 190238 148000 6 la_oenb[72]
port 417 nsew signal output
rlabel metal2 s 192758 147200 192814 148000 6 la_oenb[73]
port 418 nsew signal output
rlabel metal2 s 195334 147200 195390 148000 6 la_oenb[74]
port 419 nsew signal output
rlabel metal2 s 198002 147200 198058 148000 6 la_oenb[75]
port 420 nsew signal output
rlabel metal2 s 200578 147200 200634 148000 6 la_oenb[76]
port 421 nsew signal output
rlabel metal2 s 203154 147200 203210 148000 6 la_oenb[77]
port 422 nsew signal output
rlabel metal2 s 205822 147200 205878 148000 6 la_oenb[78]
port 423 nsew signal output
rlabel metal2 s 208398 147200 208454 148000 6 la_oenb[79]
port 424 nsew signal output
rlabel metal2 s 21086 147200 21142 148000 6 la_oenb[7]
port 425 nsew signal output
rlabel metal2 s 210974 147200 211030 148000 6 la_oenb[80]
port 426 nsew signal output
rlabel metal2 s 213550 147200 213606 148000 6 la_oenb[81]
port 427 nsew signal output
rlabel metal2 s 216218 147200 216274 148000 6 la_oenb[82]
port 428 nsew signal output
rlabel metal2 s 218794 147200 218850 148000 6 la_oenb[83]
port 429 nsew signal output
rlabel metal2 s 221370 147200 221426 148000 6 la_oenb[84]
port 430 nsew signal output
rlabel metal2 s 224038 147200 224094 148000 6 la_oenb[85]
port 431 nsew signal output
rlabel metal2 s 226614 147200 226670 148000 6 la_oenb[86]
port 432 nsew signal output
rlabel metal2 s 229190 147200 229246 148000 6 la_oenb[87]
port 433 nsew signal output
rlabel metal2 s 231766 147200 231822 148000 6 la_oenb[88]
port 434 nsew signal output
rlabel metal2 s 234434 147200 234490 148000 6 la_oenb[89]
port 435 nsew signal output
rlabel metal2 s 23662 147200 23718 148000 6 la_oenb[8]
port 436 nsew signal output
rlabel metal2 s 237010 147200 237066 148000 6 la_oenb[90]
port 437 nsew signal output
rlabel metal2 s 239586 147200 239642 148000 6 la_oenb[91]
port 438 nsew signal output
rlabel metal2 s 242254 147200 242310 148000 6 la_oenb[92]
port 439 nsew signal output
rlabel metal2 s 244830 147200 244886 148000 6 la_oenb[93]
port 440 nsew signal output
rlabel metal2 s 247406 147200 247462 148000 6 la_oenb[94]
port 441 nsew signal output
rlabel metal2 s 249982 147200 250038 148000 6 la_oenb[95]
port 442 nsew signal output
rlabel metal2 s 252650 147200 252706 148000 6 la_oenb[96]
port 443 nsew signal output
rlabel metal2 s 255226 147200 255282 148000 6 la_oenb[97]
port 444 nsew signal output
rlabel metal2 s 257802 147200 257858 148000 6 la_oenb[98]
port 445 nsew signal output
rlabel metal2 s 260378 147200 260434 148000 6 la_oenb[99]
port 446 nsew signal output
rlabel metal2 s 26238 147200 26294 148000 6 la_oenb[9]
port 447 nsew signal output
rlabel metal2 s 3514 147200 3570 148000 6 la_output[0]
port 448 nsew signal output
rlabel metal2 s 263690 147200 263746 148000 6 la_output[100]
port 449 nsew signal output
rlabel metal2 s 266266 147200 266322 148000 6 la_output[101]
port 450 nsew signal output
rlabel metal2 s 268842 147200 268898 148000 6 la_output[102]
port 451 nsew signal output
rlabel metal2 s 271510 147200 271566 148000 6 la_output[103]
port 452 nsew signal output
rlabel metal2 s 274086 147200 274142 148000 6 la_output[104]
port 453 nsew signal output
rlabel metal2 s 276662 147200 276718 148000 6 la_output[105]
port 454 nsew signal output
rlabel metal2 s 279238 147200 279294 148000 6 la_output[106]
port 455 nsew signal output
rlabel metal2 s 281906 147200 281962 148000 6 la_output[107]
port 456 nsew signal output
rlabel metal2 s 284482 147200 284538 148000 6 la_output[108]
port 457 nsew signal output
rlabel metal2 s 287058 147200 287114 148000 6 la_output[109]
port 458 nsew signal output
rlabel metal2 s 29550 147200 29606 148000 6 la_output[10]
port 459 nsew signal output
rlabel metal2 s 289726 147200 289782 148000 6 la_output[110]
port 460 nsew signal output
rlabel metal2 s 292302 147200 292358 148000 6 la_output[111]
port 461 nsew signal output
rlabel metal2 s 294878 147200 294934 148000 6 la_output[112]
port 462 nsew signal output
rlabel metal2 s 297454 147200 297510 148000 6 la_output[113]
port 463 nsew signal output
rlabel metal2 s 300122 147200 300178 148000 6 la_output[114]
port 464 nsew signal output
rlabel metal2 s 302698 147200 302754 148000 6 la_output[115]
port 465 nsew signal output
rlabel metal2 s 305274 147200 305330 148000 6 la_output[116]
port 466 nsew signal output
rlabel metal2 s 307942 147200 307998 148000 6 la_output[117]
port 467 nsew signal output
rlabel metal2 s 310518 147200 310574 148000 6 la_output[118]
port 468 nsew signal output
rlabel metal2 s 313094 147200 313150 148000 6 la_output[119]
port 469 nsew signal output
rlabel metal2 s 32126 147200 32182 148000 6 la_output[11]
port 470 nsew signal output
rlabel metal2 s 315670 147200 315726 148000 6 la_output[120]
port 471 nsew signal output
rlabel metal2 s 318338 147200 318394 148000 6 la_output[121]
port 472 nsew signal output
rlabel metal2 s 320914 147200 320970 148000 6 la_output[122]
port 473 nsew signal output
rlabel metal2 s 323490 147200 323546 148000 6 la_output[123]
port 474 nsew signal output
rlabel metal2 s 326158 147200 326214 148000 6 la_output[124]
port 475 nsew signal output
rlabel metal2 s 328734 147200 328790 148000 6 la_output[125]
port 476 nsew signal output
rlabel metal2 s 331310 147200 331366 148000 6 la_output[126]
port 477 nsew signal output
rlabel metal2 s 333886 147200 333942 148000 6 la_output[127]
port 478 nsew signal output
rlabel metal2 s 34702 147200 34758 148000 6 la_output[12]
port 479 nsew signal output
rlabel metal2 s 37278 147200 37334 148000 6 la_output[13]
port 480 nsew signal output
rlabel metal2 s 39946 147200 40002 148000 6 la_output[14]
port 481 nsew signal output
rlabel metal2 s 42522 147200 42578 148000 6 la_output[15]
port 482 nsew signal output
rlabel metal2 s 45098 147200 45154 148000 6 la_output[16]
port 483 nsew signal output
rlabel metal2 s 47766 147200 47822 148000 6 la_output[17]
port 484 nsew signal output
rlabel metal2 s 50342 147200 50398 148000 6 la_output[18]
port 485 nsew signal output
rlabel metal2 s 52918 147200 52974 148000 6 la_output[19]
port 486 nsew signal output
rlabel metal2 s 6090 147200 6146 148000 6 la_output[1]
port 487 nsew signal output
rlabel metal2 s 55494 147200 55550 148000 6 la_output[20]
port 488 nsew signal output
rlabel metal2 s 58162 147200 58218 148000 6 la_output[21]
port 489 nsew signal output
rlabel metal2 s 60738 147200 60794 148000 6 la_output[22]
port 490 nsew signal output
rlabel metal2 s 63314 147200 63370 148000 6 la_output[23]
port 491 nsew signal output
rlabel metal2 s 65982 147200 66038 148000 6 la_output[24]
port 492 nsew signal output
rlabel metal2 s 68558 147200 68614 148000 6 la_output[25]
port 493 nsew signal output
rlabel metal2 s 71134 147200 71190 148000 6 la_output[26]
port 494 nsew signal output
rlabel metal2 s 73710 147200 73766 148000 6 la_output[27]
port 495 nsew signal output
rlabel metal2 s 76378 147200 76434 148000 6 la_output[28]
port 496 nsew signal output
rlabel metal2 s 78954 147200 79010 148000 6 la_output[29]
port 497 nsew signal output
rlabel metal2 s 8666 147200 8722 148000 6 la_output[2]
port 498 nsew signal output
rlabel metal2 s 81530 147200 81586 148000 6 la_output[30]
port 499 nsew signal output
rlabel metal2 s 84198 147200 84254 148000 6 la_output[31]
port 500 nsew signal output
rlabel metal2 s 86774 147200 86830 148000 6 la_output[32]
port 501 nsew signal output
rlabel metal2 s 89350 147200 89406 148000 6 la_output[33]
port 502 nsew signal output
rlabel metal2 s 91926 147200 91982 148000 6 la_output[34]
port 503 nsew signal output
rlabel metal2 s 94594 147200 94650 148000 6 la_output[35]
port 504 nsew signal output
rlabel metal2 s 97170 147200 97226 148000 6 la_output[36]
port 505 nsew signal output
rlabel metal2 s 99746 147200 99802 148000 6 la_output[37]
port 506 nsew signal output
rlabel metal2 s 102322 147200 102378 148000 6 la_output[38]
port 507 nsew signal output
rlabel metal2 s 104990 147200 105046 148000 6 la_output[39]
port 508 nsew signal output
rlabel metal2 s 11334 147200 11390 148000 6 la_output[3]
port 509 nsew signal output
rlabel metal2 s 107566 147200 107622 148000 6 la_output[40]
port 510 nsew signal output
rlabel metal2 s 110142 147200 110198 148000 6 la_output[41]
port 511 nsew signal output
rlabel metal2 s 112810 147200 112866 148000 6 la_output[42]
port 512 nsew signal output
rlabel metal2 s 115386 147200 115442 148000 6 la_output[43]
port 513 nsew signal output
rlabel metal2 s 117962 147200 118018 148000 6 la_output[44]
port 514 nsew signal output
rlabel metal2 s 120538 147200 120594 148000 6 la_output[45]
port 515 nsew signal output
rlabel metal2 s 123206 147200 123262 148000 6 la_output[46]
port 516 nsew signal output
rlabel metal2 s 125782 147200 125838 148000 6 la_output[47]
port 517 nsew signal output
rlabel metal2 s 128358 147200 128414 148000 6 la_output[48]
port 518 nsew signal output
rlabel metal2 s 131026 147200 131082 148000 6 la_output[49]
port 519 nsew signal output
rlabel metal2 s 13910 147200 13966 148000 6 la_output[4]
port 520 nsew signal output
rlabel metal2 s 133602 147200 133658 148000 6 la_output[50]
port 521 nsew signal output
rlabel metal2 s 136178 147200 136234 148000 6 la_output[51]
port 522 nsew signal output
rlabel metal2 s 138754 147200 138810 148000 6 la_output[52]
port 523 nsew signal output
rlabel metal2 s 141422 147200 141478 148000 6 la_output[53]
port 524 nsew signal output
rlabel metal2 s 143998 147200 144054 148000 6 la_output[54]
port 525 nsew signal output
rlabel metal2 s 146574 147200 146630 148000 6 la_output[55]
port 526 nsew signal output
rlabel metal2 s 149242 147200 149298 148000 6 la_output[56]
port 527 nsew signal output
rlabel metal2 s 151818 147200 151874 148000 6 la_output[57]
port 528 nsew signal output
rlabel metal2 s 154394 147200 154450 148000 6 la_output[58]
port 529 nsew signal output
rlabel metal2 s 156970 147200 157026 148000 6 la_output[59]
port 530 nsew signal output
rlabel metal2 s 16486 147200 16542 148000 6 la_output[5]
port 531 nsew signal output
rlabel metal2 s 159638 147200 159694 148000 6 la_output[60]
port 532 nsew signal output
rlabel metal2 s 162214 147200 162270 148000 6 la_output[61]
port 533 nsew signal output
rlabel metal2 s 164790 147200 164846 148000 6 la_output[62]
port 534 nsew signal output
rlabel metal2 s 167366 147200 167422 148000 6 la_output[63]
port 535 nsew signal output
rlabel metal2 s 170034 147200 170090 148000 6 la_output[64]
port 536 nsew signal output
rlabel metal2 s 172610 147200 172666 148000 6 la_output[65]
port 537 nsew signal output
rlabel metal2 s 175186 147200 175242 148000 6 la_output[66]
port 538 nsew signal output
rlabel metal2 s 177854 147200 177910 148000 6 la_output[67]
port 539 nsew signal output
rlabel metal2 s 180430 147200 180486 148000 6 la_output[68]
port 540 nsew signal output
rlabel metal2 s 183006 147200 183062 148000 6 la_output[69]
port 541 nsew signal output
rlabel metal2 s 19154 147200 19210 148000 6 la_output[6]
port 542 nsew signal output
rlabel metal2 s 185582 147200 185638 148000 6 la_output[70]
port 543 nsew signal output
rlabel metal2 s 188250 147200 188306 148000 6 la_output[71]
port 544 nsew signal output
rlabel metal2 s 190826 147200 190882 148000 6 la_output[72]
port 545 nsew signal output
rlabel metal2 s 193402 147200 193458 148000 6 la_output[73]
port 546 nsew signal output
rlabel metal2 s 196070 147200 196126 148000 6 la_output[74]
port 547 nsew signal output
rlabel metal2 s 198646 147200 198702 148000 6 la_output[75]
port 548 nsew signal output
rlabel metal2 s 201222 147200 201278 148000 6 la_output[76]
port 549 nsew signal output
rlabel metal2 s 203798 147200 203854 148000 6 la_output[77]
port 550 nsew signal output
rlabel metal2 s 206466 147200 206522 148000 6 la_output[78]
port 551 nsew signal output
rlabel metal2 s 209042 147200 209098 148000 6 la_output[79]
port 552 nsew signal output
rlabel metal2 s 21730 147200 21786 148000 6 la_output[7]
port 553 nsew signal output
rlabel metal2 s 211618 147200 211674 148000 6 la_output[80]
port 554 nsew signal output
rlabel metal2 s 214286 147200 214342 148000 6 la_output[81]
port 555 nsew signal output
rlabel metal2 s 216862 147200 216918 148000 6 la_output[82]
port 556 nsew signal output
rlabel metal2 s 219438 147200 219494 148000 6 la_output[83]
port 557 nsew signal output
rlabel metal2 s 222014 147200 222070 148000 6 la_output[84]
port 558 nsew signal output
rlabel metal2 s 224682 147200 224738 148000 6 la_output[85]
port 559 nsew signal output
rlabel metal2 s 227258 147200 227314 148000 6 la_output[86]
port 560 nsew signal output
rlabel metal2 s 229834 147200 229890 148000 6 la_output[87]
port 561 nsew signal output
rlabel metal2 s 232410 147200 232466 148000 6 la_output[88]
port 562 nsew signal output
rlabel metal2 s 235078 147200 235134 148000 6 la_output[89]
port 563 nsew signal output
rlabel metal2 s 24306 147200 24362 148000 6 la_output[8]
port 564 nsew signal output
rlabel metal2 s 237654 147200 237710 148000 6 la_output[90]
port 565 nsew signal output
rlabel metal2 s 240230 147200 240286 148000 6 la_output[91]
port 566 nsew signal output
rlabel metal2 s 242898 147200 242954 148000 6 la_output[92]
port 567 nsew signal output
rlabel metal2 s 245474 147200 245530 148000 6 la_output[93]
port 568 nsew signal output
rlabel metal2 s 248050 147200 248106 148000 6 la_output[94]
port 569 nsew signal output
rlabel metal2 s 250626 147200 250682 148000 6 la_output[95]
port 570 nsew signal output
rlabel metal2 s 253294 147200 253350 148000 6 la_output[96]
port 571 nsew signal output
rlabel metal2 s 255870 147200 255926 148000 6 la_output[97]
port 572 nsew signal output
rlabel metal2 s 258446 147200 258502 148000 6 la_output[98]
port 573 nsew signal output
rlabel metal2 s 261114 147200 261170 148000 6 la_output[99]
port 574 nsew signal output
rlabel metal2 s 26882 147200 26938 148000 6 la_output[9]
port 575 nsew signal output
rlabel metal2 s 344466 0 344522 800 6 mgmt_soc_dff_A[0]
port 576 nsew signal output
rlabel metal3 s 399200 16600 400000 16720 6 mgmt_soc_dff_A[1]
port 577 nsew signal output
rlabel metal2 s 351182 0 351238 800 6 mgmt_soc_dff_A[2]
port 578 nsew signal output
rlabel metal3 s 0 102960 800 103080 6 mgmt_soc_dff_A[3]
port 579 nsew signal output
rlabel metal3 s 399200 36864 400000 36984 6 mgmt_soc_dff_A[4]
port 580 nsew signal output
rlabel metal2 s 390466 147200 390522 148000 6 mgmt_soc_dff_A[5]
port 581 nsew signal output
rlabel metal3 s 399200 50328 400000 50448 6 mgmt_soc_dff_A[6]
port 582 nsew signal output
rlabel metal3 s 0 112616 800 112736 6 mgmt_soc_dff_A[7]
port 583 nsew signal output
rlabel metal2 s 385958 147200 386014 148000 6 mgmt_soc_dff_Di[0]
port 584 nsew signal output
rlabel metal3 s 399200 70456 400000 70576 6 mgmt_soc_dff_Di[10]
port 585 nsew signal output
rlabel metal3 s 0 115064 800 115184 6 mgmt_soc_dff_Di[11]
port 586 nsew signal output
rlabel metal2 s 394422 147200 394478 148000 6 mgmt_soc_dff_Di[12]
port 587 nsew signal output
rlabel metal3 s 0 119824 800 119944 6 mgmt_soc_dff_Di[13]
port 588 nsew signal output
rlabel metal3 s 399200 83920 400000 84040 6 mgmt_soc_dff_Di[14]
port 589 nsew signal output
rlabel metal3 s 0 122272 800 122392 6 mgmt_soc_dff_Di[15]
port 590 nsew signal output
rlabel metal3 s 0 127168 800 127288 6 mgmt_soc_dff_Di[16]
port 591 nsew signal output
rlabel metal3 s 399200 90584 400000 90704 6 mgmt_soc_dff_Di[17]
port 592 nsew signal output
rlabel metal3 s 399200 97384 400000 97504 6 mgmt_soc_dff_Di[18]
port 593 nsew signal output
rlabel metal2 s 378138 0 378194 800 6 mgmt_soc_dff_Di[19]
port 594 nsew signal output
rlabel metal3 s 399200 23400 400000 23520 6 mgmt_soc_dff_Di[1]
port 595 nsew signal output
rlabel metal2 s 395710 147200 395766 148000 6 mgmt_soc_dff_Di[20]
port 596 nsew signal output
rlabel metal2 s 384854 0 384910 800 6 mgmt_soc_dff_Di[21]
port 597 nsew signal output
rlabel metal3 s 0 134376 800 134496 6 mgmt_soc_dff_Di[22]
port 598 nsew signal output
rlabel metal3 s 0 136824 800 136944 6 mgmt_soc_dff_Di[23]
port 599 nsew signal output
rlabel metal2 s 388166 0 388222 800 6 mgmt_soc_dff_Di[24]
port 600 nsew signal output
rlabel metal2 s 397642 147200 397698 148000 6 mgmt_soc_dff_Di[25]
port 601 nsew signal output
rlabel metal2 s 391570 0 391626 800 6 mgmt_soc_dff_Di[26]
port 602 nsew signal output
rlabel metal2 s 398930 147200 398986 148000 6 mgmt_soc_dff_Di[27]
port 603 nsew signal output
rlabel metal2 s 398286 0 398342 800 6 mgmt_soc_dff_Di[28]
port 604 nsew signal output
rlabel metal3 s 399200 137776 400000 137896 6 mgmt_soc_dff_Di[29]
port 605 nsew signal output
rlabel metal2 s 387246 147200 387302 148000 6 mgmt_soc_dff_Di[2]
port 606 nsew signal output
rlabel metal3 s 0 139272 800 139392 6 mgmt_soc_dff_Di[30]
port 607 nsew signal output
rlabel metal3 s 0 144168 800 144288 6 mgmt_soc_dff_Di[31]
port 608 nsew signal output
rlabel metal2 s 357990 0 358046 800 6 mgmt_soc_dff_Di[3]
port 609 nsew signal output
rlabel metal3 s 399200 43528 400000 43648 6 mgmt_soc_dff_Di[4]
port 610 nsew signal output
rlabel metal3 s 0 107720 800 107840 6 mgmt_soc_dff_Di[5]
port 611 nsew signal output
rlabel metal2 s 368018 0 368074 800 6 mgmt_soc_dff_Di[6]
port 612 nsew signal output
rlabel metal2 s 391846 147200 391902 148000 6 mgmt_soc_dff_Di[7]
port 613 nsew signal output
rlabel metal2 s 393134 147200 393190 148000 6 mgmt_soc_dff_Di[8]
port 614 nsew signal output
rlabel metal3 s 399200 63792 400000 63912 6 mgmt_soc_dff_Di[9]
port 615 nsew signal output
rlabel metal3 s 399200 3272 400000 3392 6 mgmt_soc_dff_Do[0]
port 616 nsew signal input
rlabel metal2 s 393778 147200 393834 148000 6 mgmt_soc_dff_Do[10]
port 617 nsew signal input
rlabel metal3 s 0 117512 800 117632 6 mgmt_soc_dff_Do[11]
port 618 nsew signal input
rlabel metal3 s 399200 77256 400000 77376 6 mgmt_soc_dff_Do[12]
port 619 nsew signal input
rlabel metal2 s 395066 147200 395122 148000 6 mgmt_soc_dff_Do[13]
port 620 nsew signal input
rlabel metal2 s 374734 0 374790 800 6 mgmt_soc_dff_Do[14]
port 621 nsew signal input
rlabel metal3 s 0 124720 800 124840 6 mgmt_soc_dff_Do[15]
port 622 nsew signal input
rlabel metal3 s 0 129616 800 129736 6 mgmt_soc_dff_Do[16]
port 623 nsew signal input
rlabel metal3 s 0 132064 800 132184 6 mgmt_soc_dff_Do[17]
port 624 nsew signal input
rlabel metal3 s 399200 104048 400000 104168 6 mgmt_soc_dff_Do[18]
port 625 nsew signal input
rlabel metal2 s 381450 0 381506 800 6 mgmt_soc_dff_Do[19]
port 626 nsew signal input
rlabel metal2 s 386602 147200 386658 148000 6 mgmt_soc_dff_Do[1]
port 627 nsew signal input
rlabel metal3 s 399200 110848 400000 110968 6 mgmt_soc_dff_Do[20]
port 628 nsew signal input
rlabel metal3 s 399200 117512 400000 117632 6 mgmt_soc_dff_Do[21]
port 629 nsew signal input
rlabel metal2 s 396354 147200 396410 148000 6 mgmt_soc_dff_Do[22]
port 630 nsew signal input
rlabel metal3 s 399200 124312 400000 124432 6 mgmt_soc_dff_Do[23]
port 631 nsew signal input
rlabel metal2 s 396998 147200 397054 148000 6 mgmt_soc_dff_Do[24]
port 632 nsew signal input
rlabel metal2 s 398286 147200 398342 148000 6 mgmt_soc_dff_Do[25]
port 633 nsew signal input
rlabel metal3 s 399200 130976 400000 131096 6 mgmt_soc_dff_Do[26]
port 634 nsew signal input
rlabel metal2 s 394882 0 394938 800 6 mgmt_soc_dff_Do[27]
port 635 nsew signal input
rlabel metal2 s 399574 147200 399630 148000 6 mgmt_soc_dff_Do[28]
port 636 nsew signal input
rlabel metal3 s 399200 144440 400000 144560 6 mgmt_soc_dff_Do[29]
port 637 nsew signal input
rlabel metal3 s 0 100512 800 100632 6 mgmt_soc_dff_Do[2]
port 638 nsew signal input
rlabel metal3 s 0 141720 800 141840 6 mgmt_soc_dff_Do[30]
port 639 nsew signal input
rlabel metal3 s 0 146616 800 146736 6 mgmt_soc_dff_Do[31]
port 640 nsew signal input
rlabel metal3 s 0 105272 800 105392 6 mgmt_soc_dff_Do[3]
port 641 nsew signal input
rlabel metal2 s 389178 147200 389234 148000 6 mgmt_soc_dff_Do[4]
port 642 nsew signal input
rlabel metal2 s 364706 0 364762 800 6 mgmt_soc_dff_Do[5]
port 643 nsew signal input
rlabel metal2 s 391202 147200 391258 148000 6 mgmt_soc_dff_Do[6]
port 644 nsew signal input
rlabel metal2 s 392490 147200 392546 148000 6 mgmt_soc_dff_Do[7]
port 645 nsew signal input
rlabel metal3 s 399200 56992 400000 57112 6 mgmt_soc_dff_Do[8]
port 646 nsew signal input
rlabel metal2 s 371422 0 371478 800 6 mgmt_soc_dff_Do[9]
port 647 nsew signal input
rlabel metal3 s 0 88408 800 88528 6 mgmt_soc_dff_EN
port 648 nsew signal output
rlabel metal3 s 0 98064 800 98184 6 mgmt_soc_dff_WE[0]
port 649 nsew signal output
rlabel metal2 s 347870 0 347926 800 6 mgmt_soc_dff_WE[1]
port 650 nsew signal output
rlabel metal2 s 387890 147200 387946 148000 6 mgmt_soc_dff_WE[2]
port 651 nsew signal output
rlabel metal2 s 361302 0 361358 800 6 mgmt_soc_dff_WE[3]
port 652 nsew signal output
rlabel metal3 s 0 83512 800 83632 6 mprj_ack_i
port 653 nsew signal input
rlabel metal2 s 336554 147200 336610 148000 6 mprj_adr_o[0]
port 654 nsew signal output
rlabel metal2 s 352102 147200 352158 148000 6 mprj_adr_o[10]
port 655 nsew signal output
rlabel metal2 s 353390 147200 353446 148000 6 mprj_adr_o[11]
port 656 nsew signal output
rlabel metal2 s 354770 147200 354826 148000 6 mprj_adr_o[12]
port 657 nsew signal output
rlabel metal2 s 356058 147200 356114 148000 6 mprj_adr_o[13]
port 658 nsew signal output
rlabel metal2 s 357346 147200 357402 148000 6 mprj_adr_o[14]
port 659 nsew signal output
rlabel metal2 s 358634 147200 358690 148000 6 mprj_adr_o[15]
port 660 nsew signal output
rlabel metal2 s 359922 147200 359978 148000 6 mprj_adr_o[16]
port 661 nsew signal output
rlabel metal2 s 361210 147200 361266 148000 6 mprj_adr_o[17]
port 662 nsew signal output
rlabel metal2 s 362498 147200 362554 148000 6 mprj_adr_o[18]
port 663 nsew signal output
rlabel metal2 s 363878 147200 363934 148000 6 mprj_adr_o[19]
port 664 nsew signal output
rlabel metal2 s 338486 147200 338542 148000 6 mprj_adr_o[1]
port 665 nsew signal output
rlabel metal2 s 365166 147200 365222 148000 6 mprj_adr_o[20]
port 666 nsew signal output
rlabel metal2 s 366454 147200 366510 148000 6 mprj_adr_o[21]
port 667 nsew signal output
rlabel metal2 s 367742 147200 367798 148000 6 mprj_adr_o[22]
port 668 nsew signal output
rlabel metal2 s 369030 147200 369086 148000 6 mprj_adr_o[23]
port 669 nsew signal output
rlabel metal2 s 370318 147200 370374 148000 6 mprj_adr_o[24]
port 670 nsew signal output
rlabel metal2 s 371606 147200 371662 148000 6 mprj_adr_o[25]
port 671 nsew signal output
rlabel metal2 s 372986 147200 373042 148000 6 mprj_adr_o[26]
port 672 nsew signal output
rlabel metal2 s 374274 147200 374330 148000 6 mprj_adr_o[27]
port 673 nsew signal output
rlabel metal2 s 375562 147200 375618 148000 6 mprj_adr_o[28]
port 674 nsew signal output
rlabel metal2 s 376850 147200 376906 148000 6 mprj_adr_o[29]
port 675 nsew signal output
rlabel metal2 s 340418 147200 340474 148000 6 mprj_adr_o[2]
port 676 nsew signal output
rlabel metal2 s 378138 147200 378194 148000 6 mprj_adr_o[30]
port 677 nsew signal output
rlabel metal2 s 379426 147200 379482 148000 6 mprj_adr_o[31]
port 678 nsew signal output
rlabel metal2 s 342350 147200 342406 148000 6 mprj_adr_o[3]
port 679 nsew signal output
rlabel metal2 s 344282 147200 344338 148000 6 mprj_adr_o[4]
port 680 nsew signal output
rlabel metal2 s 345662 147200 345718 148000 6 mprj_adr_o[5]
port 681 nsew signal output
rlabel metal2 s 346950 147200 347006 148000 6 mprj_adr_o[6]
port 682 nsew signal output
rlabel metal2 s 348238 147200 348294 148000 6 mprj_adr_o[7]
port 683 nsew signal output
rlabel metal2 s 349526 147200 349582 148000 6 mprj_adr_o[8]
port 684 nsew signal output
rlabel metal2 s 350814 147200 350870 148000 6 mprj_adr_o[9]
port 685 nsew signal output
rlabel metal2 s 334530 147200 334586 148000 6 mprj_cyc_o
port 686 nsew signal output
rlabel metal3 s 0 5856 800 5976 6 mprj_dat_i[0]
port 687 nsew signal input
rlabel metal3 s 0 30200 800 30320 6 mprj_dat_i[10]
port 688 nsew signal input
rlabel metal3 s 0 32512 800 32632 6 mprj_dat_i[11]
port 689 nsew signal input
rlabel metal3 s 0 34960 800 35080 6 mprj_dat_i[12]
port 690 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 mprj_dat_i[13]
port 691 nsew signal input
rlabel metal3 s 0 39856 800 39976 6 mprj_dat_i[14]
port 692 nsew signal input
rlabel metal3 s 0 42304 800 42424 6 mprj_dat_i[15]
port 693 nsew signal input
rlabel metal3 s 0 44752 800 44872 6 mprj_dat_i[16]
port 694 nsew signal input
rlabel metal3 s 0 47064 800 47184 6 mprj_dat_i[17]
port 695 nsew signal input
rlabel metal3 s 0 49512 800 49632 6 mprj_dat_i[18]
port 696 nsew signal input
rlabel metal3 s 0 51960 800 52080 6 mprj_dat_i[19]
port 697 nsew signal input
rlabel metal3 s 0 8304 800 8424 6 mprj_dat_i[1]
port 698 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 mprj_dat_i[20]
port 699 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 mprj_dat_i[21]
port 700 nsew signal input
rlabel metal3 s 0 59304 800 59424 6 mprj_dat_i[22]
port 701 nsew signal input
rlabel metal3 s 0 61616 800 61736 6 mprj_dat_i[23]
port 702 nsew signal input
rlabel metal3 s 0 64064 800 64184 6 mprj_dat_i[24]
port 703 nsew signal input
rlabel metal3 s 0 66512 800 66632 6 mprj_dat_i[25]
port 704 nsew signal input
rlabel metal3 s 0 68960 800 69080 6 mprj_dat_i[26]
port 705 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 mprj_dat_i[27]
port 706 nsew signal input
rlabel metal3 s 0 73856 800 73976 6 mprj_dat_i[28]
port 707 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 mprj_dat_i[29]
port 708 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 mprj_dat_i[2]
port 709 nsew signal input
rlabel metal3 s 0 78616 800 78736 6 mprj_dat_i[30]
port 710 nsew signal input
rlabel metal3 s 0 81064 800 81184 6 mprj_dat_i[31]
port 711 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 mprj_dat_i[3]
port 712 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 mprj_dat_i[4]
port 713 nsew signal input
rlabel metal3 s 0 17960 800 18080 6 mprj_dat_i[5]
port 714 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 mprj_dat_i[6]
port 715 nsew signal input
rlabel metal3 s 0 22856 800 22976 6 mprj_dat_i[7]
port 716 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 mprj_dat_i[8]
port 717 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 mprj_dat_i[9]
port 718 nsew signal input
rlabel metal2 s 337198 147200 337254 148000 6 mprj_dat_o[0]
port 719 nsew signal output
rlabel metal2 s 352746 147200 352802 148000 6 mprj_dat_o[10]
port 720 nsew signal output
rlabel metal2 s 354126 147200 354182 148000 6 mprj_dat_o[11]
port 721 nsew signal output
rlabel metal2 s 355414 147200 355470 148000 6 mprj_dat_o[12]
port 722 nsew signal output
rlabel metal2 s 356702 147200 356758 148000 6 mprj_dat_o[13]
port 723 nsew signal output
rlabel metal2 s 357990 147200 358046 148000 6 mprj_dat_o[14]
port 724 nsew signal output
rlabel metal2 s 359278 147200 359334 148000 6 mprj_dat_o[15]
port 725 nsew signal output
rlabel metal2 s 360566 147200 360622 148000 6 mprj_dat_o[16]
port 726 nsew signal output
rlabel metal2 s 361854 147200 361910 148000 6 mprj_dat_o[17]
port 727 nsew signal output
rlabel metal2 s 363234 147200 363290 148000 6 mprj_dat_o[18]
port 728 nsew signal output
rlabel metal2 s 364522 147200 364578 148000 6 mprj_dat_o[19]
port 729 nsew signal output
rlabel metal2 s 339130 147200 339186 148000 6 mprj_dat_o[1]
port 730 nsew signal output
rlabel metal2 s 365810 147200 365866 148000 6 mprj_dat_o[20]
port 731 nsew signal output
rlabel metal2 s 367098 147200 367154 148000 6 mprj_dat_o[21]
port 732 nsew signal output
rlabel metal2 s 368386 147200 368442 148000 6 mprj_dat_o[22]
port 733 nsew signal output
rlabel metal2 s 369674 147200 369730 148000 6 mprj_dat_o[23]
port 734 nsew signal output
rlabel metal2 s 370962 147200 371018 148000 6 mprj_dat_o[24]
port 735 nsew signal output
rlabel metal2 s 372250 147200 372306 148000 6 mprj_dat_o[25]
port 736 nsew signal output
rlabel metal2 s 373630 147200 373686 148000 6 mprj_dat_o[26]
port 737 nsew signal output
rlabel metal2 s 374918 147200 374974 148000 6 mprj_dat_o[27]
port 738 nsew signal output
rlabel metal2 s 376206 147200 376262 148000 6 mprj_dat_o[28]
port 739 nsew signal output
rlabel metal2 s 377494 147200 377550 148000 6 mprj_dat_o[29]
port 740 nsew signal output
rlabel metal2 s 341062 147200 341118 148000 6 mprj_dat_o[2]
port 741 nsew signal output
rlabel metal2 s 378782 147200 378838 148000 6 mprj_dat_o[30]
port 742 nsew signal output
rlabel metal2 s 380070 147200 380126 148000 6 mprj_dat_o[31]
port 743 nsew signal output
rlabel metal2 s 342994 147200 343050 148000 6 mprj_dat_o[3]
port 744 nsew signal output
rlabel metal2 s 345018 147200 345074 148000 6 mprj_dat_o[4]
port 745 nsew signal output
rlabel metal2 s 346306 147200 346362 148000 6 mprj_dat_o[5]
port 746 nsew signal output
rlabel metal2 s 347594 147200 347650 148000 6 mprj_dat_o[6]
port 747 nsew signal output
rlabel metal2 s 348882 147200 348938 148000 6 mprj_dat_o[7]
port 748 nsew signal output
rlabel metal2 s 350170 147200 350226 148000 6 mprj_dat_o[8]
port 749 nsew signal output
rlabel metal2 s 351458 147200 351514 148000 6 mprj_dat_o[9]
port 750 nsew signal output
rlabel metal2 s 337842 147200 337898 148000 6 mprj_sel_o[0]
port 751 nsew signal output
rlabel metal2 s 339774 147200 339830 148000 6 mprj_sel_o[1]
port 752 nsew signal output
rlabel metal2 s 341706 147200 341762 148000 6 mprj_sel_o[2]
port 753 nsew signal output
rlabel metal2 s 343638 147200 343694 148000 6 mprj_sel_o[3]
port 754 nsew signal output
rlabel metal2 s 335266 147200 335322 148000 6 mprj_stb_o
port 755 nsew signal output
rlabel metal2 s 380714 147200 380770 148000 6 mprj_wb_iena
port 756 nsew signal output
rlabel metal2 s 335910 147200 335966 148000 6 mprj_we_o
port 757 nsew signal output
rlabel metal2 s 58806 0 58862 800 6 qspi_enabled
port 758 nsew signal output
rlabel metal3 s 0 90720 800 90840 6 serial_rx
port 759 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 serial_tx
port 760 nsew signal output
rlabel metal2 s 384670 147200 384726 148000 6 spi_clk
port 761 nsew signal output
rlabel metal2 s 385314 147200 385370 148000 6 spi_cs_n
port 762 nsew signal output
rlabel metal2 s 324318 0 324374 800 6 spi_enabled
port 763 nsew signal output
rlabel metal2 s 341154 0 341210 800 6 spi_miso
port 764 nsew signal input
rlabel metal3 s 0 95616 800 95736 6 spi_mosi
port 765 nsew signal output
rlabel metal2 s 327722 0 327778 800 6 spi_sdoenb
port 766 nsew signal output
rlabel metal2 s 183190 0 183246 800 6 sram_ro_addr[0]
port 767 nsew signal output
rlabel metal2 s 186502 0 186558 800 6 sram_ro_addr[1]
port 768 nsew signal output
rlabel metal2 s 189906 0 189962 800 6 sram_ro_addr[2]
port 769 nsew signal output
rlabel metal2 s 193218 0 193274 800 6 sram_ro_addr[3]
port 770 nsew signal output
rlabel metal2 s 196622 0 196678 800 6 sram_ro_addr[4]
port 771 nsew signal output
rlabel metal2 s 199934 0 199990 800 6 sram_ro_addr[5]
port 772 nsew signal output
rlabel metal2 s 203338 0 203394 800 6 sram_ro_addr[6]
port 773 nsew signal output
rlabel metal2 s 206650 0 206706 800 6 sram_ro_addr[7]
port 774 nsew signal output
rlabel metal2 s 176382 0 176438 800 6 sram_ro_clk
port 775 nsew signal output
rlabel metal2 s 179786 0 179842 800 6 sram_ro_csb
port 776 nsew signal output
rlabel metal2 s 210054 0 210110 800 6 sram_ro_data[0]
port 777 nsew signal output
rlabel metal2 s 243634 0 243690 800 6 sram_ro_data[10]
port 778 nsew signal output
rlabel metal2 s 247038 0 247094 800 6 sram_ro_data[11]
port 779 nsew signal output
rlabel metal2 s 250350 0 250406 800 6 sram_ro_data[12]
port 780 nsew signal output
rlabel metal2 s 253754 0 253810 800 6 sram_ro_data[13]
port 781 nsew signal output
rlabel metal2 s 257066 0 257122 800 6 sram_ro_data[14]
port 782 nsew signal output
rlabel metal2 s 260470 0 260526 800 6 sram_ro_data[15]
port 783 nsew signal output
rlabel metal2 s 263782 0 263838 800 6 sram_ro_data[16]
port 784 nsew signal output
rlabel metal2 s 267186 0 267242 800 6 sram_ro_data[17]
port 785 nsew signal output
rlabel metal2 s 270590 0 270646 800 6 sram_ro_data[18]
port 786 nsew signal output
rlabel metal2 s 273902 0 273958 800 6 sram_ro_data[19]
port 787 nsew signal output
rlabel metal2 s 213366 0 213422 800 6 sram_ro_data[1]
port 788 nsew signal output
rlabel metal2 s 277306 0 277362 800 6 sram_ro_data[20]
port 789 nsew signal output
rlabel metal2 s 280618 0 280674 800 6 sram_ro_data[21]
port 790 nsew signal output
rlabel metal2 s 284022 0 284078 800 6 sram_ro_data[22]
port 791 nsew signal output
rlabel metal2 s 287334 0 287390 800 6 sram_ro_data[23]
port 792 nsew signal output
rlabel metal2 s 290738 0 290794 800 6 sram_ro_data[24]
port 793 nsew signal output
rlabel metal2 s 294050 0 294106 800 6 sram_ro_data[25]
port 794 nsew signal output
rlabel metal2 s 297454 0 297510 800 6 sram_ro_data[26]
port 795 nsew signal output
rlabel metal2 s 300766 0 300822 800 6 sram_ro_data[27]
port 796 nsew signal output
rlabel metal2 s 304170 0 304226 800 6 sram_ro_data[28]
port 797 nsew signal output
rlabel metal2 s 307482 0 307538 800 6 sram_ro_data[29]
port 798 nsew signal output
rlabel metal2 s 216770 0 216826 800 6 sram_ro_data[2]
port 799 nsew signal output
rlabel metal2 s 310886 0 310942 800 6 sram_ro_data[30]
port 800 nsew signal output
rlabel metal2 s 314290 0 314346 800 6 sram_ro_data[31]
port 801 nsew signal output
rlabel metal2 s 220082 0 220138 800 6 sram_ro_data[3]
port 802 nsew signal output
rlabel metal2 s 223486 0 223542 800 6 sram_ro_data[4]
port 803 nsew signal output
rlabel metal2 s 226890 0 226946 800 6 sram_ro_data[5]
port 804 nsew signal output
rlabel metal2 s 230202 0 230258 800 6 sram_ro_data[6]
port 805 nsew signal output
rlabel metal2 s 233606 0 233662 800 6 sram_ro_data[7]
port 806 nsew signal output
rlabel metal2 s 236918 0 236974 800 6 sram_ro_data[8]
port 807 nsew signal output
rlabel metal2 s 240322 0 240378 800 6 sram_ro_data[9]
port 808 nsew signal output
rlabel metal2 s 331034 0 331090 800 6 trap
port 809 nsew signal output
rlabel metal2 s 334438 0 334494 800 6 uart_enabled
port 810 nsew signal output
rlabel metal3 s 399200 9936 400000 10056 6 user_irq[0]
port 811 nsew signal input
rlabel metal3 s 399200 30064 400000 30184 6 user_irq[1]
port 812 nsew signal input
rlabel metal2 s 354586 0 354642 800 6 user_irq[2]
port 813 nsew signal input
rlabel metal2 s 388534 147200 388590 148000 6 user_irq[3]
port 814 nsew signal input
rlabel metal2 s 389822 147200 389878 148000 6 user_irq[4]
port 815 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 user_irq[5]
port 816 nsew signal input
rlabel metal2 s 381358 147200 381414 148000 6 user_irq_ena[0]
port 817 nsew signal output
rlabel metal2 s 382094 147200 382150 148000 6 user_irq_ena[1]
port 818 nsew signal output
rlabel metal2 s 382738 147200 382794 148000 6 user_irq_ena[2]
port 819 nsew signal output
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 400000 148000
string LEFview TRUE
string GDS_FILE ../gds/mgmt_core.gds
string GDS_END 108153158
string GDS_START 16753480
<< end >>

