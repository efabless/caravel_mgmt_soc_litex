VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM128
  CLASS BLOCK ;
  FOREIGN RAM128 ;
  ORIGIN 0.000 0.000 ;
  SIZE 402.500 BY 470.560 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.500 215.600 402.500 216.200 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.500 254.360 402.500 254.960 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.500 293.120 402.500 293.720 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.500 331.880 402.500 332.480 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.500 370.640 402.500 371.240 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.500 409.400 402.500 410.000 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.500 448.160 402.500 448.760 ;
    END
  END A0[6]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 2.000 235.240 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 0.000 207.370 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 0.000 219.790 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 0.000 244.630 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 0.000 257.050 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 0.000 269.470 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 0.000 281.890 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 0.000 294.310 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 0.000 306.730 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 0.000 319.150 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 0.000 381.250 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 0.000 393.670 2.000 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 2.000 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 2.000 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 2.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 468.560 8.650 470.560 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.570 468.560 132.850 470.560 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 468.560 145.270 470.560 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 468.560 157.690 470.560 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 468.560 170.110 470.560 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 468.560 182.530 470.560 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 468.560 194.950 470.560 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.090 468.560 207.370 470.560 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 468.560 219.790 470.560 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 468.560 232.210 470.560 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 468.560 244.630 470.560 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 468.560 21.070 470.560 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.770 468.560 257.050 470.560 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.190 468.560 269.470 470.560 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.610 468.560 281.890 470.560 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 468.560 294.310 470.560 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 468.560 306.730 470.560 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 468.560 319.150 470.560 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.290 468.560 331.570 470.560 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 468.560 343.990 470.560 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 468.560 356.410 470.560 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 468.560 368.830 470.560 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 468.560 33.490 470.560 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 468.560 381.250 470.560 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.390 468.560 393.670 470.560 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.630 468.560 45.910 470.560 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 468.560 58.330 470.560 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 468.560 70.750 470.560 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.890 468.560 83.170 470.560 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.310 468.560 95.590 470.560 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.730 468.560 108.010 470.560 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 468.560 120.430 470.560 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.500 21.800 402.500 22.400 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 468.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.680 2.480 250.280 468.080 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 468.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 468.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 468.080 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.500 60.560 402.500 61.160 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.500 99.320 402.500 99.920 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.500 138.080 402.500 138.680 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 400.500 176.840 402.500 177.440 ;
    END
  END WE0[3]
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 399.740 467.925 ;
      LAYER met1 ;
        RECT 0.990 0.380 402.430 470.520 ;
      LAYER met2 ;
        RECT 1.020 468.280 8.090 470.550 ;
        RECT 8.930 468.280 20.510 470.550 ;
        RECT 21.350 468.280 32.930 470.550 ;
        RECT 33.770 468.280 45.350 470.550 ;
        RECT 46.190 468.280 57.770 470.550 ;
        RECT 58.610 468.280 70.190 470.550 ;
        RECT 71.030 468.280 82.610 470.550 ;
        RECT 83.450 468.280 95.030 470.550 ;
        RECT 95.870 468.280 107.450 470.550 ;
        RECT 108.290 468.280 119.870 470.550 ;
        RECT 120.710 468.280 132.290 470.550 ;
        RECT 133.130 468.280 144.710 470.550 ;
        RECT 145.550 468.280 157.130 470.550 ;
        RECT 157.970 468.280 169.550 470.550 ;
        RECT 170.390 468.280 181.970 470.550 ;
        RECT 182.810 468.280 194.390 470.550 ;
        RECT 195.230 468.280 206.810 470.550 ;
        RECT 207.650 468.280 219.230 470.550 ;
        RECT 220.070 468.280 231.650 470.550 ;
        RECT 232.490 468.280 244.070 470.550 ;
        RECT 244.910 468.280 256.490 470.550 ;
        RECT 257.330 468.280 268.910 470.550 ;
        RECT 269.750 468.280 281.330 470.550 ;
        RECT 282.170 468.280 293.750 470.550 ;
        RECT 294.590 468.280 306.170 470.550 ;
        RECT 307.010 468.280 318.590 470.550 ;
        RECT 319.430 468.280 331.010 470.550 ;
        RECT 331.850 468.280 343.430 470.550 ;
        RECT 344.270 468.280 355.850 470.550 ;
        RECT 356.690 468.280 368.270 470.550 ;
        RECT 369.110 468.280 380.690 470.550 ;
        RECT 381.530 468.280 393.110 470.550 ;
        RECT 393.950 468.280 402.400 470.550 ;
        RECT 1.020 2.280 402.400 468.280 ;
        RECT 1.020 0.350 8.090 2.280 ;
        RECT 8.930 0.350 20.510 2.280 ;
        RECT 21.350 0.350 32.930 2.280 ;
        RECT 33.770 0.350 45.350 2.280 ;
        RECT 46.190 0.350 57.770 2.280 ;
        RECT 58.610 0.350 70.190 2.280 ;
        RECT 71.030 0.350 82.610 2.280 ;
        RECT 83.450 0.350 95.030 2.280 ;
        RECT 95.870 0.350 107.450 2.280 ;
        RECT 108.290 0.350 119.870 2.280 ;
        RECT 120.710 0.350 132.290 2.280 ;
        RECT 133.130 0.350 144.710 2.280 ;
        RECT 145.550 0.350 157.130 2.280 ;
        RECT 157.970 0.350 169.550 2.280 ;
        RECT 170.390 0.350 181.970 2.280 ;
        RECT 182.810 0.350 194.390 2.280 ;
        RECT 195.230 0.350 206.810 2.280 ;
        RECT 207.650 0.350 219.230 2.280 ;
        RECT 220.070 0.350 231.650 2.280 ;
        RECT 232.490 0.350 244.070 2.280 ;
        RECT 244.910 0.350 256.490 2.280 ;
        RECT 257.330 0.350 268.910 2.280 ;
        RECT 269.750 0.350 281.330 2.280 ;
        RECT 282.170 0.350 293.750 2.280 ;
        RECT 294.590 0.350 306.170 2.280 ;
        RECT 307.010 0.350 318.590 2.280 ;
        RECT 319.430 0.350 331.010 2.280 ;
        RECT 331.850 0.350 343.430 2.280 ;
        RECT 344.270 0.350 355.850 2.280 ;
        RECT 356.690 0.350 368.270 2.280 ;
        RECT 369.110 0.350 380.690 2.280 ;
        RECT 381.530 0.350 393.110 2.280 ;
        RECT 393.950 0.350 402.400 2.280 ;
      LAYER met3 ;
        RECT 2.000 449.160 401.975 470.540 ;
        RECT 2.000 447.760 400.100 449.160 ;
        RECT 2.000 410.400 401.975 447.760 ;
        RECT 2.000 409.000 400.100 410.400 ;
        RECT 2.000 371.640 401.975 409.000 ;
        RECT 2.000 370.240 400.100 371.640 ;
        RECT 2.000 332.880 401.975 370.240 ;
        RECT 2.000 331.480 400.100 332.880 ;
        RECT 2.000 294.120 401.975 331.480 ;
        RECT 2.000 292.720 400.100 294.120 ;
        RECT 2.000 255.360 401.975 292.720 ;
        RECT 2.000 253.960 400.100 255.360 ;
        RECT 2.000 235.640 401.975 253.960 ;
        RECT 2.400 234.240 401.975 235.640 ;
        RECT 2.000 216.600 401.975 234.240 ;
        RECT 2.000 215.200 400.100 216.600 ;
        RECT 2.000 177.840 401.975 215.200 ;
        RECT 2.000 176.440 400.100 177.840 ;
        RECT 2.000 139.080 401.975 176.440 ;
        RECT 2.000 137.680 400.100 139.080 ;
        RECT 2.000 100.320 401.975 137.680 ;
        RECT 2.000 98.920 400.100 100.320 ;
        RECT 2.000 61.560 401.975 98.920 ;
        RECT 2.000 60.160 400.100 61.560 ;
        RECT 2.000 22.800 401.975 60.160 ;
        RECT 2.000 21.400 400.100 22.800 ;
        RECT 2.000 0.855 401.975 21.400 ;
      LAYER met4 ;
        RECT 11.335 468.480 394.385 470.385 ;
        RECT 11.335 17.175 17.880 468.480 ;
        RECT 20.280 17.175 94.680 468.480 ;
        RECT 97.080 17.175 171.480 468.480 ;
        RECT 173.880 17.175 248.280 468.480 ;
        RECT 250.680 17.175 325.080 468.480 ;
        RECT 327.480 17.175 394.385 468.480 ;
  END
END RAM128
END LIBRARY

