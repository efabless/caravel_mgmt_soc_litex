VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM256
  CLASS BLOCK ;
  FOREIGN RAM256 ;
  ORIGIN 0.000 0.000 ;
  SIZE 798.100 BY 402.560 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.100 170.040 798.100 170.640 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.100 200.640 798.100 201.240 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.100 231.240 798.100 231.840 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.100 261.840 798.100 262.440 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.100 292.440 798.100 293.040 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.100 323.040 798.100 323.640 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.100 353.640 798.100 354.240 ;
    END
  END A0[6]
  PIN A0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.100 384.240 798.100 384.840 ;
    END
  END A0[7]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 2.000 201.240 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 2.000 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 2.000 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 2.000 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 0.000 312.250 2.000 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 0.000 337.090 2.000 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 0.000 361.930 2.000 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 2.000 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 2.000 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 2.000 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 0.000 461.290 2.000 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 0.000 486.130 2.000 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 2.000 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 0.000 510.970 2.000 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 0.000 535.810 2.000 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 0.000 560.650 2.000 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 2.000 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.050 0.000 610.330 2.000 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 0.000 635.170 2.000 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.730 0.000 660.010 2.000 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.570 0.000 684.850 2.000 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 0.000 709.690 2.000 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 2.000 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 2.000 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 0.000 759.370 2.000 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.930 0.000 784.210 2.000 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 2.000 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 2.000 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 2.000 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 2.000 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 2.000 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 2.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 2.000 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 400.560 14.170 402.560 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 400.560 262.570 402.560 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 400.560 287.410 402.560 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 400.560 312.250 402.560 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 400.560 337.090 402.560 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 400.560 361.930 402.560 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 400.560 386.770 402.560 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 400.560 411.610 402.560 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 400.560 436.450 402.560 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 400.560 461.290 402.560 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 400.560 486.130 402.560 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 400.560 39.010 402.560 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 400.560 510.970 402.560 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 400.560 535.810 402.560 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 400.560 560.650 402.560 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 400.560 585.490 402.560 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.050 400.560 610.330 402.560 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 400.560 635.170 402.560 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.730 400.560 660.010 402.560 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.570 400.560 684.850 402.560 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 400.560 709.690 402.560 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 400.560 734.530 402.560 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 400.560 63.850 402.560 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 400.560 759.370 402.560 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.930 400.560 784.210 402.560 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 400.560 88.690 402.560 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 400.560 113.530 402.560 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 400.560 138.370 402.560 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 400.560 163.210 402.560 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 400.560 188.050 402.560 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 400.560 212.890 402.560 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 400.560 237.730 402.560 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.100 17.040 798.100 17.640 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 95.080 2.480 96.680 400.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 248.680 2.480 250.280 400.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 402.280 2.480 403.880 400.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 555.880 2.480 557.480 400.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 709.480 2.480 711.080 400.080 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.280 2.480 19.880 400.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.880 2.480 173.480 400.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.480 2.480 327.080 400.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 479.080 2.480 480.680 400.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.680 2.480 634.280 400.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 786.280 2.480 787.880 400.080 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.100 47.640 798.100 48.240 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.100 78.240 798.100 78.840 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.100 108.840 798.100 109.440 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 796.100 139.440 798.100 140.040 ;
    END
  END WE0[3]
  OBS
      LAYER li1 ;
        RECT 2.760 2.635 795.340 399.925 ;
      LAYER met1 ;
        RECT 1.450 0.380 798.030 402.520 ;
      LAYER met2 ;
        RECT 1.470 400.280 13.610 402.550 ;
        RECT 14.450 400.280 38.450 402.550 ;
        RECT 39.290 400.280 63.290 402.550 ;
        RECT 64.130 400.280 88.130 402.550 ;
        RECT 88.970 400.280 112.970 402.550 ;
        RECT 113.810 400.280 137.810 402.550 ;
        RECT 138.650 400.280 162.650 402.550 ;
        RECT 163.490 400.280 187.490 402.550 ;
        RECT 188.330 400.280 212.330 402.550 ;
        RECT 213.170 400.280 237.170 402.550 ;
        RECT 238.010 400.280 262.010 402.550 ;
        RECT 262.850 400.280 286.850 402.550 ;
        RECT 287.690 400.280 311.690 402.550 ;
        RECT 312.530 400.280 336.530 402.550 ;
        RECT 337.370 400.280 361.370 402.550 ;
        RECT 362.210 400.280 386.210 402.550 ;
        RECT 387.050 400.280 411.050 402.550 ;
        RECT 411.890 400.280 435.890 402.550 ;
        RECT 436.730 400.280 460.730 402.550 ;
        RECT 461.570 400.280 485.570 402.550 ;
        RECT 486.410 400.280 510.410 402.550 ;
        RECT 511.250 400.280 535.250 402.550 ;
        RECT 536.090 400.280 560.090 402.550 ;
        RECT 560.930 400.280 584.930 402.550 ;
        RECT 585.770 400.280 609.770 402.550 ;
        RECT 610.610 400.280 634.610 402.550 ;
        RECT 635.450 400.280 659.450 402.550 ;
        RECT 660.290 400.280 684.290 402.550 ;
        RECT 685.130 400.280 709.130 402.550 ;
        RECT 709.970 400.280 733.970 402.550 ;
        RECT 734.810 400.280 758.810 402.550 ;
        RECT 759.650 400.280 783.650 402.550 ;
        RECT 784.490 400.280 798.000 402.550 ;
        RECT 1.470 2.280 798.000 400.280 ;
        RECT 1.470 0.155 13.610 2.280 ;
        RECT 14.450 0.155 38.450 2.280 ;
        RECT 39.290 0.155 63.290 2.280 ;
        RECT 64.130 0.155 88.130 2.280 ;
        RECT 88.970 0.155 112.970 2.280 ;
        RECT 113.810 0.155 137.810 2.280 ;
        RECT 138.650 0.155 162.650 2.280 ;
        RECT 163.490 0.155 187.490 2.280 ;
        RECT 188.330 0.155 212.330 2.280 ;
        RECT 213.170 0.155 237.170 2.280 ;
        RECT 238.010 0.155 262.010 2.280 ;
        RECT 262.850 0.155 286.850 2.280 ;
        RECT 287.690 0.155 311.690 2.280 ;
        RECT 312.530 0.155 336.530 2.280 ;
        RECT 337.370 0.155 361.370 2.280 ;
        RECT 362.210 0.155 386.210 2.280 ;
        RECT 387.050 0.155 411.050 2.280 ;
        RECT 411.890 0.155 435.890 2.280 ;
        RECT 436.730 0.155 460.730 2.280 ;
        RECT 461.570 0.155 485.570 2.280 ;
        RECT 486.410 0.155 510.410 2.280 ;
        RECT 511.250 0.155 535.250 2.280 ;
        RECT 536.090 0.155 560.090 2.280 ;
        RECT 560.930 0.155 584.930 2.280 ;
        RECT 585.770 0.155 609.770 2.280 ;
        RECT 610.610 0.155 634.610 2.280 ;
        RECT 635.450 0.155 659.450 2.280 ;
        RECT 660.290 0.155 684.290 2.280 ;
        RECT 685.130 0.155 709.130 2.280 ;
        RECT 709.970 0.155 733.970 2.280 ;
        RECT 734.810 0.155 758.810 2.280 ;
        RECT 759.650 0.155 783.650 2.280 ;
        RECT 784.490 0.155 798.000 2.280 ;
      LAYER met3 ;
        RECT 1.445 385.240 797.575 402.385 ;
        RECT 1.445 383.840 795.700 385.240 ;
        RECT 1.445 354.640 797.575 383.840 ;
        RECT 1.445 353.240 795.700 354.640 ;
        RECT 1.445 324.040 797.575 353.240 ;
        RECT 1.445 322.640 795.700 324.040 ;
        RECT 1.445 293.440 797.575 322.640 ;
        RECT 1.445 292.040 795.700 293.440 ;
        RECT 1.445 262.840 797.575 292.040 ;
        RECT 1.445 261.440 795.700 262.840 ;
        RECT 1.445 232.240 797.575 261.440 ;
        RECT 1.445 230.840 795.700 232.240 ;
        RECT 1.445 201.640 797.575 230.840 ;
        RECT 2.400 200.240 795.700 201.640 ;
        RECT 1.445 171.040 797.575 200.240 ;
        RECT 1.445 169.640 795.700 171.040 ;
        RECT 1.445 140.440 797.575 169.640 ;
        RECT 1.445 139.040 795.700 140.440 ;
        RECT 1.445 109.840 797.575 139.040 ;
        RECT 1.445 108.440 795.700 109.840 ;
        RECT 1.445 79.240 797.575 108.440 ;
        RECT 1.445 77.840 795.700 79.240 ;
        RECT 1.445 48.640 797.575 77.840 ;
        RECT 1.445 47.240 795.700 48.640 ;
        RECT 1.445 18.040 797.575 47.240 ;
        RECT 1.445 16.640 795.700 18.040 ;
        RECT 1.445 0.175 797.575 16.640 ;
      LAYER met4 ;
        RECT 5.815 400.480 785.385 402.385 ;
        RECT 5.815 4.255 17.880 400.480 ;
        RECT 20.280 4.255 94.680 400.480 ;
        RECT 97.080 4.255 171.480 400.480 ;
        RECT 173.880 4.255 248.280 400.480 ;
        RECT 250.680 4.255 325.080 400.480 ;
        RECT 327.480 4.255 401.880 400.480 ;
        RECT 404.280 4.255 478.680 400.480 ;
        RECT 481.080 4.255 555.480 400.480 ;
        RECT 557.880 4.255 632.280 400.480 ;
        RECT 634.680 4.255 709.080 400.480 ;
        RECT 711.480 4.255 785.385 400.480 ;
  END
END RAM256
END LIBRARY

