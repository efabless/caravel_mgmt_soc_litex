magic
tech sky130A
magscale 1 2
timestamp 1638474025
<< metal1 >>
rect 213178 160216 213184 160268
rect 213236 160256 213242 160268
rect 221182 160256 221188 160268
rect 213236 160228 221188 160256
rect 213236 160216 213242 160228
rect 221182 160216 221188 160228
rect 221240 160216 221246 160268
rect 126514 160080 126520 160132
rect 126572 160120 126578 160132
rect 134150 160120 134156 160132
rect 126572 160092 134156 160120
rect 126572 160080 126578 160092
rect 134150 160080 134156 160092
rect 134208 160080 134214 160132
rect 63402 160012 63408 160064
rect 63460 160052 63466 160064
rect 146478 160052 146484 160064
rect 63460 160024 146484 160052
rect 63460 160012 63466 160024
rect 146478 160012 146484 160024
rect 146536 160012 146542 160064
rect 146938 160012 146944 160064
rect 146996 160052 147002 160064
rect 154482 160052 154488 160064
rect 146996 160024 154488 160052
rect 146996 160012 147002 160024
rect 154482 160012 154488 160024
rect 154540 160012 154546 160064
rect 156782 160012 156788 160064
rect 156840 160052 156846 160064
rect 191742 160052 191748 160064
rect 156840 160024 191748 160052
rect 156840 160012 156846 160024
rect 191742 160012 191748 160024
rect 191800 160012 191806 160064
rect 197170 160012 197176 160064
rect 197228 160052 197234 160064
rect 207014 160052 207020 160064
rect 197228 160024 207020 160052
rect 197228 160012 197234 160024
rect 207014 160012 207020 160024
rect 207072 160012 207078 160064
rect 211430 160012 211436 160064
rect 211488 160052 211494 160064
rect 280338 160052 280344 160064
rect 211488 160024 280344 160052
rect 211488 160012 211494 160024
rect 280338 160012 280344 160024
rect 280396 160012 280402 160064
rect 281258 160012 281264 160064
rect 281316 160052 281322 160064
rect 332686 160052 332692 160064
rect 281316 160024 332692 160052
rect 281316 160012 281322 160024
rect 332686 160012 332692 160024
rect 332744 160012 332750 160064
rect 334250 160012 334256 160064
rect 334308 160052 334314 160064
rect 374086 160052 374092 160064
rect 334308 160024 374092 160052
rect 334308 160012 334314 160024
rect 374086 160012 374092 160024
rect 374144 160012 374150 160064
rect 378870 160012 378876 160064
rect 378928 160052 378934 160064
rect 398098 160052 398104 160064
rect 378928 160024 398104 160052
rect 378928 160012 378934 160024
rect 398098 160012 398104 160024
rect 398156 160012 398162 160064
rect 409966 160012 409972 160064
rect 410024 160052 410030 160064
rect 417878 160052 417884 160064
rect 410024 160024 417884 160052
rect 410024 160012 410030 160024
rect 417878 160012 417884 160024
rect 417936 160012 417942 160064
rect 25590 159944 25596 159996
rect 25648 159984 25654 159996
rect 109770 159984 109776 159996
rect 25648 159956 109776 159984
rect 25648 159944 25654 159956
rect 109770 159944 109776 159956
rect 109828 159944 109834 159996
rect 117222 159944 117228 159996
rect 117280 159984 117286 159996
rect 191466 159984 191472 159996
rect 117280 159956 191472 159984
rect 117280 159944 117286 159956
rect 191466 159944 191472 159956
rect 191524 159944 191530 159996
rect 197998 159944 198004 159996
rect 198056 159984 198062 159996
rect 269114 159984 269120 159996
rect 198056 159956 269120 159984
rect 198056 159944 198062 159956
rect 269114 159944 269120 159956
rect 269172 159944 269178 159996
rect 271230 159944 271236 159996
rect 271288 159984 271294 159996
rect 272794 159984 272800 159996
rect 271288 159956 272800 159984
rect 271288 159944 271294 159956
rect 272794 159944 272800 159956
rect 272852 159944 272858 159996
rect 275370 159944 275376 159996
rect 275428 159984 275434 159996
rect 328454 159984 328460 159996
rect 275428 159956 328460 159984
rect 275428 159944 275434 159956
rect 328454 159944 328460 159956
rect 328512 159944 328518 159996
rect 329190 159944 329196 159996
rect 329248 159984 329254 159996
rect 369946 159984 369952 159996
rect 329248 159956 369952 159984
rect 329248 159944 329254 159956
rect 369946 159944 369952 159956
rect 370004 159944 370010 159996
rect 374638 159944 374644 159996
rect 374696 159984 374702 159996
rect 388346 159984 388352 159996
rect 374696 159956 388352 159984
rect 374696 159944 374702 159956
rect 388346 159944 388352 159956
rect 388404 159944 388410 159996
rect 389818 159944 389824 159996
rect 389876 159984 389882 159996
rect 413830 159984 413836 159996
rect 389876 159956 413836 159984
rect 389876 159944 389882 159956
rect 413830 159944 413836 159956
rect 413888 159944 413894 159996
rect 449526 159944 449532 159996
rect 449584 159984 449590 159996
rect 456150 159984 456156 159996
rect 449584 159956 456156 159984
rect 449584 159944 449590 159956
rect 456150 159944 456156 159956
rect 456208 159944 456214 159996
rect 457070 159944 457076 159996
rect 457128 159984 457134 159996
rect 463878 159984 463884 159996
rect 457128 159956 463884 159984
rect 457128 159944 457134 159956
rect 463878 159944 463884 159956
rect 463936 159944 463942 159996
rect 469674 159944 469680 159996
rect 469732 159984 469738 159996
rect 477402 159984 477408 159996
rect 469732 159956 477408 159984
rect 469732 159944 469738 159956
rect 477402 159944 477408 159956
rect 477460 159944 477466 159996
rect 76926 159876 76932 159928
rect 76984 159916 76990 159928
rect 162486 159916 162492 159928
rect 76984 159888 162492 159916
rect 76984 159876 76990 159888
rect 162486 159876 162492 159888
rect 162544 159876 162550 159928
rect 166902 159876 166908 159928
rect 166960 159916 166966 159928
rect 186406 159916 186412 159928
rect 166960 159888 186412 159916
rect 166960 159876 166966 159888
rect 186406 159876 186412 159888
rect 186464 159876 186470 159928
rect 191282 159876 191288 159928
rect 191340 159916 191346 159928
rect 264882 159916 264888 159928
rect 191340 159888 264888 159916
rect 191340 159876 191346 159888
rect 264882 159876 264888 159888
rect 264940 159876 264946 159928
rect 268654 159876 268660 159928
rect 268712 159916 268718 159928
rect 324038 159916 324044 159928
rect 268712 159888 324044 159916
rect 268712 159876 268718 159888
rect 324038 159876 324044 159888
rect 324096 159876 324102 159928
rect 328362 159876 328368 159928
rect 328420 159916 328426 159928
rect 369486 159916 369492 159928
rect 328420 159888 369492 159916
rect 328420 159876 328426 159888
rect 369486 159876 369492 159888
rect 369544 159876 369550 159928
rect 372154 159876 372160 159928
rect 372212 159916 372218 159928
rect 396166 159916 396172 159928
rect 372212 159888 396172 159916
rect 372212 159876 372218 159888
rect 396166 159876 396172 159888
rect 396224 159876 396230 159928
rect 403250 159876 403256 159928
rect 403308 159916 403314 159928
rect 416590 159916 416596 159928
rect 403308 159888 416596 159916
rect 403308 159876 403314 159888
rect 416590 159876 416596 159888
rect 416648 159876 416654 159928
rect 480622 159876 480628 159928
rect 480680 159916 480686 159928
rect 485958 159916 485964 159928
rect 480680 159888 485964 159916
rect 480680 159876 480686 159888
rect 485958 159876 485964 159888
rect 486016 159876 486022 159928
rect 70118 159808 70124 159860
rect 70176 159848 70182 159860
rect 153378 159848 153384 159860
rect 70176 159820 153384 159848
rect 70176 159808 70182 159820
rect 153378 159808 153384 159820
rect 153436 159808 153442 159860
rect 153470 159808 153476 159860
rect 153528 159848 153534 159860
rect 179414 159848 179420 159860
rect 153528 159820 179420 159848
rect 153528 159808 153534 159820
rect 179414 159808 179420 159820
rect 179472 159808 179478 159860
rect 184566 159808 184572 159860
rect 184624 159848 184630 159860
rect 259546 159848 259552 159860
rect 184624 159820 259552 159848
rect 184624 159808 184630 159820
rect 259546 159808 259552 159820
rect 259604 159808 259610 159860
rect 261938 159808 261944 159860
rect 261996 159848 262002 159860
rect 312354 159848 312360 159860
rect 261996 159820 312360 159848
rect 261996 159808 262002 159820
rect 312354 159808 312360 159820
rect 312412 159808 312418 159860
rect 312446 159808 312452 159860
rect 312504 159848 312510 159860
rect 313366 159848 313372 159860
rect 312504 159820 313372 159848
rect 312504 159808 312510 159820
rect 313366 159808 313372 159820
rect 313424 159808 313430 159860
rect 322474 159808 322480 159860
rect 322532 159848 322538 159860
rect 365162 159848 365168 159860
rect 322532 159820 365168 159848
rect 322532 159808 322538 159820
rect 365162 159808 365168 159820
rect 365220 159808 365226 159860
rect 376294 159808 376300 159860
rect 376352 159848 376358 159860
rect 406194 159848 406200 159860
rect 376352 159820 406200 159848
rect 376352 159808 376358 159820
rect 406194 159808 406200 159820
rect 406252 159808 406258 159860
rect 424318 159808 424324 159860
rect 424376 159848 424382 159860
rect 442718 159848 442724 159860
rect 424376 159820 442724 159848
rect 424376 159808 424382 159820
rect 442718 159808 442724 159820
rect 442776 159808 442782 159860
rect 450354 159808 450360 159860
rect 450412 159848 450418 159860
rect 456886 159848 456892 159860
rect 450412 159820 456892 159848
rect 450412 159808 450418 159820
rect 456886 159808 456892 159820
rect 456944 159808 456950 159860
rect 458726 159808 458732 159860
rect 458784 159848 458790 159860
rect 465074 159848 465080 159860
rect 458784 159820 465080 159848
rect 458784 159808 458790 159820
rect 465074 159808 465080 159820
rect 465132 159808 465138 159860
rect 468018 159808 468024 159860
rect 468076 159848 468082 159860
rect 476022 159848 476028 159860
rect 468076 159820 476028 159848
rect 468076 159808 468082 159820
rect 476022 159808 476028 159820
rect 476080 159808 476086 159860
rect 479794 159808 479800 159860
rect 479852 159848 479858 159860
rect 485222 159848 485228 159860
rect 479852 159820 485228 159848
rect 479852 159808 479858 159820
rect 485222 159808 485228 159820
rect 485280 159808 485286 159860
rect 56686 159740 56692 159792
rect 56744 159780 56750 159792
rect 131206 159780 131212 159792
rect 56744 159752 131212 159780
rect 56744 159740 56750 159752
rect 131206 159740 131212 159752
rect 131264 159740 131270 159792
rect 143258 159780 143264 159792
rect 131408 159752 143264 159780
rect 18874 159672 18880 159724
rect 18932 159712 18938 159724
rect 109126 159712 109132 159724
rect 18932 159684 109132 159712
rect 18932 159672 18938 159684
rect 109126 159672 109132 159684
rect 109184 159672 109190 159724
rect 113082 159672 113088 159724
rect 113140 159712 113146 159724
rect 126422 159712 126428 159724
rect 113140 159684 126428 159712
rect 113140 159672 113146 159684
rect 126422 159672 126428 159684
rect 126480 159672 126486 159724
rect 49970 159604 49976 159656
rect 50028 159644 50034 159656
rect 131408 159644 131436 159752
rect 143258 159740 143264 159752
rect 143316 159740 143322 159792
rect 143350 159740 143356 159792
rect 143408 159780 143414 159792
rect 160094 159780 160100 159792
rect 143408 159752 160100 159780
rect 143408 159740 143414 159752
rect 160094 159740 160100 159752
rect 160152 159740 160158 159792
rect 171134 159740 171140 159792
rect 171192 159780 171198 159792
rect 173250 159780 173256 159792
rect 171192 159752 173256 159780
rect 171192 159740 171198 159752
rect 173250 159740 173256 159752
rect 173308 159740 173314 159792
rect 177850 159740 177856 159792
rect 177908 159780 177914 159792
rect 253934 159780 253940 159792
rect 177908 159752 253940 159780
rect 177908 159740 177914 159752
rect 253934 159740 253940 159752
rect 253992 159740 253998 159792
rect 255222 159740 255228 159792
rect 255280 159780 255286 159792
rect 313458 159780 313464 159792
rect 255280 159752 313464 159780
rect 255280 159740 255286 159752
rect 313458 159740 313464 159752
rect 313516 159740 313522 159792
rect 314102 159740 314108 159792
rect 314160 159780 314166 159792
rect 357986 159780 357992 159792
rect 314160 159752 357992 159780
rect 314160 159740 314166 159752
rect 357986 159740 357992 159752
rect 358044 159740 358050 159792
rect 365438 159740 365444 159792
rect 365496 159780 365502 159792
rect 395522 159780 395528 159792
rect 365496 159752 395528 159780
rect 365496 159740 365502 159752
rect 395522 159740 395528 159752
rect 395580 159740 395586 159792
rect 396534 159740 396540 159792
rect 396592 159780 396598 159792
rect 413738 159780 413744 159792
rect 396592 159752 413744 159780
rect 396592 159740 396598 159752
rect 413738 159740 413744 159752
rect 413796 159740 413802 159792
rect 420914 159740 420920 159792
rect 420972 159780 420978 159792
rect 440418 159780 440424 159792
rect 420972 159752 440424 159780
rect 420972 159740 420978 159752
rect 440418 159740 440424 159752
rect 440476 159740 440482 159792
rect 134150 159672 134156 159724
rect 134208 159712 134214 159724
rect 156506 159712 156512 159724
rect 134208 159684 156512 159712
rect 134208 159672 134214 159684
rect 156506 159672 156512 159684
rect 156564 159672 156570 159724
rect 163774 159712 163780 159724
rect 156616 159684 163780 159712
rect 50028 159616 131436 159644
rect 50028 159604 50034 159616
rect 131666 159604 131672 159656
rect 131724 159644 131730 159656
rect 136542 159644 136548 159656
rect 131724 159616 136548 159644
rect 131724 159604 131730 159616
rect 136542 159604 136548 159616
rect 136600 159604 136606 159656
rect 136634 159604 136640 159656
rect 136692 159644 136698 159656
rect 139394 159644 139400 159656
rect 136692 159616 139400 159644
rect 136692 159604 136698 159616
rect 139394 159604 139400 159616
rect 139452 159604 139458 159656
rect 139946 159604 139952 159656
rect 140004 159644 140010 159656
rect 156616 159644 156644 159684
rect 163774 159672 163780 159684
rect 163832 159672 163838 159724
rect 167730 159672 167736 159724
rect 167788 159712 167794 159724
rect 246942 159712 246948 159724
rect 167788 159684 246948 159712
rect 167788 159672 167794 159684
rect 246942 159672 246948 159684
rect 247000 159672 247006 159724
rect 248506 159672 248512 159724
rect 248564 159712 248570 159724
rect 248564 159684 306374 159712
rect 248564 159672 248570 159684
rect 140004 159616 156644 159644
rect 140004 159604 140010 159616
rect 161014 159604 161020 159656
rect 161072 159644 161078 159656
rect 240226 159644 240232 159656
rect 161072 159616 240232 159644
rect 161072 159604 161078 159616
rect 240226 159604 240232 159616
rect 240284 159604 240290 159656
rect 244274 159604 244280 159656
rect 244332 159644 244338 159656
rect 305362 159644 305368 159656
rect 244332 159616 305368 159644
rect 244332 159604 244338 159616
rect 305362 159604 305368 159616
rect 305420 159604 305426 159656
rect 306346 159644 306374 159684
rect 308214 159672 308220 159724
rect 308272 159712 308278 159724
rect 342622 159712 342628 159724
rect 308272 159684 342628 159712
rect 308272 159672 308278 159684
rect 342622 159672 342628 159684
rect 342680 159672 342686 159724
rect 342714 159672 342720 159724
rect 342772 159712 342778 159724
rect 343818 159712 343824 159724
rect 342772 159684 343824 159712
rect 342772 159672 342778 159684
rect 343818 159672 343824 159684
rect 343876 159672 343882 159724
rect 347774 159672 347780 159724
rect 347832 159712 347838 159724
rect 378778 159712 378784 159724
rect 347832 159684 378784 159712
rect 347832 159672 347838 159684
rect 378778 159672 378784 159684
rect 378836 159672 378842 159724
rect 379698 159672 379704 159724
rect 379756 159712 379762 159724
rect 405826 159712 405832 159724
rect 379756 159684 405832 159712
rect 379756 159672 379762 159684
rect 405826 159672 405832 159684
rect 405884 159672 405890 159724
rect 417510 159672 417516 159724
rect 417568 159712 417574 159724
rect 437658 159712 437664 159724
rect 417568 159684 437664 159712
rect 417568 159672 417574 159684
rect 437658 159672 437664 159684
rect 437716 159672 437722 159724
rect 308582 159644 308588 159656
rect 306346 159616 308588 159644
rect 308582 159604 308588 159616
rect 308640 159604 308646 159656
rect 309042 159604 309048 159656
rect 309100 159644 309106 159656
rect 341610 159644 341616 159656
rect 309100 159616 341616 159644
rect 309100 159604 309106 159616
rect 341610 159604 341616 159616
rect 341668 159604 341674 159656
rect 342456 159616 342668 159644
rect 43254 159536 43260 159588
rect 43312 159576 43318 159588
rect 43312 159548 128354 159576
rect 43312 159536 43318 159548
rect 32306 159468 32312 159520
rect 32364 159508 32370 159520
rect 32364 159480 126376 159508
rect 32364 159468 32370 159480
rect 36538 159400 36544 159452
rect 36596 159440 36602 159452
rect 126238 159440 126244 159452
rect 36596 159412 126244 159440
rect 36596 159400 36602 159412
rect 126238 159400 126244 159412
rect 126296 159400 126302 159452
rect 126348 159440 126376 159480
rect 126422 159468 126428 159520
rect 126480 159508 126486 159520
rect 127802 159508 127808 159520
rect 126480 159480 127808 159508
rect 126480 159468 126486 159480
rect 127802 159468 127808 159480
rect 127860 159468 127866 159520
rect 128326 159508 128354 159548
rect 129918 159536 129924 159588
rect 129976 159576 129982 159588
rect 146938 159576 146944 159588
rect 129976 159548 146944 159576
rect 129976 159536 129982 159548
rect 146938 159536 146944 159548
rect 146996 159536 147002 159588
rect 153378 159536 153384 159588
rect 153436 159576 153442 159588
rect 156782 159576 156788 159588
rect 153436 159548 156788 159576
rect 153436 159536 153442 159548
rect 156782 159536 156788 159548
rect 156840 159536 156846 159588
rect 157610 159536 157616 159588
rect 157668 159576 157674 159588
rect 239306 159576 239312 159588
rect 157668 159548 239312 159576
rect 157668 159536 157674 159548
rect 239306 159536 239312 159548
rect 239364 159536 239370 159588
rect 250990 159536 250996 159588
rect 251048 159576 251054 159588
rect 310606 159576 310612 159588
rect 251048 159548 310612 159576
rect 251048 159536 251054 159548
rect 310606 159536 310612 159548
rect 310664 159536 310670 159588
rect 315758 159536 315764 159588
rect 315816 159576 315822 159588
rect 342456 159576 342484 159616
rect 315816 159548 342484 159576
rect 342640 159576 342668 159616
rect 342806 159604 342812 159656
rect 342864 159644 342870 159656
rect 354214 159644 354220 159656
rect 342864 159616 354220 159644
rect 342864 159604 342870 159616
rect 354214 159604 354220 159616
rect 354272 159604 354278 159656
rect 357434 159604 357440 159656
rect 357492 159644 357498 159656
rect 363138 159644 363144 159656
rect 357492 159616 363144 159644
rect 357492 159604 357498 159616
rect 363138 159604 363144 159616
rect 363196 159604 363202 159656
rect 369578 159604 369584 159656
rect 369636 159644 369642 159656
rect 401042 159644 401048 159656
rect 369636 159616 401048 159644
rect 369636 159604 369642 159616
rect 401042 159604 401048 159616
rect 401100 159604 401106 159656
rect 407482 159604 407488 159656
rect 407540 159644 407546 159656
rect 429930 159644 429936 159656
rect 407540 159616 429936 159644
rect 407540 159604 407546 159616
rect 429930 159604 429936 159616
rect 429988 159604 429994 159656
rect 478966 159604 478972 159656
rect 479024 159644 479030 159656
rect 484578 159644 484584 159656
rect 479024 159616 484584 159644
rect 479024 159604 479030 159616
rect 484578 159604 484584 159616
rect 484636 159604 484642 159656
rect 358906 159576 358912 159588
rect 342640 159548 358912 159576
rect 315816 159536 315822 159548
rect 358906 159536 358912 159548
rect 358964 159536 358970 159588
rect 362862 159536 362868 159588
rect 362920 159576 362926 159588
rect 394970 159576 394976 159588
rect 362920 159548 394976 159576
rect 362920 159536 362926 159548
rect 394970 159536 394976 159548
rect 395028 159536 395034 159588
rect 399018 159536 399024 159588
rect 399076 159576 399082 159588
rect 408494 159576 408500 159588
rect 399076 159548 408500 159576
rect 399076 159536 399082 159548
rect 408494 159536 408500 159548
rect 408552 159536 408558 159588
rect 410794 159536 410800 159588
rect 410852 159576 410858 159588
rect 432506 159576 432512 159588
rect 410852 159548 432512 159576
rect 410852 159536 410858 159548
rect 432506 159536 432512 159548
rect 432564 159536 432570 159588
rect 467190 159536 467196 159588
rect 467248 159576 467254 159588
rect 473354 159576 473360 159588
rect 467248 159548 473360 159576
rect 467248 159536 467254 159548
rect 473354 159536 473360 159548
rect 473412 159536 473418 159588
rect 131114 159508 131120 159520
rect 128326 159480 131120 159508
rect 131114 159468 131120 159480
rect 131172 159468 131178 159520
rect 131206 159468 131212 159520
rect 131264 159508 131270 159520
rect 144086 159508 144092 159520
rect 131264 159480 144092 159508
rect 131264 159468 131270 159480
rect 144086 159468 144092 159480
rect 144144 159468 144150 159520
rect 144178 159468 144184 159520
rect 144236 159508 144242 159520
rect 225322 159508 225328 159520
rect 144236 159480 225328 159508
rect 144236 159468 144242 159480
rect 225322 159468 225328 159480
rect 225380 159468 225386 159520
rect 230842 159468 230848 159520
rect 230900 159508 230906 159520
rect 293954 159508 293960 159520
rect 230900 159480 293960 159508
rect 230900 159468 230906 159480
rect 293954 159468 293960 159480
rect 294012 159468 294018 159520
rect 294782 159468 294788 159520
rect 294840 159508 294846 159520
rect 294840 159480 341564 159508
rect 294840 159468 294846 159480
rect 126790 159440 126796 159452
rect 126348 159412 126796 159440
rect 126790 159400 126796 159412
rect 126848 159400 126854 159452
rect 147490 159440 147496 159452
rect 128326 159412 147496 159440
rect 6270 159332 6276 159384
rect 6328 159372 6334 159384
rect 122834 159372 122840 159384
rect 6328 159344 122840 159372
rect 6328 159332 6334 159344
rect 122834 159332 122840 159344
rect 122892 159332 122898 159384
rect 123110 159332 123116 159384
rect 123168 159372 123174 159384
rect 128326 159372 128354 159412
rect 147490 159400 147496 159412
rect 147548 159400 147554 159452
rect 147582 159400 147588 159452
rect 147640 159440 147646 159452
rect 149514 159440 149520 159452
rect 147640 159412 149520 159440
rect 147640 159400 147646 159412
rect 149514 159400 149520 159412
rect 149572 159400 149578 159452
rect 150894 159400 150900 159452
rect 150952 159440 150958 159452
rect 233234 159440 233240 159452
rect 150952 159412 233240 159440
rect 150952 159400 150958 159412
rect 233234 159400 233240 159412
rect 233292 159400 233298 159452
rect 234982 159400 234988 159452
rect 235040 159440 235046 159452
rect 298002 159440 298008 159452
rect 235040 159412 298008 159440
rect 235040 159400 235046 159412
rect 298002 159400 298008 159412
rect 298060 159400 298066 159452
rect 301498 159400 301504 159452
rect 301556 159440 301562 159452
rect 341426 159440 341432 159452
rect 301556 159412 341432 159440
rect 301556 159400 301562 159412
rect 341426 159400 341432 159412
rect 341484 159400 341490 159452
rect 341536 159440 341564 159480
rect 341610 159468 341616 159520
rect 341668 159508 341674 159520
rect 354858 159508 354864 159520
rect 341668 159480 354864 159508
rect 341668 159468 341674 159480
rect 354858 159468 354864 159480
rect 354916 159468 354922 159520
rect 356146 159468 356152 159520
rect 356204 159508 356210 159520
rect 390554 159508 390560 159520
rect 356204 159480 390560 159508
rect 356204 159468 356210 159480
rect 390554 159468 390560 159480
rect 390612 159468 390618 159520
rect 400766 159468 400772 159520
rect 400824 159508 400830 159520
rect 424870 159508 424876 159520
rect 400824 159480 424876 159508
rect 400824 159468 400830 159480
rect 424870 159468 424876 159480
rect 424928 159468 424934 159520
rect 448698 159468 448704 159520
rect 448756 159508 448762 159520
rect 456058 159508 456064 159520
rect 448756 159480 456064 159508
rect 448756 159468 448762 159480
rect 456058 159468 456064 159480
rect 456116 159468 456122 159520
rect 457898 159468 457904 159520
rect 457956 159508 457962 159520
rect 464706 159508 464712 159520
rect 457956 159480 464712 159508
rect 457956 159468 457962 159480
rect 464706 159468 464712 159480
rect 464764 159468 464770 159520
rect 342254 159440 342260 159452
rect 341536 159412 342260 159440
rect 342254 159400 342260 159412
rect 342312 159400 342318 159452
rect 342346 159400 342352 159452
rect 342404 159440 342410 159452
rect 349338 159440 349344 159452
rect 342404 159412 349344 159440
rect 342404 159400 342410 159412
rect 349338 159400 349344 159412
rect 349396 159400 349402 159452
rect 358630 159400 358636 159452
rect 358688 159440 358694 159452
rect 392762 159440 392768 159452
rect 358688 159412 392768 159440
rect 358688 159400 358694 159412
rect 392762 159400 392768 159412
rect 392820 159400 392826 159452
rect 404078 159400 404084 159452
rect 404136 159440 404142 159452
rect 427354 159440 427360 159452
rect 404136 159412 427360 159440
rect 404136 159400 404142 159412
rect 427354 159400 427360 159412
rect 427412 159400 427418 159452
rect 427630 159400 427636 159452
rect 427688 159440 427694 159452
rect 445386 159440 445392 159452
rect 427688 159412 445392 159440
rect 427688 159400 427694 159412
rect 445386 159400 445392 159412
rect 445444 159400 445450 159452
rect 451182 159400 451188 159452
rect 451240 159440 451246 159452
rect 456794 159440 456800 159452
rect 451240 159412 456800 159440
rect 451240 159400 451246 159412
rect 456794 159400 456800 159412
rect 456852 159400 456858 159452
rect 459646 159400 459652 159452
rect 459704 159440 459710 159452
rect 466454 159440 466460 159452
rect 459704 159412 466460 159440
rect 459704 159400 459710 159412
rect 466454 159400 466460 159412
rect 466512 159400 466518 159452
rect 468846 159400 468852 159452
rect 468904 159440 468910 159452
rect 474826 159440 474832 159452
rect 468904 159412 474832 159440
rect 468904 159400 468910 159412
rect 474826 159400 474832 159412
rect 474884 159400 474890 159452
rect 477310 159400 477316 159452
rect 477368 159440 477374 159452
rect 483290 159440 483296 159452
rect 477368 159412 483296 159440
rect 477368 159400 477374 159412
rect 483290 159400 483296 159412
rect 483348 159400 483354 159452
rect 518802 159400 518808 159452
rect 518860 159440 518866 159452
rect 522666 159440 522672 159452
rect 518860 159412 522672 159440
rect 518860 159400 518866 159412
rect 522666 159400 522672 159412
rect 522724 159400 522730 159452
rect 123168 159344 128354 159372
rect 123168 159332 123174 159344
rect 129918 159332 129924 159384
rect 129976 159372 129982 159384
rect 137094 159372 137100 159384
rect 129976 159344 137100 159372
rect 129976 159332 129982 159344
rect 137094 159332 137100 159344
rect 137152 159332 137158 159384
rect 137462 159332 137468 159384
rect 137520 159372 137526 159384
rect 223574 159372 223580 159384
rect 137520 159344 223580 159372
rect 137520 159332 137526 159344
rect 223574 159332 223580 159344
rect 223632 159332 223638 159384
rect 231670 159332 231676 159384
rect 231728 159372 231734 159384
rect 295518 159372 295524 159384
rect 231728 159344 295524 159372
rect 231728 159332 231734 159344
rect 295518 159332 295524 159344
rect 295576 159332 295582 159384
rect 295610 159332 295616 159384
rect 295668 159372 295674 159384
rect 342438 159372 342444 159384
rect 295668 159344 342444 159372
rect 295668 159332 295674 159344
rect 342438 159332 342444 159344
rect 342496 159332 342502 159384
rect 346026 159332 346032 159384
rect 346084 159372 346090 159384
rect 382826 159372 382832 159384
rect 346084 159344 382832 159372
rect 346084 159332 346090 159344
rect 382826 159332 382832 159344
rect 382884 159332 382890 159384
rect 383102 159332 383108 159384
rect 383160 159372 383166 159384
rect 411346 159372 411352 159384
rect 383160 159344 411352 159372
rect 383160 159332 383166 159344
rect 411346 159332 411352 159344
rect 411404 159332 411410 159384
rect 414198 159332 414204 159384
rect 414256 159372 414262 159384
rect 435082 159372 435088 159384
rect 414256 159344 435088 159372
rect 414256 159332 414262 159344
rect 435082 159332 435088 159344
rect 435140 159332 435146 159384
rect 447870 159332 447876 159384
rect 447928 159372 447934 159384
rect 456978 159372 456984 159384
rect 447928 159344 456984 159372
rect 447928 159332 447934 159344
rect 456978 159332 456984 159344
rect 457036 159332 457042 159384
rect 470502 159332 470508 159384
rect 470560 159372 470566 159384
rect 476114 159372 476120 159384
rect 470560 159344 476120 159372
rect 470560 159332 470566 159344
rect 476114 159332 476120 159344
rect 476172 159332 476178 159384
rect 478138 159332 478144 159384
rect 478196 159372 478202 159384
rect 483198 159372 483204 159384
rect 478196 159344 483204 159372
rect 478196 159332 478202 159344
rect 483198 159332 483204 159344
rect 483256 159332 483262 159384
rect 518710 159332 518716 159384
rect 518768 159372 518774 159384
rect 523494 159372 523500 159384
rect 518768 159344 523500 159372
rect 518768 159332 518774 159344
rect 523494 159332 523500 159344
rect 523552 159332 523558 159384
rect 73522 159264 73528 159316
rect 73580 159304 73586 159316
rect 80054 159304 80060 159316
rect 73580 159276 80060 159304
rect 73580 159264 73586 159276
rect 80054 159264 80060 159276
rect 80112 159264 80118 159316
rect 83642 159264 83648 159316
rect 83700 159304 83706 159316
rect 166994 159304 167000 159316
rect 83700 159276 167000 159304
rect 83700 159264 83706 159276
rect 166994 159264 167000 159276
rect 167052 159264 167058 159316
rect 170214 159264 170220 159316
rect 170272 159304 170278 159316
rect 198918 159304 198924 159316
rect 170272 159276 198924 159304
rect 170272 159264 170278 159276
rect 198918 159264 198924 159276
rect 198976 159264 198982 159316
rect 201402 159264 201408 159316
rect 201460 159304 201466 159316
rect 212626 159304 212632 159316
rect 201460 159276 212632 159304
rect 201460 159264 201466 159276
rect 212626 159264 212632 159276
rect 212684 159264 212690 159316
rect 214006 159264 214012 159316
rect 214064 159304 214070 159316
rect 281534 159304 281540 159316
rect 214064 159276 281540 159304
rect 214064 159264 214070 159276
rect 281534 159264 281540 159276
rect 281592 159264 281598 159316
rect 282086 159264 282092 159316
rect 282144 159304 282150 159316
rect 334342 159304 334348 159316
rect 282144 159276 334348 159304
rect 282144 159264 282150 159276
rect 334342 159264 334348 159276
rect 334400 159264 334406 159316
rect 335078 159264 335084 159316
rect 335136 159304 335142 159316
rect 374730 159304 374736 159316
rect 335136 159276 374736 159304
rect 335136 159264 335142 159276
rect 374730 159264 374736 159276
rect 374788 159264 374794 159316
rect 388990 159264 388996 159316
rect 389048 159304 389054 159316
rect 403894 159304 403900 159316
rect 389048 159276 403900 159304
rect 389048 159264 389054 159276
rect 403894 159264 403900 159276
rect 403952 159264 403958 159316
rect 460474 159264 460480 159316
rect 460532 159304 460538 159316
rect 466638 159304 466644 159316
rect 460532 159276 466644 159304
rect 460532 159264 460538 159276
rect 466638 159264 466644 159276
rect 466696 159264 466702 159316
rect 80238 159196 80244 159248
rect 80296 159236 80302 159248
rect 91094 159236 91100 159248
rect 80296 159208 91100 159236
rect 80296 159196 80302 159208
rect 91094 159196 91100 159208
rect 91152 159196 91158 159248
rect 100478 159196 100484 159248
rect 100536 159236 100542 159248
rect 184382 159236 184388 159248
rect 100536 159208 184388 159236
rect 100536 159196 100542 159208
rect 184382 159196 184388 159208
rect 184440 159196 184446 159248
rect 187050 159196 187056 159248
rect 187108 159236 187114 159248
rect 214650 159236 214656 159248
rect 187108 159208 214656 159236
rect 187108 159196 187114 159208
rect 214650 159196 214656 159208
rect 214708 159196 214714 159248
rect 218238 159196 218244 159248
rect 218296 159236 218302 159248
rect 284386 159236 284392 159248
rect 218296 159208 284392 159236
rect 218296 159196 218302 159208
rect 284386 159196 284392 159208
rect 284444 159196 284450 159248
rect 287974 159196 287980 159248
rect 288032 159236 288038 159248
rect 338758 159236 338764 159248
rect 288032 159208 338764 159236
rect 288032 159196 288038 159208
rect 338758 159196 338764 159208
rect 338816 159196 338822 159248
rect 339310 159196 339316 159248
rect 339368 159236 339374 159248
rect 377950 159236 377956 159248
rect 339368 159208 377956 159236
rect 339368 159196 339374 159208
rect 377950 159196 377956 159208
rect 378008 159196 378014 159248
rect 385494 159236 385500 159248
rect 378796 159208 385500 159236
rect 86954 159128 86960 159180
rect 87012 159168 87018 159180
rect 87012 159140 162992 159168
rect 87012 159128 87018 159140
rect 93670 159060 93676 159112
rect 93728 159100 93734 159112
rect 162854 159100 162860 159112
rect 93728 159072 162860 159100
rect 93728 159060 93734 159072
rect 162854 159060 162860 159072
rect 162912 159060 162918 159112
rect 162964 159100 162992 159140
rect 163038 159128 163044 159180
rect 163096 159168 163102 159180
rect 172146 159168 172152 159180
rect 163096 159140 172152 159168
rect 163096 159128 163102 159140
rect 172146 159128 172152 159140
rect 172204 159128 172210 159180
rect 193766 159128 193772 159180
rect 193824 159168 193830 159180
rect 218054 159168 218060 159180
rect 193824 159140 218060 159168
rect 193824 159128 193830 159140
rect 218054 159128 218060 159140
rect 218112 159128 218118 159180
rect 224954 159128 224960 159180
rect 225012 159168 225018 159180
rect 290642 159168 290648 159180
rect 225012 159140 290648 159168
rect 225012 159128 225018 159140
rect 290642 159128 290648 159140
rect 290700 159128 290706 159180
rect 293954 159128 293960 159180
rect 294012 159168 294018 159180
rect 295150 159168 295156 159180
rect 294012 159140 295156 159168
rect 294012 159128 294018 159140
rect 295150 159128 295156 159140
rect 295208 159128 295214 159180
rect 302326 159128 302332 159180
rect 302384 159168 302390 159180
rect 302384 159140 340874 159168
rect 302384 159128 302390 159140
rect 169754 159100 169760 159112
rect 162964 159072 169760 159100
rect 169754 159060 169760 159072
rect 169812 159060 169818 159112
rect 173618 159060 173624 159112
rect 173676 159100 173682 159112
rect 197354 159100 197360 159112
rect 173676 159072 197360 159100
rect 173676 159060 173682 159072
rect 197354 159060 197360 159072
rect 197412 159060 197418 159112
rect 203886 159060 203892 159112
rect 203944 159100 203950 159112
rect 212718 159100 212724 159112
rect 203944 159072 212724 159100
rect 203944 159060 203950 159072
rect 212718 159060 212724 159072
rect 212776 159060 212782 159112
rect 220722 159060 220728 159112
rect 220780 159100 220786 159112
rect 283190 159100 283196 159112
rect 220780 159072 283196 159100
rect 220780 159060 220786 159072
rect 283190 159060 283196 159072
rect 283248 159060 283254 159112
rect 284662 159060 284668 159112
rect 284720 159100 284726 159112
rect 285766 159100 285772 159112
rect 284720 159072 285772 159100
rect 284720 159060 284726 159072
rect 285766 159060 285772 159072
rect 285824 159060 285830 159112
rect 288066 159100 288072 159112
rect 287026 159072 288072 159100
rect 107194 158992 107200 159044
rect 107252 159032 107258 159044
rect 183462 159032 183468 159044
rect 107252 159004 183468 159032
rect 107252 158992 107258 159004
rect 183462 158992 183468 159004
rect 183520 158992 183526 159044
rect 183738 158992 183744 159044
rect 183796 159032 183802 159044
rect 201402 159032 201408 159044
rect 183796 159004 201408 159032
rect 183796 158992 183802 159004
rect 201402 158992 201408 159004
rect 201460 158992 201466 159044
rect 214834 158992 214840 159044
rect 214892 159032 214898 159044
rect 222102 159032 222108 159044
rect 214892 159004 222108 159032
rect 214892 158992 214898 159004
rect 222102 158992 222108 159004
rect 222160 158992 222166 159044
rect 224126 158992 224132 159044
rect 224184 159032 224190 159044
rect 287026 159032 287054 159072
rect 288066 159060 288072 159072
rect 288124 159060 288130 159112
rect 288894 159060 288900 159112
rect 288952 159100 288958 159112
rect 338390 159100 338396 159112
rect 288952 159072 338396 159100
rect 288952 159060 288958 159072
rect 338390 159060 338396 159072
rect 338448 159060 338454 159112
rect 338482 159060 338488 159112
rect 338540 159100 338546 159112
rect 339678 159100 339684 159112
rect 338540 159072 339684 159100
rect 338540 159060 338546 159072
rect 339678 159060 339684 159072
rect 339736 159060 339742 159112
rect 340846 159100 340874 159140
rect 341426 159128 341432 159180
rect 341484 159168 341490 159180
rect 345658 159168 345664 159180
rect 341484 159140 345664 159168
rect 341484 159128 341490 159140
rect 345658 159128 345664 159140
rect 345716 159128 345722 159180
rect 345750 159128 345756 159180
rect 345808 159168 345814 159180
rect 351822 159168 351828 159180
rect 345808 159140 351828 159168
rect 345808 159128 345814 159140
rect 351822 159128 351828 159140
rect 351880 159128 351886 159180
rect 351914 159128 351920 159180
rect 351972 159168 351978 159180
rect 378796 159168 378824 159208
rect 385494 159196 385500 159208
rect 385552 159196 385558 159248
rect 385586 159196 385592 159248
rect 385644 159236 385650 159248
rect 398834 159236 398840 159248
rect 385644 159208 398840 159236
rect 385644 159196 385650 159208
rect 398834 159196 398840 159208
rect 398892 159196 398898 159248
rect 388438 159168 388444 159180
rect 351972 159140 378824 159168
rect 383626 159140 388444 159168
rect 351972 159128 351978 159140
rect 349246 159100 349252 159112
rect 340846 159072 349252 159100
rect 349246 159060 349252 159072
rect 349304 159060 349310 159112
rect 349338 159060 349344 159112
rect 349396 159100 349402 159112
rect 376938 159100 376944 159112
rect 349396 159072 376944 159100
rect 349396 159060 349402 159072
rect 376938 159060 376944 159072
rect 376996 159060 377002 159112
rect 378042 159060 378048 159112
rect 378100 159100 378106 159112
rect 383626 159100 383654 159140
rect 388438 159128 388444 159140
rect 388496 159128 388502 159180
rect 392302 159128 392308 159180
rect 392360 159168 392366 159180
rect 404262 159168 404268 159180
rect 392360 159140 404268 159168
rect 392360 159128 392366 159140
rect 404262 159128 404268 159140
rect 404320 159128 404326 159180
rect 461302 159128 461308 159180
rect 461360 159168 461366 159180
rect 467834 159168 467840 159180
rect 461360 159140 467840 159168
rect 461360 159128 461366 159140
rect 467834 159128 467840 159140
rect 467892 159128 467898 159180
rect 472250 159128 472256 159180
rect 472308 159168 472314 159180
rect 479426 159168 479432 159180
rect 472308 159140 479432 159168
rect 472308 159128 472314 159140
rect 479426 159128 479432 159140
rect 479484 159128 479490 159180
rect 378100 159072 383654 159100
rect 378100 159060 378106 159072
rect 395706 159060 395712 159112
rect 395764 159100 395770 159112
rect 404630 159100 404636 159112
rect 395764 159072 404636 159100
rect 395764 159060 395770 159072
rect 404630 159060 404636 159072
rect 404688 159060 404694 159112
rect 452010 159060 452016 159112
rect 452068 159100 452074 159112
rect 458174 159100 458180 159112
rect 452068 159072 458180 159100
rect 452068 159060 452074 159072
rect 458174 159060 458180 159072
rect 458232 159060 458238 159112
rect 462130 159060 462136 159112
rect 462188 159100 462194 159112
rect 467926 159100 467932 159112
rect 462188 159072 467932 159100
rect 462188 159060 462194 159072
rect 467926 159060 467932 159072
rect 467984 159060 467990 159112
rect 471422 159060 471428 159112
rect 471480 159100 471486 159112
rect 477678 159100 477684 159112
rect 471480 159072 477684 159100
rect 471480 159060 471486 159072
rect 477678 159060 477684 159072
rect 477736 159060 477742 159112
rect 224184 159004 287054 159032
rect 224184 158992 224190 159004
rect 298094 158992 298100 159044
rect 298152 159032 298158 159044
rect 300394 159032 300400 159044
rect 298152 159004 300400 159032
rect 298152 158992 298158 159004
rect 300394 158992 300400 159004
rect 300452 158992 300458 159044
rect 307386 158992 307392 159044
rect 307444 159032 307450 159044
rect 345566 159032 345572 159044
rect 307444 159004 345572 159032
rect 307444 158992 307450 159004
rect 345566 158992 345572 159004
rect 345624 158992 345630 159044
rect 345842 158992 345848 159044
rect 345900 159032 345906 159044
rect 349062 159032 349068 159044
rect 345900 159004 349068 159032
rect 345900 158992 345906 159004
rect 349062 158992 349068 159004
rect 349120 158992 349126 159044
rect 351086 158992 351092 159044
rect 351144 159032 351150 159044
rect 382550 159032 382556 159044
rect 351144 159004 382556 159032
rect 351144 158992 351150 159004
rect 382550 158992 382556 159004
rect 382608 158992 382614 159044
rect 455414 158992 455420 159044
rect 455472 159032 455478 159044
rect 463510 159032 463516 159044
rect 455472 159004 463516 159032
rect 455472 158992 455478 159004
rect 463510 158992 463516 159004
rect 463568 158992 463574 159044
rect 465534 158992 465540 159044
rect 465592 159032 465598 159044
rect 472526 159032 472532 159044
rect 465592 159004 472532 159032
rect 465592 158992 465598 159004
rect 472526 158992 472532 159004
rect 472584 158992 472590 159044
rect 473906 158992 473912 159044
rect 473964 159032 473970 159044
rect 480714 159032 480720 159044
rect 473964 159004 480720 159032
rect 473964 158992 473970 159004
rect 480714 158992 480720 159004
rect 480772 158992 480778 159044
rect 96246 158924 96252 158976
rect 96304 158964 96310 158976
rect 121914 158964 121920 158976
rect 96304 158936 121920 158964
rect 96304 158924 96310 158936
rect 121914 158924 121920 158936
rect 121972 158924 121978 158976
rect 124030 158924 124036 158976
rect 124088 158964 124094 158976
rect 194134 158964 194140 158976
rect 124088 158936 194140 158964
rect 124088 158924 124094 158936
rect 194134 158924 194140 158936
rect 194192 158924 194198 158976
rect 200574 158924 200580 158976
rect 200632 158964 200638 158976
rect 224954 158964 224960 158976
rect 200632 158936 224960 158964
rect 200632 158924 200638 158936
rect 224954 158924 224960 158936
rect 225012 158924 225018 158976
rect 237558 158924 237564 158976
rect 237616 158964 237622 158976
rect 299474 158964 299480 158976
rect 237616 158936 299480 158964
rect 237616 158924 237622 158936
rect 299474 158924 299480 158936
rect 299532 158924 299538 158976
rect 314930 158924 314936 158976
rect 314988 158964 314994 158976
rect 357526 158964 357532 158976
rect 314988 158936 357532 158964
rect 314988 158924 314994 158936
rect 357526 158924 357532 158936
rect 357584 158924 357590 158976
rect 357802 158924 357808 158976
rect 357860 158964 357866 158976
rect 384942 158964 384948 158976
rect 357860 158936 384948 158964
rect 357860 158924 357866 158936
rect 384942 158924 384948 158936
rect 385000 158924 385006 158976
rect 420086 158924 420092 158976
rect 420144 158964 420150 158976
rect 423490 158964 423496 158976
rect 420144 158936 423496 158964
rect 420144 158924 420150 158936
rect 423490 158924 423496 158936
rect 423548 158924 423554 158976
rect 446122 158924 446128 158976
rect 446180 158964 446186 158976
rect 453942 158964 453948 158976
rect 446180 158936 453948 158964
rect 446180 158924 446186 158936
rect 453942 158924 453948 158936
rect 454000 158924 454006 158976
rect 456242 158924 456248 158976
rect 456300 158964 456306 158976
rect 463602 158964 463608 158976
rect 456300 158936 463608 158964
rect 456300 158924 456306 158936
rect 463602 158924 463608 158936
rect 463660 158924 463666 158976
rect 464614 158924 464620 158976
rect 464672 158964 464678 158976
rect 471422 158964 471428 158976
rect 464672 158936 471428 158964
rect 464672 158924 464678 158936
rect 471422 158924 471428 158936
rect 471480 158924 471486 158976
rect 475562 158924 475568 158976
rect 475620 158964 475626 158976
rect 481634 158964 481640 158976
rect 475620 158936 481640 158964
rect 475620 158924 475626 158936
rect 481634 158924 481640 158936
rect 481692 158924 481698 158976
rect 102962 158856 102968 158908
rect 103020 158896 103026 158908
rect 125502 158896 125508 158908
rect 103020 158868 125508 158896
rect 103020 158856 103026 158868
rect 125502 158856 125508 158868
rect 125560 158856 125566 158908
rect 126238 158856 126244 158908
rect 126296 158896 126302 158908
rect 129734 158896 129740 158908
rect 126296 158868 129740 158896
rect 126296 158856 126302 158868
rect 129734 158856 129740 158868
rect 129792 158856 129798 158908
rect 130746 158856 130752 158908
rect 130804 158896 130810 158908
rect 194594 158896 194600 158908
rect 130804 158868 194600 158896
rect 130804 158856 130810 158868
rect 194594 158856 194600 158868
rect 194652 158856 194658 158908
rect 194686 158856 194692 158908
rect 194744 158896 194750 158908
rect 203702 158896 203708 158908
rect 194744 158868 203708 158896
rect 194744 158856 194750 158868
rect 203702 158856 203708 158868
rect 203760 158856 203766 158908
rect 208118 158856 208124 158908
rect 208176 158896 208182 158908
rect 212442 158896 212448 158908
rect 208176 158868 212448 158896
rect 208176 158856 208182 158868
rect 212442 158856 212448 158868
rect 212500 158856 212506 158908
rect 230750 158896 230756 158908
rect 215266 158868 230756 158896
rect 109678 158788 109684 158840
rect 109736 158828 109742 158840
rect 129918 158828 129924 158840
rect 109736 158800 129924 158828
rect 109736 158788 109742 158800
rect 129918 158788 129924 158800
rect 129976 158788 129982 158840
rect 133230 158788 133236 158840
rect 133288 158828 133294 158840
rect 158714 158828 158720 158840
rect 133288 158800 158720 158828
rect 133288 158788 133294 158800
rect 158714 158788 158720 158800
rect 158772 158788 158778 158840
rect 163498 158788 163504 158840
rect 163556 158828 163562 158840
rect 195974 158828 195980 158840
rect 163556 158800 195980 158828
rect 163556 158788 163562 158800
rect 195974 158788 195980 158800
rect 196032 158788 196038 158840
rect 207290 158788 207296 158840
rect 207348 158828 207354 158840
rect 215266 158828 215294 158868
rect 230750 158856 230756 158868
rect 230808 158856 230814 158908
rect 241790 158856 241796 158908
rect 241848 158896 241854 158908
rect 303522 158896 303528 158908
rect 241848 158868 303528 158896
rect 241848 158856 241854 158868
rect 303522 158856 303528 158868
rect 303580 158856 303586 158908
rect 305638 158856 305644 158908
rect 305696 158896 305702 158908
rect 307386 158896 307392 158908
rect 305696 158868 307392 158896
rect 305696 158856 305702 158868
rect 307386 158856 307392 158868
rect 307444 158856 307450 158908
rect 310698 158856 310704 158908
rect 310756 158896 310762 158908
rect 312170 158896 312176 158908
rect 310756 158868 312176 158896
rect 310756 158856 310762 158868
rect 312170 158856 312176 158868
rect 312228 158856 312234 158908
rect 312354 158856 312360 158908
rect 312412 158896 312418 158908
rect 318886 158896 318892 158908
rect 312412 158868 318892 158896
rect 312412 158856 312418 158868
rect 318886 158856 318892 158868
rect 318944 158856 318950 158908
rect 320818 158856 320824 158908
rect 320876 158896 320882 158908
rect 320876 158868 357572 158896
rect 320876 158856 320882 158868
rect 207348 158800 215294 158828
rect 207348 158788 207354 158800
rect 217318 158788 217324 158840
rect 217376 158828 217382 158840
rect 220354 158828 220360 158840
rect 217376 158800 220360 158828
rect 217376 158788 217382 158800
rect 220354 158788 220360 158800
rect 220412 158788 220418 158840
rect 238386 158788 238392 158840
rect 238444 158828 238450 158840
rect 241606 158828 241612 158840
rect 238444 158800 241612 158828
rect 238444 158788 238450 158800
rect 241606 158788 241612 158800
rect 241664 158788 241670 158840
rect 261110 158788 261116 158840
rect 261168 158828 261174 158840
rect 317046 158828 317052 158840
rect 261168 158800 317052 158828
rect 261168 158788 261174 158800
rect 317046 158788 317052 158800
rect 317104 158788 317110 158840
rect 319162 158788 319168 158840
rect 319220 158828 319226 158840
rect 319220 158800 321600 158828
rect 319220 158788 319226 158800
rect 90358 158720 90364 158772
rect 90416 158760 90422 158772
rect 92566 158760 92572 158772
rect 90416 158732 92572 158760
rect 90416 158720 90422 158732
rect 92566 158720 92572 158732
rect 92624 158720 92630 158772
rect 92842 158720 92848 158772
rect 92900 158760 92906 158772
rect 114462 158760 114468 158772
rect 92900 158732 114468 158760
rect 92900 158720 92906 158732
rect 114462 158720 114468 158732
rect 114520 158720 114526 158772
rect 119798 158720 119804 158772
rect 119856 158760 119862 158772
rect 146570 158760 146576 158772
rect 119856 158732 146576 158760
rect 119856 158720 119862 158732
rect 146570 158720 146576 158732
rect 146628 158720 146634 158772
rect 146662 158720 146668 158772
rect 146720 158760 146726 158772
rect 176654 158760 176660 158772
rect 146720 158732 176660 158760
rect 146720 158720 146726 158732
rect 176654 158720 176660 158732
rect 176712 158720 176718 158772
rect 180334 158720 180340 158772
rect 180392 158760 180398 158772
rect 204898 158760 204904 158772
rect 180392 158732 204904 158760
rect 180392 158720 180398 158732
rect 204898 158720 204904 158732
rect 204956 158720 204962 158772
rect 210602 158720 210608 158772
rect 210660 158760 210666 158772
rect 215386 158760 215392 158772
rect 210660 158732 215392 158760
rect 210660 158720 210666 158732
rect 215386 158720 215392 158732
rect 215444 158720 215450 158772
rect 221550 158720 221556 158772
rect 221608 158760 221614 158772
rect 224402 158760 224408 158772
rect 221608 158732 224408 158760
rect 221608 158720 221614 158732
rect 224402 158720 224408 158732
rect 224460 158720 224466 158772
rect 240870 158720 240876 158772
rect 240928 158760 240934 158772
rect 243354 158760 243360 158772
rect 240928 158732 243360 158760
rect 240928 158720 240934 158732
rect 243354 158720 243360 158732
rect 243412 158720 243418 158772
rect 254394 158720 254400 158772
rect 254452 158760 254458 158772
rect 255406 158760 255412 158772
rect 254452 158732 255412 158760
rect 254452 158720 254458 158732
rect 255406 158720 255412 158732
rect 255464 158720 255470 158772
rect 258534 158720 258540 158772
rect 258592 158760 258598 158772
rect 260926 158760 260932 158772
rect 258592 158732 260932 158760
rect 258592 158720 258598 158732
rect 260926 158720 260932 158732
rect 260984 158720 260990 158772
rect 264422 158720 264428 158772
rect 264480 158760 264486 158772
rect 266354 158760 266360 158772
rect 264480 158732 266360 158760
rect 264480 158720 264486 158732
rect 266354 158720 266360 158732
rect 266412 158720 266418 158772
rect 267826 158720 267832 158772
rect 267884 158760 267890 158772
rect 320266 158760 320272 158772
rect 267884 158732 320272 158760
rect 267884 158720 267890 158732
rect 320266 158720 320272 158732
rect 320324 158720 320330 158772
rect 321572 158704 321600 158800
rect 321646 158788 321652 158840
rect 321704 158828 321710 158840
rect 357434 158828 357440 158840
rect 321704 158800 357440 158828
rect 321704 158788 321710 158800
rect 357434 158788 357440 158800
rect 357492 158788 357498 158840
rect 357544 158828 357572 158868
rect 361206 158856 361212 158908
rect 361264 158896 361270 158908
rect 376754 158896 376760 158908
rect 361264 158868 376760 158896
rect 361264 158856 361270 158868
rect 376754 158856 376760 158868
rect 376812 158856 376818 158908
rect 376938 158856 376944 158908
rect 376996 158896 377002 158908
rect 378226 158896 378232 158908
rect 376996 158868 378232 158896
rect 376996 158856 377002 158868
rect 378226 158856 378232 158868
rect 378284 158856 378290 158908
rect 386138 158896 386144 158908
rect 383626 158868 386144 158896
rect 362954 158828 362960 158840
rect 357544 158800 362960 158828
rect 362954 158788 362960 158800
rect 363012 158788 363018 158840
rect 367922 158788 367928 158840
rect 367980 158828 367986 158840
rect 383626 158828 383654 158868
rect 386138 158856 386144 158868
rect 386196 158856 386202 158908
rect 391474 158856 391480 158908
rect 391532 158896 391538 158908
rect 393682 158896 393688 158908
rect 391532 158868 393688 158896
rect 391532 158856 391538 158868
rect 393682 158856 393688 158868
rect 393740 158856 393746 158908
rect 412542 158856 412548 158908
rect 412600 158896 412606 158908
rect 412910 158896 412916 158908
rect 412600 158868 412916 158896
rect 412600 158856 412606 158868
rect 412910 158856 412916 158868
rect 412968 158856 412974 158908
rect 454586 158856 454592 158908
rect 454644 158896 454650 158908
rect 462222 158896 462228 158908
rect 454644 158868 462228 158896
rect 454644 158856 454650 158868
rect 462222 158856 462228 158868
rect 462280 158856 462286 158908
rect 466362 158856 466368 158908
rect 466420 158896 466426 158908
rect 472434 158896 472440 158908
rect 466420 158868 472440 158896
rect 466420 158856 466426 158868
rect 472434 158856 472440 158868
rect 472492 158856 472498 158908
rect 476390 158856 476396 158908
rect 476448 158896 476454 158908
rect 482646 158896 482652 158908
rect 476448 158868 482652 158896
rect 476448 158856 476454 158868
rect 482646 158856 482652 158868
rect 482704 158856 482710 158908
rect 508314 158856 508320 158908
rect 508372 158896 508378 158908
rect 510062 158896 510068 158908
rect 508372 158868 510068 158896
rect 508372 158856 508378 158868
rect 510062 158856 510068 158868
rect 510120 158856 510126 158908
rect 386230 158828 386236 158840
rect 367980 158800 373994 158828
rect 367980 158788 367986 158800
rect 327534 158720 327540 158772
rect 327592 158760 327598 158772
rect 367186 158760 367192 158772
rect 327592 158732 367192 158760
rect 327592 158720 327598 158732
rect 367186 158720 367192 158732
rect 367244 158720 367250 158772
rect 373966 158760 373994 158800
rect 376956 158800 383654 158828
rect 384684 158800 386236 158828
rect 373966 158732 376800 158760
rect 81066 158652 81072 158704
rect 81124 158692 81130 158704
rect 180886 158692 180892 158704
rect 81124 158664 180892 158692
rect 81124 158652 81130 158664
rect 180886 158652 180892 158664
rect 180944 158652 180950 158704
rect 181990 158652 181996 158704
rect 182048 158692 182054 158704
rect 256786 158692 256792 158704
rect 182048 158664 256792 158692
rect 182048 158652 182054 158664
rect 256786 158652 256792 158664
rect 256844 158652 256850 158704
rect 321554 158652 321560 158704
rect 321612 158652 321618 158704
rect 376772 158692 376800 158732
rect 376956 158692 376984 158800
rect 384684 158760 384712 158800
rect 386230 158788 386236 158800
rect 386288 158788 386294 158840
rect 388070 158788 388076 158840
rect 388128 158828 388134 158840
rect 390370 158828 390376 158840
rect 388128 158800 390376 158828
rect 388128 158788 388134 158800
rect 390370 158788 390376 158800
rect 390428 158788 390434 158840
rect 409138 158788 409144 158840
rect 409196 158828 409202 158840
rect 410794 158828 410800 158840
rect 409196 158800 410800 158828
rect 409196 158788 409202 158800
rect 410794 158788 410800 158800
rect 410852 158788 410858 158840
rect 416682 158788 416688 158840
rect 416740 158828 416746 158840
rect 419534 158828 419540 158840
rect 416740 158800 419540 158828
rect 416740 158788 416746 158800
rect 419534 158788 419540 158800
rect 419592 158788 419598 158840
rect 452838 158788 452844 158840
rect 452896 158828 452902 158840
rect 459646 158828 459652 158840
rect 452896 158800 459652 158828
rect 452896 158788 452902 158800
rect 459646 158788 459652 158800
rect 459704 158788 459710 158840
rect 463786 158788 463792 158840
rect 463844 158828 463850 158840
rect 471330 158828 471336 158840
rect 463844 158800 471336 158828
rect 463844 158788 463850 158800
rect 471330 158788 471336 158800
rect 471388 158788 471394 158840
rect 474734 158788 474740 158840
rect 474792 158828 474798 158840
rect 480254 158828 480260 158840
rect 474792 158800 480260 158828
rect 474792 158788 474798 158800
rect 480254 158788 480260 158800
rect 480312 158788 480318 158840
rect 482278 158788 482284 158840
rect 482336 158828 482342 158840
rect 487246 158828 487252 158840
rect 482336 158800 487252 158828
rect 482336 158788 482342 158800
rect 487246 158788 487252 158800
rect 487304 158788 487310 158840
rect 506382 158788 506388 158840
rect 506440 158828 506446 158840
rect 507578 158828 507584 158840
rect 506440 158800 507584 158828
rect 506440 158788 506446 158800
rect 507578 158788 507584 158800
rect 507636 158788 507642 158840
rect 376772 158664 376984 158692
rect 377048 158732 384712 158760
rect 67634 158584 67640 158636
rect 67692 158624 67698 158636
rect 170306 158624 170312 158636
rect 67692 158596 170312 158624
rect 67692 158584 67698 158596
rect 170306 158584 170312 158596
rect 170364 158584 170370 158636
rect 171962 158584 171968 158636
rect 172020 158624 172026 158636
rect 250070 158624 250076 158636
rect 172020 158596 250076 158624
rect 172020 158584 172026 158596
rect 250070 158584 250076 158596
rect 250128 158584 250134 158636
rect 376754 158584 376760 158636
rect 376812 158624 376818 158636
rect 377048 158624 377076 158732
rect 384758 158720 384764 158772
rect 384816 158760 384822 158772
rect 389174 158760 389180 158772
rect 384816 158732 389180 158760
rect 384816 158720 384822 158732
rect 389174 158720 389180 158732
rect 389232 158720 389238 158772
rect 405734 158720 405740 158772
rect 405792 158760 405798 158772
rect 409230 158760 409236 158772
rect 405792 158732 409236 158760
rect 405792 158720 405798 158732
rect 409230 158720 409236 158732
rect 409288 158720 409294 158772
rect 413370 158720 413376 158772
rect 413428 158760 413434 158772
rect 419626 158760 419632 158772
rect 413428 158732 419632 158760
rect 413428 158720 413434 158732
rect 419626 158720 419632 158732
rect 419684 158720 419690 158772
rect 453758 158720 453764 158772
rect 453816 158760 453822 158772
rect 459554 158760 459560 158772
rect 453816 158732 459560 158760
rect 453816 158720 453822 158732
rect 459554 158720 459560 158732
rect 459612 158720 459618 158772
rect 462958 158720 462964 158772
rect 463016 158760 463022 158772
rect 469214 158760 469220 158772
rect 463016 158732 469220 158760
rect 463016 158720 463022 158732
rect 469214 158720 469220 158732
rect 469272 158720 469278 158772
rect 473078 158720 473084 158772
rect 473136 158760 473142 158772
rect 478966 158760 478972 158772
rect 473136 158732 478972 158760
rect 473136 158720 473142 158732
rect 478966 158720 478972 158732
rect 479024 158720 479030 158772
rect 481450 158720 481456 158772
rect 481508 158760 481514 158772
rect 486510 158760 486516 158772
rect 481508 158732 486516 158760
rect 481508 158720 481514 158732
rect 486510 158720 486516 158732
rect 486568 158720 486574 158772
rect 505278 158720 505284 158772
rect 505336 158760 505342 158772
rect 506750 158760 506756 158772
rect 505336 158732 506756 158760
rect 505336 158720 505342 158732
rect 506750 158720 506756 158732
rect 506808 158720 506814 158772
rect 507026 158720 507032 158772
rect 507084 158760 507090 158772
rect 508406 158760 508412 158772
rect 507084 158732 508412 158760
rect 507084 158720 507090 158732
rect 508406 158720 508412 158732
rect 508464 158720 508470 158772
rect 509418 158720 509424 158772
rect 509476 158760 509482 158772
rect 511718 158760 511724 158772
rect 509476 158732 511724 158760
rect 509476 158720 509482 158732
rect 511718 158720 511724 158732
rect 511776 158720 511782 158772
rect 514938 158720 514944 158772
rect 514996 158760 515002 158772
rect 518526 158760 518532 158772
rect 514996 158732 518532 158760
rect 514996 158720 515002 158732
rect 518526 158720 518532 158732
rect 518584 158720 518590 158772
rect 376812 158596 377076 158624
rect 376812 158584 376818 158596
rect 74350 158516 74356 158568
rect 74408 158556 74414 158568
rect 175182 158556 175188 158568
rect 74408 158528 175188 158556
rect 74408 158516 74414 158528
rect 175182 158516 175188 158528
rect 175240 158516 175246 158568
rect 175274 158516 175280 158568
rect 175332 158556 175338 158568
rect 252738 158556 252744 158568
rect 175332 158528 252744 158556
rect 175332 158516 175338 158528
rect 252738 158516 252744 158528
rect 252796 158516 252802 158568
rect 71038 158448 71044 158500
rect 71096 158488 71102 158500
rect 71096 158460 170076 158488
rect 71096 158448 71102 158460
rect 64230 158380 64236 158432
rect 64288 158420 64294 158432
rect 167546 158420 167552 158432
rect 64288 158392 167552 158420
rect 64288 158380 64294 158392
rect 167546 158380 167552 158392
rect 167604 158380 167610 158432
rect 168558 158380 168564 158432
rect 168616 158420 168622 158432
rect 169662 158420 169668 158432
rect 168616 158392 169668 158420
rect 168616 158380 168622 158392
rect 169662 158380 169668 158392
rect 169720 158380 169726 158432
rect 170048 158420 170076 158460
rect 171778 158448 171784 158500
rect 171836 158488 171842 158500
rect 178034 158488 178040 158500
rect 171836 158460 178040 158488
rect 171836 158448 171842 158460
rect 178034 158448 178040 158460
rect 178092 158448 178098 158500
rect 178678 158448 178684 158500
rect 178736 158488 178742 158500
rect 255590 158488 255596 158500
rect 178736 158460 255596 158488
rect 178736 158448 178742 158460
rect 255590 158448 255596 158460
rect 255648 158448 255654 158500
rect 173066 158420 173072 158432
rect 170048 158392 173072 158420
rect 173066 158380 173072 158392
rect 173124 158380 173130 158432
rect 173158 158380 173164 158432
rect 173216 158420 173222 158432
rect 247126 158420 247132 158432
rect 173216 158392 247132 158420
rect 173216 158380 173222 158392
rect 247126 158380 247132 158392
rect 247184 158380 247190 158432
rect 60918 158312 60924 158364
rect 60976 158352 60982 158364
rect 164326 158352 164332 158364
rect 60976 158324 164332 158352
rect 60976 158312 60982 158324
rect 164326 158312 164332 158324
rect 164384 158312 164390 158364
rect 165246 158312 165252 158364
rect 165304 158352 165310 158364
rect 245010 158352 245016 158364
rect 165304 158324 245016 158352
rect 165304 158312 165310 158324
rect 245010 158312 245016 158324
rect 245068 158312 245074 158364
rect 54202 158244 54208 158296
rect 54260 158284 54266 158296
rect 160278 158284 160284 158296
rect 54260 158256 160284 158284
rect 54260 158244 54266 158256
rect 160278 158244 160284 158256
rect 160336 158244 160342 158296
rect 161842 158244 161848 158296
rect 161900 158284 161906 158296
rect 242066 158284 242072 158296
rect 161900 158256 242072 158284
rect 161900 158244 161906 158256
rect 242066 158244 242072 158256
rect 242124 158244 242130 158296
rect 50798 158176 50804 158228
rect 50856 158216 50862 158228
rect 157702 158216 157708 158228
rect 50856 158188 157708 158216
rect 50856 158176 50862 158188
rect 157702 158176 157708 158188
rect 157760 158176 157766 158228
rect 158438 158176 158444 158228
rect 158496 158216 158502 158228
rect 238938 158216 238944 158228
rect 158496 158188 238944 158216
rect 158496 158176 158502 158188
rect 238938 158176 238944 158188
rect 238996 158176 239002 158228
rect 256878 158176 256884 158228
rect 256936 158216 256942 158228
rect 315022 158216 315028 158228
rect 256936 158188 315028 158216
rect 256936 158176 256942 158188
rect 315022 158176 315028 158188
rect 315080 158176 315086 158228
rect 47486 158108 47492 158160
rect 47544 158148 47550 158160
rect 155034 158148 155040 158160
rect 47544 158120 155040 158148
rect 47544 158108 47550 158120
rect 155034 158108 155040 158120
rect 155092 158108 155098 158160
rect 155126 158108 155132 158160
rect 155184 158148 155190 158160
rect 237374 158148 237380 158160
rect 155184 158120 237380 158148
rect 155184 158108 155190 158120
rect 237374 158108 237380 158120
rect 237432 158108 237438 158160
rect 246758 158108 246764 158160
rect 246816 158148 246822 158160
rect 306926 158148 306932 158160
rect 246816 158120 306932 158148
rect 246816 158108 246822 158120
rect 306926 158108 306932 158120
rect 306984 158108 306990 158160
rect 37366 158040 37372 158092
rect 37424 158080 37430 158092
rect 146386 158080 146392 158092
rect 37424 158052 146392 158080
rect 37424 158040 37430 158052
rect 146386 158040 146392 158052
rect 146444 158040 146450 158092
rect 148410 158040 148416 158092
rect 148468 158080 148474 158092
rect 231946 158080 231952 158092
rect 148468 158052 231952 158080
rect 148468 158040 148474 158052
rect 231946 158040 231952 158052
rect 232004 158040 232010 158092
rect 243446 158040 243452 158092
rect 243504 158080 243510 158092
rect 304718 158080 304724 158092
rect 243504 158052 304724 158080
rect 243504 158040 243510 158052
rect 304718 158040 304724 158052
rect 304776 158040 304782 158092
rect 382 157972 388 158024
rect 440 158012 446 158024
rect 118878 158012 118884 158024
rect 440 157984 118884 158012
rect 440 157972 446 157984
rect 118878 157972 118884 157984
rect 118936 157972 118942 158024
rect 131758 157972 131764 158024
rect 131816 158012 131822 158024
rect 219342 158012 219348 158024
rect 131816 157984 219348 158012
rect 131816 157972 131822 157984
rect 219342 157972 219348 157984
rect 219400 157972 219406 158024
rect 236730 157972 236736 158024
rect 236788 158012 236794 158024
rect 299658 158012 299664 158024
rect 236788 157984 299664 158012
rect 236788 157972 236794 157984
rect 299658 157972 299664 157984
rect 299716 157972 299722 158024
rect 77754 157904 77760 157956
rect 77812 157944 77818 157956
rect 171778 157944 171784 157956
rect 77812 157916 171784 157944
rect 77812 157904 77818 157916
rect 171778 157904 171784 157916
rect 171836 157904 171842 157956
rect 171870 157904 171876 157956
rect 171928 157944 171934 157956
rect 182266 157944 182272 157956
rect 171928 157916 182272 157944
rect 171928 157904 171934 157916
rect 182266 157904 182272 157916
rect 182324 157904 182330 157956
rect 185302 157944 185308 157956
rect 185228 157916 185308 157944
rect 87782 157836 87788 157888
rect 87840 157876 87846 157888
rect 185118 157876 185124 157888
rect 87840 157848 171916 157876
rect 87840 157836 87846 157848
rect 84470 157768 84476 157820
rect 84528 157808 84534 157820
rect 171778 157808 171784 157820
rect 84528 157780 171784 157808
rect 84528 157768 84534 157780
rect 171778 157768 171784 157780
rect 171836 157768 171842 157820
rect 171888 157808 171916 157848
rect 173866 157848 185124 157876
rect 173866 157808 173894 157848
rect 185118 157836 185124 157848
rect 185176 157836 185182 157888
rect 171888 157780 173894 157808
rect 179414 157768 179420 157820
rect 179472 157808 179478 157820
rect 185228 157808 185256 157916
rect 185302 157904 185308 157916
rect 185360 157904 185366 157956
rect 185394 157904 185400 157956
rect 185452 157944 185458 157956
rect 260466 157944 260472 157956
rect 185452 157916 260472 157944
rect 185452 157904 185458 157916
rect 260466 157904 260472 157916
rect 260524 157904 260530 157956
rect 188798 157836 188804 157888
rect 188856 157876 188862 157888
rect 263042 157876 263048 157888
rect 188856 157848 263048 157876
rect 188856 157836 188862 157848
rect 263042 157836 263048 157848
rect 263100 157836 263106 157888
rect 190638 157808 190644 157820
rect 179472 157780 185256 157808
rect 185504 157780 190644 157808
rect 179472 157768 179478 157780
rect 91186 157700 91192 157752
rect 91244 157740 91250 157752
rect 185302 157740 185308 157752
rect 91244 157712 185308 157740
rect 91244 157700 91250 157712
rect 185302 157700 185308 157712
rect 185360 157700 185366 157752
rect 94590 157632 94596 157684
rect 94648 157672 94654 157684
rect 185504 157672 185532 157780
rect 190638 157768 190644 157780
rect 190696 157768 190702 157820
rect 195514 157768 195520 157820
rect 195572 157808 195578 157820
rect 267734 157808 267740 157820
rect 195572 157780 267740 157808
rect 195572 157768 195578 157780
rect 267734 157768 267740 157780
rect 267792 157768 267798 157820
rect 185670 157700 185676 157752
rect 185728 157740 185734 157752
rect 188522 157740 188528 157752
rect 185728 157712 188528 157740
rect 185728 157700 185734 157712
rect 188522 157700 188528 157712
rect 188580 157700 188586 157752
rect 190454 157700 190460 157752
rect 190512 157740 190518 157752
rect 263686 157740 263692 157752
rect 190512 157712 263692 157740
rect 190512 157700 190518 157712
rect 263686 157700 263692 157712
rect 263744 157700 263750 157752
rect 94648 157644 185532 157672
rect 94648 157632 94654 157644
rect 185578 157632 185584 157684
rect 185636 157672 185642 157684
rect 236086 157672 236092 157684
rect 185636 157644 236092 157672
rect 185636 157632 185642 157644
rect 236086 157632 236092 157644
rect 236144 157632 236150 157684
rect 97902 157564 97908 157616
rect 97960 157604 97966 157616
rect 193214 157604 193220 157616
rect 97960 157576 193220 157604
rect 97960 157564 97966 157576
rect 193214 157564 193220 157576
rect 193272 157564 193278 157616
rect 197354 157564 197360 157616
rect 197412 157604 197418 157616
rect 251450 157604 251456 157616
rect 197412 157576 251456 157604
rect 197412 157564 197418 157576
rect 251450 157564 251456 157576
rect 251508 157564 251514 157616
rect 111334 157496 111340 157548
rect 111392 157536 111398 157548
rect 203426 157536 203432 157548
rect 111392 157508 203432 157536
rect 111392 157496 111398 157508
rect 203426 157496 203432 157508
rect 203484 157496 203490 157548
rect 204898 157496 204904 157548
rect 204956 157536 204962 157548
rect 255866 157536 255872 157548
rect 204956 157508 255872 157536
rect 204956 157496 204962 157508
rect 255866 157496 255872 157508
rect 255924 157496 255930 157548
rect 114738 157428 114744 157480
rect 114796 157468 114802 157480
rect 206554 157468 206560 157480
rect 114796 157440 206560 157468
rect 114796 157428 114802 157440
rect 206554 157428 206560 157440
rect 206612 157428 206618 157480
rect 214558 157428 214564 157480
rect 214616 157468 214622 157480
rect 214616 157440 222194 157468
rect 214616 157428 214622 157440
rect 141694 157360 141700 157412
rect 141752 157400 141758 157412
rect 222166 157400 222194 157440
rect 227070 157400 227076 157412
rect 141752 157372 212534 157400
rect 222166 157372 227076 157400
rect 141752 157360 141758 157372
rect 49142 157292 49148 157344
rect 49200 157332 49206 157344
rect 156414 157332 156420 157344
rect 49200 157304 156420 157332
rect 49200 157292 49206 157304
rect 156414 157292 156420 157304
rect 156472 157292 156478 157344
rect 158714 157292 158720 157344
rect 158772 157332 158778 157344
rect 210510 157332 210516 157344
rect 158772 157304 210516 157332
rect 158772 157292 158778 157304
rect 210510 157292 210516 157304
rect 210568 157292 210574 157344
rect 212506 157332 212534 157372
rect 227070 157360 227076 157372
rect 227128 157360 227134 157412
rect 214374 157332 214380 157344
rect 212506 157304 214380 157332
rect 214374 157292 214380 157304
rect 214432 157292 214438 157344
rect 221182 157292 221188 157344
rect 221240 157332 221246 157344
rect 221240 157304 273254 157332
rect 221240 157292 221246 157304
rect 45738 157224 45744 157276
rect 45796 157264 45802 157276
rect 153746 157264 153752 157276
rect 45796 157236 153752 157264
rect 45796 157224 45802 157236
rect 153746 157224 153752 157236
rect 153804 157224 153810 157276
rect 163774 157224 163780 157276
rect 163832 157264 163838 157276
rect 166442 157264 166448 157276
rect 163832 157236 166448 157264
rect 163832 157224 163838 157236
rect 166442 157224 166448 157236
rect 166500 157224 166506 157276
rect 192110 157224 192116 157276
rect 192168 157264 192174 157276
rect 265158 157264 265164 157276
rect 192168 157236 265164 157264
rect 192168 157224 192174 157236
rect 265158 157224 265164 157236
rect 265216 157224 265222 157276
rect 42426 157156 42432 157208
rect 42484 157196 42490 157208
rect 151262 157196 151268 157208
rect 42484 157168 151268 157196
rect 42484 157156 42490 157168
rect 151262 157156 151268 157168
rect 151320 157156 151326 157208
rect 156506 157156 156512 157208
rect 156564 157196 156570 157208
rect 159082 157196 159088 157208
rect 156564 157168 159088 157196
rect 156564 157156 156570 157168
rect 159082 157156 159088 157168
rect 159140 157156 159146 157208
rect 160094 157156 160100 157208
rect 160152 157196 160158 157208
rect 166166 157196 166172 157208
rect 160152 157168 166172 157196
rect 160152 157156 160158 157168
rect 166166 157156 166172 157168
rect 166224 157156 166230 157208
rect 166258 157156 166264 157208
rect 166316 157196 166322 157208
rect 171134 157196 171140 157208
rect 166316 157168 171140 157196
rect 166316 157156 166322 157168
rect 171134 157156 171140 157168
rect 171192 157156 171198 157208
rect 177022 157156 177028 157208
rect 177080 157196 177086 157208
rect 254026 157196 254032 157208
rect 177080 157168 254032 157196
rect 177080 157156 177086 157168
rect 254026 157156 254032 157168
rect 254084 157156 254090 157208
rect 273226 157196 273254 157304
rect 283834 157224 283840 157276
rect 283892 157264 283898 157276
rect 335538 157264 335544 157276
rect 283892 157236 335544 157264
rect 283892 157224 283898 157236
rect 335538 157224 335544 157236
rect 335596 157224 335602 157276
rect 281626 157196 281632 157208
rect 273226 157168 281632 157196
rect 281626 157156 281632 157168
rect 281684 157156 281690 157208
rect 300670 157156 300676 157208
rect 300728 157196 300734 157208
rect 348050 157196 348056 157208
rect 300728 157168 348056 157196
rect 300728 157156 300734 157168
rect 348050 157156 348056 157168
rect 348108 157156 348114 157208
rect 39022 157088 39028 157140
rect 39080 157128 39086 157140
rect 147674 157128 147680 157140
rect 39080 157100 147680 157128
rect 39080 157088 39086 157100
rect 147674 157088 147680 157100
rect 147732 157088 147738 157140
rect 150066 157088 150072 157140
rect 150124 157128 150130 157140
rect 233510 157128 233516 157140
rect 150124 157100 233516 157128
rect 150124 157088 150130 157100
rect 233510 157088 233516 157100
rect 233568 157088 233574 157140
rect 287146 157088 287152 157140
rect 287204 157128 287210 157140
rect 338114 157128 338120 157140
rect 287204 157100 338120 157128
rect 287204 157088 287210 157100
rect 338114 157088 338120 157100
rect 338172 157088 338178 157140
rect 35710 157020 35716 157072
rect 35768 157060 35774 157072
rect 146202 157060 146208 157072
rect 35768 157032 146208 157060
rect 35768 157020 35774 157032
rect 146202 157020 146208 157032
rect 146260 157020 146266 157072
rect 151722 157020 151728 157072
rect 151780 157060 151786 157072
rect 234798 157060 234804 157072
rect 151780 157032 234804 157060
rect 151780 157020 151786 157032
rect 234798 157020 234804 157032
rect 234856 157020 234862 157072
rect 280430 157020 280436 157072
rect 280488 157060 280494 157072
rect 333054 157060 333060 157072
rect 280488 157032 333060 157060
rect 280488 157020 280494 157032
rect 333054 157020 333060 157032
rect 333112 157020 333118 157072
rect 24762 156952 24768 157004
rect 24820 156992 24826 157004
rect 137370 156992 137376 157004
rect 24820 156964 137376 156992
rect 24820 156952 24826 156964
rect 137370 156952 137376 156964
rect 137428 156952 137434 157004
rect 138290 156952 138296 157004
rect 138348 156992 138354 157004
rect 224126 156992 224132 157004
rect 138348 156964 224132 156992
rect 138348 156952 138354 156964
rect 224126 156952 224132 156964
rect 224184 156952 224190 157004
rect 273714 156952 273720 157004
rect 273772 156992 273778 157004
rect 327902 156992 327908 157004
rect 273772 156964 327908 156992
rect 273772 156952 273778 156964
rect 327902 156952 327908 156964
rect 327960 156952 327966 157004
rect 21358 156884 21364 156936
rect 21416 156924 21422 156936
rect 135254 156924 135260 156936
rect 21416 156896 135260 156924
rect 21416 156884 21422 156896
rect 135254 156884 135260 156896
rect 135312 156884 135318 156936
rect 135806 156884 135812 156936
rect 135864 156924 135870 156936
rect 222562 156924 222568 156936
rect 135864 156896 222568 156924
rect 135864 156884 135870 156896
rect 222562 156884 222568 156896
rect 222620 156884 222626 156936
rect 224954 156884 224960 156936
rect 225012 156924 225018 156936
rect 272058 156924 272064 156936
rect 225012 156896 272064 156924
rect 225012 156884 225018 156896
rect 272058 156884 272064 156896
rect 272116 156884 272122 156936
rect 277118 156884 277124 156936
rect 277176 156924 277182 156936
rect 330478 156924 330484 156936
rect 277176 156896 330484 156924
rect 277176 156884 277182 156896
rect 330478 156884 330484 156896
rect 330536 156884 330542 156936
rect 18046 156816 18052 156868
rect 18104 156856 18110 156868
rect 132494 156856 132500 156868
rect 18104 156828 132500 156856
rect 18104 156816 18110 156828
rect 132494 156816 132500 156828
rect 132552 156816 132558 156868
rect 134886 156816 134892 156868
rect 134944 156856 134950 156868
rect 210418 156856 210424 156868
rect 134944 156828 210424 156856
rect 134944 156816 134950 156828
rect 210418 156816 210424 156828
rect 210476 156816 210482 156868
rect 210602 156816 210608 156868
rect 210660 156856 210666 156868
rect 214190 156856 214196 156868
rect 210660 156828 214196 156856
rect 210660 156816 210666 156828
rect 214190 156816 214196 156828
rect 214248 156816 214254 156868
rect 219710 156816 219716 156868
rect 219768 156856 219774 156868
rect 219768 156828 225276 156856
rect 219768 156816 219774 156828
rect 14642 156748 14648 156800
rect 14700 156788 14706 156800
rect 130102 156788 130108 156800
rect 14700 156760 130108 156788
rect 14700 156748 14706 156760
rect 130102 156748 130108 156760
rect 130160 156748 130166 156800
rect 139118 156748 139124 156800
rect 139176 156788 139182 156800
rect 225138 156788 225144 156800
rect 139176 156760 225144 156788
rect 139176 156748 139182 156760
rect 225138 156748 225144 156760
rect 225196 156748 225202 156800
rect 225248 156788 225276 156828
rect 226610 156816 226616 156868
rect 226668 156856 226674 156868
rect 291930 156856 291936 156868
rect 226668 156828 291936 156856
rect 226668 156816 226674 156828
rect 291930 156816 291936 156828
rect 291988 156816 291994 156868
rect 293862 156816 293868 156868
rect 293920 156856 293926 156868
rect 342530 156856 342536 156868
rect 293920 156828 342536 156856
rect 293920 156816 293926 156828
rect 342530 156816 342536 156828
rect 342588 156816 342594 156868
rect 228358 156788 228364 156800
rect 225248 156760 228364 156788
rect 228358 156748 228364 156760
rect 228416 156748 228422 156800
rect 230014 156748 230020 156800
rect 230072 156788 230078 156800
rect 294046 156788 294052 156800
rect 230072 156760 294052 156788
rect 230072 156748 230078 156760
rect 294046 156748 294052 156760
rect 294104 156748 294110 156800
rect 297266 156748 297272 156800
rect 297324 156788 297330 156800
rect 345106 156788 345112 156800
rect 297324 156760 345112 156788
rect 297324 156748 297330 156760
rect 345106 156748 345112 156760
rect 345164 156748 345170 156800
rect 11238 156680 11244 156732
rect 11296 156720 11302 156732
rect 127526 156720 127532 156732
rect 11296 156692 127532 156720
rect 11296 156680 11302 156692
rect 127526 156680 127532 156692
rect 127584 156680 127590 156732
rect 128170 156680 128176 156732
rect 128228 156720 128234 156732
rect 216766 156720 216772 156732
rect 128228 156692 216772 156720
rect 128228 156680 128234 156692
rect 216766 156680 216772 156692
rect 216824 156680 216830 156732
rect 223206 156680 223212 156732
rect 223264 156720 223270 156732
rect 289354 156720 289360 156732
rect 223264 156692 289360 156720
rect 223264 156680 223270 156692
rect 289354 156680 289360 156692
rect 289412 156680 289418 156732
rect 290550 156680 290556 156732
rect 290608 156720 290614 156732
rect 340046 156720 340052 156732
rect 290608 156692 340052 156720
rect 290608 156680 290614 156692
rect 340046 156680 340052 156692
rect 340104 156680 340110 156732
rect 2038 156612 2044 156664
rect 2096 156652 2102 156664
rect 120442 156652 120448 156664
rect 2096 156624 120448 156652
rect 2096 156612 2102 156624
rect 120442 156612 120448 156624
rect 120500 156612 120506 156664
rect 124858 156612 124864 156664
rect 124916 156652 124922 156664
rect 209774 156652 209780 156664
rect 124916 156624 209780 156652
rect 124916 156612 124922 156624
rect 209774 156612 209780 156624
rect 209832 156612 209838 156664
rect 209958 156612 209964 156664
rect 210016 156652 210022 156664
rect 211614 156652 211620 156664
rect 210016 156624 211620 156652
rect 210016 156612 210022 156624
rect 211614 156612 211620 156624
rect 211672 156612 211678 156664
rect 216490 156612 216496 156664
rect 216548 156652 216554 156664
rect 283098 156652 283104 156664
rect 216548 156624 283104 156652
rect 216548 156612 216554 156624
rect 283098 156612 283104 156624
rect 283156 156612 283162 156664
rect 498286 156612 498292 156664
rect 498344 156652 498350 156664
rect 499298 156652 499304 156664
rect 498344 156624 499304 156652
rect 498344 156612 498350 156624
rect 499298 156612 499304 156624
rect 499356 156612 499362 156664
rect 502334 156612 502340 156664
rect 502392 156652 502398 156664
rect 503346 156652 503352 156664
rect 502392 156624 503352 156652
rect 502392 156612 502398 156624
rect 503346 156612 503352 156624
rect 503404 156612 503410 156664
rect 52454 156544 52460 156596
rect 52512 156584 52518 156596
rect 158990 156584 158996 156596
rect 52512 156556 158996 156584
rect 52512 156544 52518 156556
rect 158990 156544 158996 156556
rect 159048 156544 159054 156596
rect 159082 156544 159088 156596
rect 159140 156584 159146 156596
rect 200758 156584 200764 156596
rect 159140 156556 200764 156584
rect 159140 156544 159146 156556
rect 200758 156544 200764 156556
rect 200816 156544 200822 156596
rect 200942 156544 200948 156596
rect 201000 156584 201006 156596
rect 270494 156584 270500 156596
rect 201000 156556 270500 156584
rect 201000 156544 201006 156556
rect 270494 156544 270500 156556
rect 270552 156544 270558 156596
rect 59262 156476 59268 156528
rect 59320 156516 59326 156528
rect 164142 156516 164148 156528
rect 59320 156488 164148 156516
rect 59320 156476 59326 156488
rect 164142 156476 164148 156488
rect 164200 156476 164206 156528
rect 166166 156476 166172 156528
rect 166224 156516 166230 156528
rect 166224 156488 166396 156516
rect 166224 156476 166230 156488
rect 69290 156408 69296 156460
rect 69348 156448 69354 156460
rect 166258 156448 166264 156460
rect 69348 156420 166264 156448
rect 69348 156408 69354 156420
rect 166258 156408 166264 156420
rect 166316 156408 166322 156460
rect 166368 156448 166396 156488
rect 166442 156476 166448 156528
rect 166500 156516 166506 156528
rect 225046 156516 225052 156528
rect 166500 156488 225052 156516
rect 166500 156476 166506 156488
rect 225046 156476 225052 156488
rect 225104 156476 225110 156528
rect 219710 156448 219716 156460
rect 166368 156420 219716 156448
rect 219710 156408 219716 156420
rect 219768 156408 219774 156460
rect 219802 156408 219808 156460
rect 219860 156448 219866 156460
rect 221366 156448 221372 156460
rect 219860 156420 221372 156448
rect 219860 156408 219866 156420
rect 221366 156408 221372 156420
rect 221424 156408 221430 156460
rect 82814 156340 82820 156392
rect 82872 156380 82878 156392
rect 182082 156380 182088 156392
rect 82872 156352 182088 156380
rect 82872 156340 82878 156352
rect 182082 156340 182088 156352
rect 182140 156340 182146 156392
rect 198826 156340 198832 156392
rect 198884 156380 198890 156392
rect 200942 156380 200948 156392
rect 198884 156352 200948 156380
rect 198884 156340 198890 156352
rect 200942 156340 200948 156352
rect 201000 156340 201006 156392
rect 209866 156340 209872 156392
rect 209924 156380 209930 156392
rect 279050 156380 279056 156392
rect 209924 156352 279056 156380
rect 209924 156340 209930 156352
rect 279050 156340 279056 156352
rect 279108 156340 279114 156392
rect 99558 156272 99564 156324
rect 99616 156312 99622 156324
rect 194962 156312 194968 156324
rect 99616 156284 194968 156312
rect 99616 156272 99622 156284
rect 194962 156272 194968 156284
rect 195020 156272 195026 156324
rect 195974 156272 195980 156324
rect 196032 156312 196038 156324
rect 196986 156312 196992 156324
rect 196032 156284 196992 156312
rect 196032 156272 196038 156284
rect 196986 156272 196992 156284
rect 197044 156272 197050 156324
rect 200758 156272 200764 156324
rect 200816 156312 200822 156324
rect 200816 156284 210372 156312
rect 200816 156272 200822 156284
rect 101306 156204 101312 156256
rect 101364 156244 101370 156256
rect 196250 156244 196256 156256
rect 101364 156216 196256 156244
rect 101364 156204 101370 156216
rect 196250 156204 196256 156216
rect 196308 156204 196314 156256
rect 197998 156204 198004 156256
rect 198056 156244 198062 156256
rect 209958 156244 209964 156256
rect 198056 156216 209964 156244
rect 198056 156204 198062 156216
rect 209958 156204 209964 156216
rect 210016 156204 210022 156256
rect 108022 156136 108028 156188
rect 108080 156176 108086 156188
rect 200666 156176 200672 156188
rect 108080 156148 200672 156176
rect 108080 156136 108086 156148
rect 200666 156136 200672 156148
rect 200724 156136 200730 156188
rect 209130 156176 209136 156188
rect 201236 156148 209136 156176
rect 118142 156068 118148 156120
rect 118200 156108 118206 156120
rect 201236 156108 201264 156148
rect 209130 156136 209136 156148
rect 209188 156136 209194 156188
rect 210344 156176 210372 156284
rect 210418 156272 210424 156324
rect 210476 156312 210482 156324
rect 219802 156312 219808 156324
rect 210476 156284 219808 156312
rect 210476 156272 210482 156284
rect 219802 156272 219808 156284
rect 219860 156272 219866 156324
rect 219894 156272 219900 156324
rect 219952 156312 219958 156324
rect 286226 156312 286232 156324
rect 219952 156284 286232 156312
rect 219952 156272 219958 156284
rect 286226 156272 286232 156284
rect 286284 156272 286290 156324
rect 210510 156204 210516 156256
rect 210568 156244 210574 156256
rect 219986 156244 219992 156256
rect 210568 156216 219992 156244
rect 210568 156204 210574 156216
rect 219986 156204 219992 156216
rect 220044 156204 220050 156256
rect 266906 156244 266912 156256
rect 229066 156216 266912 156244
rect 215478 156176 215484 156188
rect 210344 156148 215484 156176
rect 215478 156136 215484 156148
rect 215536 156136 215542 156188
rect 218054 156136 218060 156188
rect 218112 156176 218118 156188
rect 229066 156176 229094 156216
rect 266906 156204 266912 156216
rect 266964 156204 266970 156256
rect 218112 156148 229094 156176
rect 218112 156136 218118 156148
rect 230750 156136 230756 156188
rect 230808 156176 230814 156188
rect 277118 156176 277124 156188
rect 230808 156148 277124 156176
rect 230808 156136 230814 156148
rect 277118 156136 277124 156148
rect 277176 156136 277182 156188
rect 118200 156080 201264 156108
rect 118200 156068 118206 156080
rect 203058 156068 203064 156120
rect 203116 156108 203122 156120
rect 273898 156108 273904 156120
rect 203116 156080 273904 156108
rect 203116 156068 203122 156080
rect 273898 156068 273904 156080
rect 273956 156068 273962 156120
rect 121454 156000 121460 156052
rect 121512 156040 121518 156052
rect 197998 156040 198004 156052
rect 121512 156012 198004 156040
rect 121512 156000 121518 156012
rect 197998 156000 198004 156012
rect 198056 156000 198062 156052
rect 202230 156000 202236 156052
rect 202288 156040 202294 156052
rect 273254 156040 273260 156052
rect 202288 156012 273260 156040
rect 202288 156000 202294 156012
rect 273254 156000 273260 156012
rect 273312 156000 273318 156052
rect 145006 155932 145012 155984
rect 145064 155972 145070 155984
rect 229646 155972 229652 155984
rect 145064 155944 229652 155972
rect 145064 155932 145070 155944
rect 229646 155932 229652 155944
rect 229704 155932 229710 155984
rect 66806 155864 66812 155916
rect 66864 155904 66870 155916
rect 82906 155904 82912 155916
rect 66864 155876 82912 155904
rect 66864 155864 66870 155876
rect 82906 155864 82912 155876
rect 82964 155864 82970 155916
rect 88702 155864 88708 155916
rect 88760 155904 88766 155916
rect 186866 155904 186872 155916
rect 88760 155876 186872 155904
rect 88760 155864 88766 155876
rect 186866 155864 186872 155876
rect 186924 155864 186930 155916
rect 192938 155864 192944 155916
rect 192996 155904 193002 155916
rect 266262 155904 266268 155916
rect 192996 155876 266268 155904
rect 192996 155864 193002 155876
rect 266262 155864 266268 155876
rect 266320 155864 266326 155916
rect 296438 155864 296444 155916
rect 296496 155904 296502 155916
rect 345198 155904 345204 155916
rect 296496 155876 345204 155904
rect 296496 155864 296502 155876
rect 345198 155864 345204 155876
rect 345256 155864 345262 155916
rect 60090 155796 60096 155848
rect 60148 155836 60154 155848
rect 78766 155836 78772 155848
rect 60148 155808 78772 155836
rect 60148 155796 60154 155808
rect 78766 155796 78772 155808
rect 78824 155796 78830 155848
rect 89530 155796 89536 155848
rect 89588 155836 89594 155848
rect 186314 155836 186320 155848
rect 89588 155808 186320 155836
rect 89588 155796 89594 155808
rect 186314 155796 186320 155808
rect 186372 155796 186378 155848
rect 186406 155796 186412 155848
rect 186464 155836 186470 155848
rect 189534 155836 189540 155848
rect 186464 155808 189540 155836
rect 186464 155796 186470 155808
rect 189534 155796 189540 155808
rect 189592 155796 189598 155848
rect 189626 155796 189632 155848
rect 189684 155836 189690 155848
rect 263778 155836 263784 155848
rect 189684 155808 263784 155836
rect 189684 155796 189690 155808
rect 263778 155796 263784 155808
rect 263836 155796 263842 155848
rect 293034 155796 293040 155848
rect 293092 155836 293098 155848
rect 342346 155836 342352 155848
rect 293092 155808 342352 155836
rect 293092 155796 293098 155808
rect 342346 155796 342352 155808
rect 342404 155796 342410 155848
rect 12158 155728 12164 155780
rect 12216 155768 12222 155780
rect 110322 155768 110328 155780
rect 12216 155740 110328 155768
rect 12216 155728 12222 155740
rect 110322 155728 110328 155740
rect 110380 155728 110386 155780
rect 112254 155728 112260 155780
rect 112312 155768 112318 155780
rect 204622 155768 204628 155780
rect 112312 155740 204628 155768
rect 112312 155728 112318 155740
rect 204622 155728 204628 155740
rect 204680 155728 204686 155780
rect 206462 155728 206468 155780
rect 206520 155768 206526 155780
rect 276474 155768 276480 155780
rect 206520 155740 276480 155768
rect 206520 155728 206526 155740
rect 276474 155728 276480 155740
rect 276532 155728 276538 155780
rect 289722 155728 289728 155780
rect 289780 155768 289786 155780
rect 339586 155768 339592 155780
rect 289780 155740 339592 155768
rect 289780 155728 289786 155740
rect 339586 155728 339592 155740
rect 339644 155728 339650 155780
rect 46566 155660 46572 155712
rect 46624 155700 46630 155712
rect 75086 155700 75092 155712
rect 46624 155672 75092 155700
rect 46624 155660 46630 155672
rect 75086 155660 75092 155672
rect 75144 155660 75150 155712
rect 81894 155660 81900 155712
rect 81952 155700 81958 155712
rect 180978 155700 180984 155712
rect 81952 155672 180984 155700
rect 81952 155660 81958 155672
rect 180978 155660 180984 155672
rect 181036 155660 181042 155712
rect 186222 155660 186228 155712
rect 186280 155700 186286 155712
rect 260834 155700 260840 155712
rect 186280 155672 260840 155700
rect 186280 155660 186286 155672
rect 260834 155660 260840 155672
rect 260892 155660 260898 155712
rect 270310 155660 270316 155712
rect 270368 155700 270374 155712
rect 325326 155700 325332 155712
rect 270368 155672 325332 155700
rect 270368 155660 270374 155672
rect 325326 155660 325332 155672
rect 325384 155660 325390 155712
rect 344370 155660 344376 155712
rect 344428 155700 344434 155712
rect 381814 155700 381820 155712
rect 344428 155672 381820 155700
rect 344428 155660 344434 155672
rect 381814 155660 381820 155672
rect 381872 155660 381878 155712
rect 53374 155592 53380 155644
rect 53432 155632 53438 155644
rect 66622 155632 66628 155644
rect 53432 155604 66628 155632
rect 53432 155592 53438 155604
rect 66622 155592 66628 155604
rect 66680 155592 66686 155644
rect 71866 155592 71872 155644
rect 71924 155632 71930 155644
rect 172698 155632 172704 155644
rect 71924 155604 172704 155632
rect 71924 155592 71930 155604
rect 172698 155592 172704 155604
rect 172756 155592 172762 155644
rect 176102 155592 176108 155644
rect 176160 155632 176166 155644
rect 253382 155632 253388 155644
rect 176160 155604 253388 155632
rect 176160 155592 176166 155604
rect 253382 155592 253388 155604
rect 253440 155592 253446 155644
rect 266998 155592 267004 155644
rect 267056 155632 267062 155644
rect 322106 155632 322112 155644
rect 267056 155604 322112 155632
rect 267056 155592 267062 155604
rect 322106 155592 322112 155604
rect 322164 155592 322170 155644
rect 340966 155592 340972 155644
rect 341024 155632 341030 155644
rect 378134 155632 378140 155644
rect 341024 155604 378140 155632
rect 341024 155592 341030 155604
rect 378134 155592 378140 155604
rect 378192 155592 378198 155644
rect 39850 155524 39856 155576
rect 39908 155564 39914 155576
rect 68922 155564 68928 155576
rect 39908 155536 68928 155564
rect 39908 155524 39914 155536
rect 68922 155524 68928 155536
rect 68980 155524 68986 155576
rect 75178 155524 75184 155576
rect 75236 155564 75242 155576
rect 176378 155564 176384 155576
rect 75236 155536 176384 155564
rect 75236 155524 75242 155536
rect 176378 155524 176384 155536
rect 176436 155524 176442 155576
rect 179506 155524 179512 155576
rect 179564 155564 179570 155576
rect 255682 155564 255688 155576
rect 179564 155536 255688 155564
rect 179564 155524 179570 155536
rect 255682 155524 255688 155536
rect 255740 155524 255746 155576
rect 263594 155524 263600 155576
rect 263652 155564 263658 155576
rect 320174 155564 320180 155576
rect 263652 155536 320180 155564
rect 263652 155524 263658 155536
rect 320174 155524 320180 155536
rect 320232 155524 320238 155576
rect 337654 155524 337660 155576
rect 337712 155564 337718 155576
rect 375558 155564 375564 155576
rect 337712 155536 375564 155564
rect 337712 155524 337718 155536
rect 375558 155524 375564 155536
rect 375616 155524 375622 155576
rect 65150 155456 65156 155508
rect 65208 155496 65214 155508
rect 168650 155496 168656 155508
rect 65208 155468 168656 155496
rect 65208 155456 65214 155468
rect 168650 155456 168656 155468
rect 168708 155456 168714 155508
rect 169386 155456 169392 155508
rect 169444 155496 169450 155508
rect 248230 155496 248236 155508
rect 169444 155468 248236 155496
rect 169444 155456 169450 155468
rect 248230 155456 248236 155468
rect 248288 155456 248294 155508
rect 260282 155456 260288 155508
rect 260340 155496 260346 155508
rect 317598 155496 317604 155508
rect 260340 155468 317604 155496
rect 260340 155456 260346 155468
rect 317598 155456 317604 155468
rect 317656 155456 317662 155508
rect 333422 155456 333428 155508
rect 333480 155496 333486 155508
rect 373442 155496 373448 155508
rect 333480 155468 373448 155496
rect 333480 155456 333486 155468
rect 373442 155456 373448 155468
rect 373500 155456 373506 155508
rect 7926 155388 7932 155440
rect 7984 155428 7990 155440
rect 124674 155428 124680 155440
rect 7984 155400 124680 155428
rect 7984 155388 7990 155400
rect 124674 155388 124680 155400
rect 124732 155388 124738 155440
rect 149238 155388 149244 155440
rect 149296 155428 149302 155440
rect 232866 155428 232872 155440
rect 149296 155400 232872 155428
rect 149296 155388 149302 155400
rect 232866 155388 232872 155400
rect 232924 155388 232930 155440
rect 253566 155388 253572 155440
rect 253624 155428 253630 155440
rect 312446 155428 312452 155440
rect 253624 155400 312452 155428
rect 253624 155388 253630 155400
rect 312446 155388 312452 155400
rect 312504 155388 312510 155440
rect 330110 155388 330116 155440
rect 330168 155428 330174 155440
rect 370866 155428 370872 155440
rect 330168 155400 370872 155428
rect 330168 155388 330174 155400
rect 370866 155388 370872 155400
rect 370924 155388 370930 155440
rect 8754 155320 8760 155372
rect 8812 155360 8818 155372
rect 125686 155360 125692 155372
rect 8812 155332 125692 155360
rect 8812 155320 8818 155332
rect 125686 155320 125692 155332
rect 125744 155320 125750 155372
rect 145834 155320 145840 155372
rect 145892 155360 145898 155372
rect 229186 155360 229192 155372
rect 145892 155332 229192 155360
rect 145892 155320 145898 155332
rect 229186 155320 229192 155332
rect 229244 155320 229250 155372
rect 250162 155320 250168 155372
rect 250220 155360 250226 155372
rect 309870 155360 309876 155372
rect 250220 155332 309876 155360
rect 250220 155320 250226 155332
rect 309870 155320 309876 155332
rect 309928 155320 309934 155372
rect 319990 155320 319996 155372
rect 320048 155360 320054 155372
rect 363230 155360 363236 155372
rect 320048 155332 363236 155360
rect 320048 155320 320054 155332
rect 363230 155320 363236 155332
rect 363288 155320 363294 155372
rect 4522 155252 4528 155304
rect 4580 155292 4586 155304
rect 122006 155292 122012 155304
rect 4580 155264 122012 155292
rect 4580 155252 4586 155264
rect 122006 155252 122012 155264
rect 122064 155252 122070 155304
rect 142522 155252 142528 155304
rect 142580 155292 142586 155304
rect 227806 155292 227812 155304
rect 142580 155264 227812 155292
rect 142580 155252 142586 155264
rect 227806 155252 227812 155264
rect 227864 155252 227870 155304
rect 233326 155252 233332 155304
rect 233384 155292 233390 155304
rect 297082 155292 297088 155304
rect 233384 155264 297088 155292
rect 233384 155252 233390 155264
rect 297082 155252 297088 155264
rect 297140 155252 297146 155304
rect 299750 155252 299756 155304
rect 299808 155292 299814 155304
rect 347866 155292 347872 155304
rect 299808 155264 347872 155292
rect 299808 155252 299814 155264
rect 347866 155252 347872 155264
rect 347924 155252 347930 155304
rect 373810 155252 373816 155304
rect 373868 155292 373874 155304
rect 403158 155292 403164 155304
rect 373868 155264 403164 155292
rect 373868 155252 373874 155264
rect 403158 155252 403164 155264
rect 403216 155252 403222 155304
rect 5350 155184 5356 155236
rect 5408 155224 5414 155236
rect 123018 155224 123024 155236
rect 5408 155196 123024 155224
rect 5408 155184 5414 155196
rect 123018 155184 123024 155196
rect 123076 155184 123082 155236
rect 128998 155184 129004 155236
rect 129056 155224 129062 155236
rect 217410 155224 217416 155236
rect 129056 155196 217416 155224
rect 129056 155184 129062 155196
rect 217410 155184 217416 155196
rect 217468 155184 217474 155236
rect 240042 155184 240048 155236
rect 240100 155224 240106 155236
rect 302510 155224 302516 155236
rect 240100 155196 302516 155224
rect 240100 155184 240106 155196
rect 302510 155184 302516 155196
rect 302568 155184 302574 155236
rect 306558 155184 306564 155236
rect 306616 155224 306622 155236
rect 352466 155224 352472 155236
rect 306616 155196 352472 155224
rect 306616 155184 306622 155196
rect 352466 155184 352472 155196
rect 352524 155184 352530 155236
rect 370406 155184 370412 155236
rect 370464 155224 370470 155236
rect 401778 155224 401784 155236
rect 370464 155196 401784 155224
rect 370464 155184 370470 155196
rect 401778 155184 401784 155196
rect 401836 155184 401842 155236
rect 92014 155116 92020 155168
rect 92072 155156 92078 155168
rect 189166 155156 189172 155168
rect 92072 155128 189172 155156
rect 92072 155116 92078 155128
rect 189166 155116 189172 155128
rect 189224 155116 189230 155168
rect 189534 155116 189540 155168
rect 189592 155156 189598 155168
rect 194318 155156 194324 155168
rect 189592 155128 194324 155156
rect 189592 155116 189598 155128
rect 194318 155116 194324 155128
rect 194376 155116 194382 155168
rect 196342 155116 196348 155168
rect 196400 155156 196406 155168
rect 268838 155156 268844 155168
rect 196400 155128 268844 155156
rect 196400 155116 196406 155128
rect 268838 155116 268844 155128
rect 268896 155116 268902 155168
rect 95418 155048 95424 155100
rect 95476 155088 95482 155100
rect 95476 155060 186452 155088
rect 95476 155048 95482 155060
rect 98730 154980 98736 155032
rect 98788 155020 98794 155032
rect 186314 155020 186320 155032
rect 98788 154992 186320 155020
rect 98788 154980 98794 154992
rect 186314 154980 186320 154992
rect 186372 154980 186378 155032
rect 186424 155020 186452 155060
rect 186774 155048 186780 155100
rect 186832 155088 186838 155100
rect 186832 155060 195974 155088
rect 186832 155048 186838 155060
rect 191742 155020 191748 155032
rect 186424 154992 191748 155020
rect 191742 154980 191748 154992
rect 191800 154980 191806 155032
rect 195946 155020 195974 155060
rect 199654 155048 199660 155100
rect 199712 155088 199718 155100
rect 271414 155088 271420 155100
rect 199712 155060 271420 155088
rect 199712 155048 199718 155060
rect 271414 155048 271420 155060
rect 271472 155048 271478 155100
rect 303154 155048 303160 155100
rect 303212 155088 303218 155100
rect 350350 155088 350356 155100
rect 303212 155060 350356 155088
rect 303212 155048 303218 155060
rect 350350 155048 350356 155060
rect 350408 155048 350414 155100
rect 200114 155020 200120 155032
rect 195946 154992 200120 155020
rect 200114 154980 200120 154992
rect 200172 154980 200178 155032
rect 207014 154980 207020 155032
rect 207072 155020 207078 155032
rect 269482 155020 269488 155032
rect 207072 154992 269488 155020
rect 207072 154980 207078 154992
rect 269482 154980 269488 154992
rect 269540 154980 269546 155032
rect 15470 154912 15476 154964
rect 15528 154952 15534 154964
rect 109034 154952 109040 154964
rect 15528 154924 109040 154952
rect 15528 154912 15534 154924
rect 109034 154912 109040 154924
rect 109092 154912 109098 154964
rect 122282 154912 122288 154964
rect 122340 154952 122346 154964
rect 212258 154952 212264 154964
rect 122340 154924 212264 154952
rect 122340 154912 122346 154924
rect 212258 154912 212264 154924
rect 212316 154912 212322 154964
rect 214650 154912 214656 154964
rect 214708 154952 214714 154964
rect 261386 154952 261392 154964
rect 214708 154924 261392 154952
rect 214708 154912 214714 154924
rect 261386 154912 261392 154924
rect 261444 154912 261450 154964
rect 106366 154844 106372 154896
rect 106424 154884 106430 154896
rect 186406 154884 186412 154896
rect 106424 154856 186412 154884
rect 106424 154844 106430 154856
rect 186406 154844 186412 154856
rect 186464 154844 186470 154896
rect 186682 154844 186688 154896
rect 186740 154884 186746 154896
rect 245838 154884 245844 154896
rect 186740 154856 245844 154884
rect 186740 154844 186746 154856
rect 245838 154844 245844 154856
rect 245896 154844 245902 154896
rect 125778 154776 125784 154828
rect 125836 154816 125842 154828
rect 214834 154816 214840 154828
rect 125836 154788 214840 154816
rect 125836 154776 125842 154788
rect 214834 154776 214840 154788
rect 214892 154776 214898 154828
rect 275462 154816 275468 154828
rect 275112 154788 275468 154816
rect 110506 154708 110512 154760
rect 110564 154748 110570 154760
rect 139302 154748 139308 154760
rect 110564 154720 139308 154748
rect 110564 154708 110570 154720
rect 139302 154708 139308 154720
rect 139360 154708 139366 154760
rect 155954 154708 155960 154760
rect 156012 154748 156018 154760
rect 238018 154748 238024 154760
rect 156012 154720 238024 154748
rect 156012 154708 156018 154720
rect 238018 154708 238024 154720
rect 238076 154708 238082 154760
rect 109126 154640 109132 154692
rect 109184 154680 109190 154692
rect 133046 154680 133052 154692
rect 109184 154652 133052 154680
rect 109184 154640 109190 154652
rect 133046 154640 133052 154652
rect 133104 154640 133110 154692
rect 159358 154640 159364 154692
rect 159416 154680 159422 154692
rect 240594 154680 240600 154692
rect 159416 154652 240600 154680
rect 159416 154640 159422 154652
rect 240594 154640 240600 154652
rect 240652 154640 240658 154692
rect 114462 154572 114468 154624
rect 114520 154612 114526 154624
rect 119982 154612 119988 154624
rect 114520 154584 119988 154612
rect 114520 154572 114526 154584
rect 119982 154572 119988 154584
rect 120040 154572 120046 154624
rect 137094 154572 137100 154624
rect 137152 154612 137158 154624
rect 138198 154612 138204 154624
rect 137152 154584 138204 154612
rect 137152 154572 137158 154584
rect 138198 154572 138204 154584
rect 138256 154572 138262 154624
rect 154482 154572 154488 154624
rect 154540 154612 154546 154624
rect 156690 154612 156696 154624
rect 154540 154584 155172 154612
rect 154540 154572 154546 154584
rect 51074 154504 51080 154556
rect 51132 154544 51138 154556
rect 155034 154544 155040 154556
rect 51132 154516 155040 154544
rect 51132 154504 51138 154516
rect 155034 154504 155040 154516
rect 155092 154504 155098 154556
rect 155144 154544 155172 154584
rect 156524 154584 156696 154612
rect 156524 154544 156552 154584
rect 156690 154572 156696 154584
rect 156748 154572 156754 154624
rect 162670 154572 162676 154624
rect 162728 154612 162734 154624
rect 243078 154612 243084 154624
rect 162728 154584 243084 154612
rect 162728 154572 162734 154584
rect 243078 154572 243084 154584
rect 243136 154572 243142 154624
rect 155144 154516 156552 154544
rect 156598 154504 156604 154556
rect 156656 154544 156662 154556
rect 212902 154544 212908 154556
rect 156656 154516 212908 154544
rect 156656 154504 156662 154516
rect 212902 154504 212908 154516
rect 212960 154504 212966 154556
rect 215294 154504 215300 154556
rect 215352 154544 215358 154556
rect 275112 154544 275140 154788
rect 275462 154776 275468 154788
rect 275520 154776 275526 154828
rect 275388 154720 275600 154748
rect 275388 154544 275416 154720
rect 275462 154640 275468 154692
rect 275520 154640 275526 154692
rect 215352 154516 275140 154544
rect 275296 154516 275416 154544
rect 215352 154504 215358 154516
rect 44174 154436 44180 154488
rect 44232 154476 44238 154488
rect 142522 154476 142528 154488
rect 44232 154448 142528 154476
rect 44232 154436 44238 154448
rect 142522 154436 142528 154448
rect 142580 154436 142586 154488
rect 142798 154436 142804 154488
rect 142856 154476 142862 154488
rect 188430 154476 188436 154488
rect 142856 154448 188436 154476
rect 142856 154436 142862 154448
rect 188430 154436 188436 154448
rect 188488 154436 188494 154488
rect 202690 154476 202696 154488
rect 188632 154448 202696 154476
rect 115934 154368 115940 154420
rect 115992 154408 115998 154420
rect 119890 154408 119896 154420
rect 115992 154380 119896 154408
rect 115992 154368 115998 154380
rect 119890 154368 119896 154380
rect 119948 154368 119954 154420
rect 119982 154368 119988 154420
rect 120040 154408 120046 154420
rect 185394 154408 185400 154420
rect 120040 154380 185400 154408
rect 120040 154368 120046 154380
rect 185394 154368 185400 154380
rect 185452 154368 185458 154420
rect 185504 154380 185808 154408
rect 34514 154300 34520 154352
rect 34572 154340 34578 154352
rect 142614 154340 142620 154352
rect 34572 154312 142620 154340
rect 34572 154300 34578 154312
rect 142614 154300 142620 154312
rect 142672 154300 142678 154352
rect 142706 154300 142712 154352
rect 142764 154340 142770 154352
rect 185504 154340 185532 154380
rect 142764 154312 185532 154340
rect 185780 154340 185808 154380
rect 185854 154368 185860 154420
rect 185912 154408 185918 154420
rect 188632 154408 188660 154448
rect 202690 154436 202696 154448
rect 202748 154436 202754 154488
rect 218330 154436 218336 154488
rect 218388 154476 218394 154488
rect 275296 154476 275324 154516
rect 218388 154448 275324 154476
rect 275480 154476 275508 154640
rect 275572 154544 275600 154720
rect 282932 154584 283880 154612
rect 282932 154544 282960 154584
rect 275572 154516 282960 154544
rect 283006 154504 283012 154556
rect 283064 154544 283070 154556
rect 283742 154544 283748 154556
rect 283064 154516 283748 154544
rect 283064 154504 283070 154516
rect 283742 154504 283748 154516
rect 283800 154504 283806 154556
rect 283650 154476 283656 154488
rect 275480 154448 283656 154476
rect 218388 154436 218394 154448
rect 283650 154436 283656 154448
rect 283708 154436 283714 154488
rect 283852 154476 283880 154584
rect 283926 154504 283932 154556
rect 283984 154544 283990 154556
rect 334894 154544 334900 154556
rect 283984 154516 334900 154544
rect 283984 154504 283990 154516
rect 334894 154504 334900 154516
rect 334952 154504 334958 154556
rect 353662 154504 353668 154556
rect 353720 154544 353726 154556
rect 388898 154544 388904 154556
rect 353720 154516 388904 154544
rect 353720 154504 353726 154516
rect 388898 154504 388904 154516
rect 388956 154504 388962 154556
rect 285582 154476 285588 154488
rect 283852 154448 285588 154476
rect 285582 154436 285588 154448
rect 285640 154436 285646 154488
rect 285674 154436 285680 154488
rect 285732 154476 285738 154488
rect 337470 154476 337476 154488
rect 285732 154448 337476 154476
rect 285732 154436 285738 154448
rect 337470 154436 337476 154448
rect 337528 154436 337534 154488
rect 349522 154436 349528 154488
rect 349580 154476 349586 154488
rect 386322 154476 386328 154488
rect 349580 154448 386328 154476
rect 349580 154436 349586 154448
rect 386322 154436 386328 154448
rect 386380 154436 386386 154488
rect 390646 154436 390652 154488
rect 390704 154476 390710 154488
rect 417142 154476 417148 154488
rect 390704 154448 417148 154476
rect 390704 154436 390710 154448
rect 417142 154436 417148 154448
rect 417200 154436 417206 154488
rect 185912 154380 188660 154408
rect 185912 154368 185918 154380
rect 191006 154368 191012 154420
rect 191064 154408 191070 154420
rect 202046 154408 202052 154420
rect 191064 154380 202052 154408
rect 191064 154368 191070 154380
rect 202046 154368 202052 154380
rect 202104 154368 202110 154420
rect 204990 154368 204996 154420
rect 205048 154408 205054 154420
rect 275278 154408 275284 154420
rect 205048 154380 275284 154408
rect 205048 154368 205054 154380
rect 275278 154368 275284 154380
rect 275336 154368 275342 154420
rect 276198 154368 276204 154420
rect 276256 154408 276262 154420
rect 329926 154408 329932 154420
rect 276256 154380 329932 154408
rect 276256 154368 276262 154380
rect 329926 154368 329932 154380
rect 329984 154368 329990 154420
rect 346394 154368 346400 154420
rect 346452 154408 346458 154420
rect 383746 154408 383752 154420
rect 346452 154380 383752 154408
rect 346452 154368 346458 154380
rect 383746 154368 383752 154380
rect 383804 154368 383810 154420
rect 393314 154368 393320 154420
rect 393372 154408 393378 154420
rect 419718 154408 419724 154420
rect 393372 154380 419724 154408
rect 393372 154368 393378 154380
rect 419718 154368 419724 154380
rect 419776 154368 419782 154420
rect 205266 154340 205272 154352
rect 185780 154312 205272 154340
rect 142764 154300 142770 154312
rect 205266 154300 205272 154312
rect 205324 154300 205330 154352
rect 208394 154300 208400 154352
rect 208452 154340 208458 154352
rect 278406 154340 278412 154352
rect 208452 154312 278412 154340
rect 208452 154300 208458 154312
rect 278406 154300 278412 154312
rect 278464 154300 278470 154352
rect 278866 154300 278872 154352
rect 278924 154340 278930 154352
rect 332410 154340 332416 154352
rect 278924 154312 332416 154340
rect 278924 154300 278930 154312
rect 332410 154300 332416 154312
rect 332468 154300 332474 154352
rect 336826 154300 336832 154352
rect 336884 154340 336890 154352
rect 376018 154340 376024 154352
rect 336884 154312 376024 154340
rect 336884 154300 336890 154312
rect 376018 154300 376024 154312
rect 376076 154300 376082 154352
rect 397362 154300 397368 154352
rect 397420 154340 397426 154352
rect 422478 154340 422484 154352
rect 397420 154312 422484 154340
rect 397420 154300 397426 154312
rect 422478 154300 422484 154312
rect 422536 154300 422542 154352
rect 37918 154232 37924 154284
rect 37976 154272 37982 154284
rect 37976 154244 142936 154272
rect 37976 154232 37982 154244
rect 27246 154164 27252 154216
rect 27304 154204 27310 154216
rect 136910 154204 136916 154216
rect 27304 154176 136916 154204
rect 27304 154164 27310 154176
rect 136910 154164 136916 154176
rect 136968 154164 136974 154216
rect 142798 154204 142804 154216
rect 137112 154176 142804 154204
rect 23474 154096 23480 154148
rect 23532 154136 23538 154148
rect 137002 154136 137008 154148
rect 23532 154108 137008 154136
rect 23532 154096 23538 154108
rect 137002 154096 137008 154108
rect 137060 154096 137066 154148
rect 13814 154028 13820 154080
rect 13872 154068 13878 154080
rect 129458 154068 129464 154080
rect 13872 154040 129464 154068
rect 13872 154028 13878 154040
rect 129458 154028 129464 154040
rect 129516 154028 129522 154080
rect 137112 154068 137140 154176
rect 142798 154164 142804 154176
rect 142856 154164 142862 154216
rect 142430 154136 142436 154148
rect 129568 154040 137140 154068
rect 137204 154108 142436 154136
rect 9674 153960 9680 154012
rect 9732 154000 9738 154012
rect 126882 154000 126888 154012
rect 9732 153972 126888 154000
rect 9732 153960 9738 153972
rect 126882 153960 126888 153972
rect 126940 153960 126946 154012
rect 129568 154000 129596 154040
rect 137204 154000 137232 154108
rect 142430 154096 142436 154108
rect 142488 154096 142494 154148
rect 142908 154136 142936 154244
rect 143166 154232 143172 154284
rect 143224 154272 143230 154284
rect 185302 154272 185308 154284
rect 143224 154244 185308 154272
rect 143224 154232 143230 154244
rect 185302 154232 185308 154244
rect 185360 154232 185366 154284
rect 185762 154232 185768 154284
rect 185820 154272 185826 154284
rect 186866 154272 186872 154284
rect 185820 154244 186872 154272
rect 185820 154232 185826 154244
rect 186866 154232 186872 154244
rect 186924 154232 186930 154284
rect 186958 154232 186964 154284
rect 187016 154272 187022 154284
rect 258534 154272 258540 154284
rect 187016 154244 258540 154272
rect 187016 154232 187022 154244
rect 258534 154232 258540 154244
rect 258592 154232 258598 154284
rect 262214 154232 262220 154284
rect 262272 154272 262278 154284
rect 319530 154272 319536 154284
rect 262272 154244 319536 154272
rect 262272 154232 262278 154244
rect 319530 154232 319536 154244
rect 319588 154232 319594 154284
rect 339494 154232 339500 154284
rect 339552 154272 339558 154284
rect 378594 154272 378600 154284
rect 339552 154244 378600 154272
rect 339552 154232 339558 154244
rect 378594 154232 378600 154244
rect 378652 154232 378658 154284
rect 386506 154232 386512 154284
rect 386564 154272 386570 154284
rect 414566 154272 414572 154284
rect 386564 154244 414572 154272
rect 386564 154232 386570 154244
rect 414566 154232 414572 154244
rect 414624 154232 414630 154284
rect 147582 154204 147588 154216
rect 143276 154176 147588 154204
rect 143276 154136 143304 154176
rect 147582 154164 147588 154176
rect 147640 154164 147646 154216
rect 147766 154164 147772 154216
rect 147824 154204 147830 154216
rect 156598 154204 156604 154216
rect 147824 154176 156604 154204
rect 147824 154164 147830 154176
rect 156598 154164 156604 154176
rect 156656 154164 156662 154216
rect 172514 154164 172520 154216
rect 172572 154204 172578 154216
rect 250806 154204 250812 154216
rect 172572 154176 250812 154204
rect 172572 154164 172578 154176
rect 250806 154164 250812 154176
rect 250864 154164 250870 154216
rect 255314 154164 255320 154216
rect 255372 154204 255378 154216
rect 314378 154204 314384 154216
rect 255372 154176 314384 154204
rect 255372 154164 255378 154176
rect 314378 154164 314384 154176
rect 314436 154164 314442 154216
rect 343542 154164 343548 154216
rect 343600 154204 343606 154216
rect 381170 154204 381176 154216
rect 343600 154176 381176 154204
rect 343600 154164 343606 154176
rect 381170 154164 381176 154176
rect 381228 154164 381234 154216
rect 383654 154164 383660 154216
rect 383712 154204 383718 154216
rect 411990 154204 411996 154216
rect 383712 154176 411996 154204
rect 383712 154164 383718 154176
rect 411990 154164 411996 154176
rect 412048 154164 412054 154216
rect 142908 154108 143304 154136
rect 143442 154096 143448 154148
rect 143500 154136 143506 154148
rect 145558 154136 145564 154148
rect 143500 154108 145564 154136
rect 143500 154096 143506 154108
rect 145558 154096 145564 154108
rect 145616 154096 145622 154148
rect 147122 154096 147128 154148
rect 147180 154136 147186 154148
rect 147180 154108 156460 154136
rect 147180 154096 147186 154108
rect 138382 154028 138388 154080
rect 138440 154068 138446 154080
rect 143166 154068 143172 154080
rect 138440 154040 143172 154068
rect 138440 154028 138446 154040
rect 143166 154028 143172 154040
rect 143224 154028 143230 154080
rect 143350 154028 143356 154080
rect 143408 154068 143414 154080
rect 150618 154068 150624 154080
rect 143408 154040 150624 154068
rect 143408 154028 143414 154040
rect 150618 154028 150624 154040
rect 150676 154028 150682 154080
rect 151814 154028 151820 154080
rect 151872 154068 151878 154080
rect 155862 154068 155868 154080
rect 151872 154040 155868 154068
rect 151872 154028 151878 154040
rect 155862 154028 155868 154040
rect 155920 154028 155926 154080
rect 156432 154068 156460 154108
rect 156506 154096 156512 154148
rect 156564 154136 156570 154148
rect 163498 154136 163504 154148
rect 156564 154108 163504 154136
rect 156564 154096 156570 154108
rect 163498 154096 163504 154108
rect 163556 154096 163562 154148
rect 165614 154096 165620 154148
rect 165672 154136 165678 154148
rect 245654 154136 245660 154148
rect 165672 154108 245660 154136
rect 165672 154096 165678 154108
rect 245654 154096 245660 154108
rect 245712 154096 245718 154148
rect 245930 154096 245936 154148
rect 245988 154136 245994 154148
rect 306650 154136 306656 154148
rect 245988 154108 306656 154136
rect 245988 154096 245994 154108
rect 306650 154096 306656 154108
rect 306708 154096 306714 154148
rect 326706 154096 326712 154148
rect 326764 154136 326770 154148
rect 368290 154136 368296 154148
rect 326764 154108 368296 154136
rect 326764 154096 326770 154108
rect 368290 154096 368296 154108
rect 368348 154096 368354 154148
rect 376846 154096 376852 154148
rect 376904 154136 376910 154148
rect 406838 154136 406844 154148
rect 376904 154108 406844 154136
rect 376904 154096 376910 154108
rect 406838 154096 406844 154108
rect 406896 154096 406902 154148
rect 156598 154068 156604 154080
rect 156432 154040 156604 154068
rect 156598 154028 156604 154040
rect 156656 154028 156662 154080
rect 156690 154028 156696 154080
rect 156748 154068 156754 154080
rect 158530 154068 158536 154080
rect 156748 154040 158536 154068
rect 156748 154028 156754 154040
rect 158530 154028 158536 154040
rect 158588 154028 158594 154080
rect 160186 154028 160192 154080
rect 160244 154068 160250 154080
rect 241238 154068 241244 154080
rect 160244 154040 241244 154068
rect 160244 154028 160250 154040
rect 241238 154028 241244 154040
rect 241296 154028 241302 154080
rect 248598 154028 248604 154080
rect 248656 154068 248662 154080
rect 309226 154068 309232 154080
rect 248656 154040 309232 154068
rect 248656 154028 248662 154040
rect 309226 154028 309232 154040
rect 309284 154028 309290 154080
rect 323302 154028 323308 154080
rect 323360 154068 323366 154080
rect 365806 154068 365812 154080
rect 323360 154040 365812 154068
rect 323360 154028 323366 154040
rect 365806 154028 365812 154040
rect 365864 154028 365870 154080
rect 380158 154028 380164 154080
rect 380216 154068 380222 154080
rect 409414 154068 409420 154080
rect 380216 154040 409420 154068
rect 380216 154028 380222 154040
rect 409414 154028 409420 154040
rect 409472 154028 409478 154080
rect 219894 154000 219900 154012
rect 126992 153972 129596 154000
rect 129660 153972 137232 154000
rect 139780 153972 219900 154000
rect 7098 153892 7104 153944
rect 7156 153932 7162 153944
rect 124306 153932 124312 153944
rect 7156 153904 124312 153932
rect 7156 153892 7162 153904
rect 124306 153892 124312 153904
rect 124364 153892 124370 153944
rect 125502 153892 125508 153944
rect 125560 153932 125566 153944
rect 126992 153932 127020 153972
rect 127710 153932 127716 153944
rect 125560 153904 127020 153932
rect 127544 153904 127716 153932
rect 125560 153892 125566 153904
rect 474 153824 480 153876
rect 532 153864 538 153876
rect 119798 153864 119804 153876
rect 532 153836 119804 153864
rect 532 153824 538 153836
rect 119798 153824 119804 153836
rect 119856 153824 119862 153876
rect 119890 153824 119896 153876
rect 119948 153864 119954 153876
rect 127544 153864 127572 153904
rect 127710 153892 127716 153904
rect 127768 153892 127774 153944
rect 127802 153892 127808 153944
rect 127860 153932 127866 153944
rect 129660 153932 129688 153972
rect 127860 153904 129688 153932
rect 127860 153892 127866 153904
rect 132402 153892 132408 153944
rect 132460 153932 132466 153944
rect 139780 153932 139808 153972
rect 219894 153960 219900 153972
rect 219952 153960 219958 154012
rect 222378 153960 222384 154012
rect 222436 154000 222442 154012
rect 288710 154000 288716 154012
rect 222436 153972 288716 154000
rect 222436 153960 222442 153972
rect 288710 153960 288716 153972
rect 288768 153960 288774 154012
rect 313274 153960 313280 154012
rect 313332 154000 313338 154012
rect 357894 154000 357900 154012
rect 313332 153972 357900 154000
rect 313332 153960 313338 153972
rect 357894 153960 357900 153972
rect 357952 153960 357958 154012
rect 367094 153960 367100 154012
rect 367152 154000 367158 154012
rect 399110 154000 399116 154012
rect 367152 153972 399116 154000
rect 367152 153960 367158 153972
rect 399110 153960 399116 153972
rect 399168 153960 399174 154012
rect 132460 153904 139808 153932
rect 132460 153892 132466 153904
rect 139854 153892 139860 153944
rect 139912 153932 139918 153944
rect 142430 153932 142436 153944
rect 139912 153904 142436 153932
rect 139912 153892 139918 153904
rect 142430 153892 142436 153904
rect 142488 153892 142494 153944
rect 142522 153892 142528 153944
rect 142580 153932 142586 153944
rect 142580 153904 142936 153932
rect 142580 153892 142586 153904
rect 119948 153836 127572 153864
rect 119948 153824 119954 153836
rect 127618 153824 127624 153876
rect 127676 153864 127682 153876
rect 142798 153864 142804 153876
rect 127676 153836 142804 153864
rect 127676 153824 127682 153836
rect 142798 153824 142804 153836
rect 142856 153824 142862 153876
rect 142908 153864 142936 153904
rect 142982 153892 142988 153944
rect 143040 153932 143046 153944
rect 223206 153932 223212 153944
rect 143040 153904 223212 153932
rect 143040 153892 143046 153904
rect 223206 153892 223212 153904
rect 223264 153892 223270 153944
rect 225230 153892 225236 153944
rect 225288 153932 225294 153944
rect 291286 153932 291292 153944
rect 225288 153904 291292 153932
rect 225288 153892 225294 153904
rect 291286 153892 291292 153904
rect 291344 153892 291350 153944
rect 316034 153892 316040 153944
rect 316092 153932 316098 153944
rect 360654 153932 360660 153944
rect 316092 153904 360660 153932
rect 316092 153892 316098 153904
rect 360654 153892 360660 153904
rect 360712 153892 360718 153944
rect 363046 153892 363052 153944
rect 363104 153932 363110 153944
rect 396534 153932 396540 153944
rect 363104 153904 396540 153932
rect 363104 153892 363110 153904
rect 396534 153892 396540 153904
rect 396592 153892 396598 153944
rect 401594 153892 401600 153944
rect 401652 153932 401658 153944
rect 425514 153932 425520 153944
rect 401652 153904 425520 153932
rect 401652 153892 401658 153904
rect 425514 153892 425520 153904
rect 425572 153892 425578 153944
rect 153286 153864 153292 153876
rect 142908 153836 153292 153864
rect 153286 153824 153292 153836
rect 153344 153824 153350 153876
rect 155034 153824 155040 153876
rect 155092 153864 155098 153876
rect 158346 153864 158352 153876
rect 155092 153836 158352 153864
rect 155092 153824 155098 153836
rect 158346 153824 158352 153836
rect 158404 153824 158410 153876
rect 235442 153864 235448 153876
rect 158456 153836 235448 153864
rect 48314 153756 48320 153808
rect 48372 153796 48378 153808
rect 155770 153796 155776 153808
rect 48372 153768 155776 153796
rect 48372 153756 48378 153768
rect 155770 153756 155776 153768
rect 155828 153756 155834 153808
rect 155862 153756 155868 153808
rect 155920 153796 155926 153808
rect 158456 153796 158484 153836
rect 235442 153824 235448 153836
rect 235500 153824 235506 153876
rect 241882 153824 241888 153876
rect 241940 153864 241946 153876
rect 304074 153864 304080 153876
rect 241940 153836 304080 153864
rect 241940 153824 241946 153836
rect 304074 153824 304080 153836
rect 304132 153824 304138 153876
rect 309134 153824 309140 153876
rect 309192 153864 309198 153876
rect 355502 153864 355508 153876
rect 309192 153836 355508 153864
rect 309192 153824 309198 153836
rect 355502 153824 355508 153836
rect 355560 153824 355566 153876
rect 356238 153824 356244 153876
rect 356296 153864 356302 153876
rect 391474 153864 391480 153876
rect 356296 153836 391480 153864
rect 356296 153824 356302 153836
rect 391474 153824 391480 153836
rect 391532 153824 391538 153876
rect 397454 153824 397460 153876
rect 397512 153864 397518 153876
rect 423030 153864 423036 153876
rect 397512 153836 423036 153864
rect 397512 153824 397518 153836
rect 423030 153824 423036 153836
rect 423088 153824 423094 153876
rect 155920 153768 158484 153796
rect 155920 153756 155926 153768
rect 158530 153756 158536 153808
rect 158588 153796 158594 153808
rect 218054 153796 218060 153808
rect 158588 153768 218060 153796
rect 158588 153756 158594 153768
rect 218054 153756 218060 153768
rect 218112 153756 218118 153808
rect 231854 153756 231860 153808
rect 231912 153796 231918 153808
rect 296438 153796 296444 153808
rect 231912 153768 296444 153796
rect 231912 153756 231918 153768
rect 296438 153756 296444 153768
rect 296496 153756 296502 153808
rect 360378 153756 360384 153808
rect 360436 153796 360442 153808
rect 394050 153796 394056 153808
rect 360436 153768 394056 153796
rect 360436 153756 360442 153768
rect 394050 153756 394056 153768
rect 394108 153756 394114 153808
rect 61102 153688 61108 153740
rect 61160 153728 61166 153740
rect 166074 153728 166080 153740
rect 61160 153700 166080 153728
rect 61160 153688 61166 153700
rect 166074 153688 166080 153700
rect 166132 153688 166138 153740
rect 210418 153728 210424 153740
rect 171106 153700 210424 153728
rect 57974 153620 57980 153672
rect 58032 153660 58038 153672
rect 156506 153660 156512 153672
rect 58032 153632 156512 153660
rect 58032 153620 58038 153632
rect 156506 153620 156512 153632
rect 156564 153620 156570 153672
rect 156598 153620 156604 153672
rect 156656 153660 156662 153672
rect 171106 153660 171134 153700
rect 210418 153688 210424 153700
rect 210476 153688 210482 153740
rect 229094 153688 229100 153740
rect 229152 153728 229158 153740
rect 293862 153728 293868 153740
rect 229152 153700 293868 153728
rect 229152 153688 229158 153700
rect 293862 153688 293868 153700
rect 293920 153688 293926 153740
rect 156656 153632 171134 153660
rect 156656 153620 156662 153632
rect 176654 153620 176660 153672
rect 176712 153660 176718 153672
rect 176712 153632 180794 153660
rect 176712 153620 176718 153632
rect 78674 153552 78680 153604
rect 78732 153592 78738 153604
rect 179598 153592 179604 153604
rect 78732 153564 179604 153592
rect 78732 153552 78738 153564
rect 179598 153552 179604 153564
rect 179656 153552 179662 153604
rect 180766 153592 180794 153632
rect 182174 153620 182180 153672
rect 182232 153660 182238 153672
rect 186958 153660 186964 153672
rect 182232 153632 186964 153660
rect 182232 153620 182238 153632
rect 186958 153620 186964 153632
rect 187016 153620 187022 153672
rect 188430 153620 188436 153672
rect 188488 153660 188494 153672
rect 195974 153660 195980 153672
rect 188488 153632 195980 153660
rect 188488 153620 188494 153632
rect 195974 153620 195980 153632
rect 196032 153620 196038 153672
rect 196066 153620 196072 153672
rect 196124 153660 196130 153672
rect 196124 153632 233924 153660
rect 196124 153620 196130 153632
rect 230934 153592 230940 153604
rect 180766 153564 230940 153592
rect 230934 153552 230940 153564
rect 230992 153552 230998 153604
rect 233896 153592 233924 153632
rect 235074 153620 235080 153672
rect 235132 153660 235138 153672
rect 299014 153660 299020 153672
rect 235132 153632 299020 153660
rect 235132 153620 235138 153632
rect 299014 153620 299020 153632
rect 299072 153620 299078 153672
rect 238662 153592 238668 153604
rect 233896 153564 238668 153592
rect 238662 153552 238668 153564
rect 238720 153552 238726 153604
rect 238846 153552 238852 153604
rect 238904 153592 238910 153604
rect 301590 153592 301596 153604
rect 238904 153564 301596 153592
rect 238904 153552 238910 153564
rect 301590 153552 301596 153564
rect 301648 153552 301654 153604
rect 102134 153484 102140 153536
rect 102192 153524 102198 153536
rect 196894 153524 196900 153536
rect 102192 153496 196900 153524
rect 102192 153484 102198 153496
rect 196894 153484 196900 153496
rect 196952 153484 196958 153536
rect 198918 153484 198924 153536
rect 198976 153524 198982 153536
rect 248874 153524 248880 153536
rect 198976 153496 248880 153524
rect 198976 153484 198982 153496
rect 248874 153484 248880 153496
rect 248932 153484 248938 153536
rect 252646 153484 252652 153536
rect 252704 153524 252710 153536
rect 311802 153524 311808 153536
rect 252704 153496 311808 153524
rect 252704 153484 252710 153496
rect 311802 153484 311808 153496
rect 311860 153484 311866 153536
rect 104894 153416 104900 153468
rect 104952 153456 104958 153468
rect 196526 153456 196532 153468
rect 104952 153428 196532 153456
rect 104952 153416 104958 153428
rect 196526 153416 196532 153428
rect 196584 153416 196590 153468
rect 196986 153416 196992 153468
rect 197044 153456 197050 153468
rect 197044 153428 197676 153456
rect 197044 153416 197050 153428
rect 108298 153348 108304 153400
rect 108356 153388 108362 153400
rect 191006 153388 191012 153400
rect 108356 153360 191012 153388
rect 108356 153348 108362 153360
rect 191006 153348 191012 153360
rect 191064 153348 191070 153400
rect 191650 153348 191656 153400
rect 191708 153388 191714 153400
rect 195882 153388 195888 153400
rect 191708 153360 195888 153388
rect 191708 153348 191714 153360
rect 195882 153348 195888 153360
rect 195940 153348 195946 153400
rect 195974 153348 195980 153400
rect 196032 153388 196038 153400
rect 197538 153388 197544 153400
rect 196032 153360 197544 153388
rect 196032 153348 196038 153360
rect 197538 153348 197544 153360
rect 197596 153348 197602 153400
rect 197648 153388 197676 153428
rect 201402 153416 201408 153468
rect 201460 153456 201466 153468
rect 259178 153456 259184 153468
rect 201460 153428 259184 153456
rect 201460 153416 201466 153428
rect 259178 153416 259184 153428
rect 259236 153416 259242 153468
rect 265434 153416 265440 153468
rect 265492 153456 265498 153468
rect 322014 153456 322020 153468
rect 265492 153428 322020 153456
rect 265492 153416 265498 153428
rect 322014 153416 322020 153428
rect 322072 153416 322078 153468
rect 243722 153388 243728 153400
rect 197648 153360 243728 153388
rect 243722 153348 243728 153360
rect 243780 153348 243786 153400
rect 259454 153348 259460 153400
rect 259512 153388 259518 153400
rect 316954 153388 316960 153400
rect 259512 153360 316960 153388
rect 259512 153348 259518 153360
rect 316954 153348 316960 153360
rect 317012 153348 317018 153400
rect 41598 153280 41604 153332
rect 41656 153320 41662 153332
rect 142706 153320 142712 153332
rect 41656 153292 142712 153320
rect 41656 153280 41662 153292
rect 142706 153280 142712 153292
rect 142764 153280 142770 153332
rect 142798 153280 142804 153332
rect 142856 153320 142862 153332
rect 209774 153320 209780 153332
rect 142856 153292 209780 153320
rect 142856 153280 142862 153292
rect 209774 153280 209780 153292
rect 209832 153280 209838 153332
rect 269206 153280 269212 153332
rect 269264 153320 269270 153332
rect 324682 153320 324688 153332
rect 269264 153292 324688 153320
rect 269264 153280 269270 153292
rect 324682 153280 324688 153292
rect 324740 153280 324746 153332
rect 118694 153212 118700 153264
rect 118752 153252 118758 153264
rect 127618 153252 127624 153264
rect 118752 153224 127624 153252
rect 118752 153212 118758 153224
rect 127618 153212 127624 153224
rect 127676 153212 127682 153264
rect 127710 153212 127716 153264
rect 127768 153252 127774 153264
rect 207842 153252 207848 153264
rect 127768 153224 207848 153252
rect 127768 153212 127774 153224
rect 207842 153212 207848 153224
rect 207900 153212 207906 153264
rect 272886 153212 272892 153264
rect 272944 153252 272950 153264
rect 327258 153252 327264 153264
rect 272944 153224 327264 153252
rect 272944 153212 272950 153224
rect 327258 153212 327264 153224
rect 327316 153212 327322 153264
rect 442920 153224 444328 153252
rect 23290 153144 23296 153196
rect 23348 153184 23354 153196
rect 110966 153184 110972 153196
rect 23348 153156 110972 153184
rect 23348 153144 23354 153156
rect 110966 153144 110972 153156
rect 111024 153144 111030 153196
rect 113174 153144 113180 153196
rect 113232 153184 113238 153196
rect 205910 153184 205916 153196
rect 113232 153156 205916 153184
rect 113232 153144 113238 153156
rect 205910 153144 205916 153156
rect 205968 153144 205974 153196
rect 215386 153144 215392 153196
rect 215444 153184 215450 153196
rect 279694 153184 279700 153196
rect 215444 153156 279700 153184
rect 215444 153144 215450 153156
rect 279694 153144 279700 153156
rect 279752 153144 279758 153196
rect 285490 153144 285496 153196
rect 285548 153184 285554 153196
rect 336826 153184 336832 153196
rect 285548 153156 336832 153184
rect 285548 153144 285554 153156
rect 336826 153144 336832 153156
rect 336884 153144 336890 153196
rect 339678 153144 339684 153196
rect 339736 153184 339742 153196
rect 377306 153184 377312 153196
rect 339736 153156 377312 153184
rect 339736 153144 339742 153156
rect 377306 153144 377312 153156
rect 377364 153144 377370 153196
rect 378226 153144 378232 153196
rect 378284 153184 378290 153196
rect 379882 153184 379888 153196
rect 378284 153156 379888 153184
rect 378284 153144 378290 153156
rect 379882 153144 379888 153156
rect 379940 153144 379946 153196
rect 380986 153144 380992 153196
rect 381044 153184 381050 153196
rect 410058 153184 410064 153196
rect 381044 153156 410064 153184
rect 381044 153144 381050 153156
rect 410058 153144 410064 153156
rect 410116 153144 410122 153196
rect 412910 153144 412916 153196
rect 412968 153184 412974 153196
rect 433794 153184 433800 153196
rect 412968 153156 433800 153184
rect 412968 153144 412974 153156
rect 433794 153144 433800 153156
rect 433852 153144 433858 153196
rect 434346 153144 434352 153196
rect 434404 153184 434410 153196
rect 441614 153184 441620 153196
rect 434404 153156 441620 153184
rect 434404 153144 434410 153156
rect 441614 153144 441620 153156
rect 441672 153144 441678 153196
rect 441706 153144 441712 153196
rect 441764 153184 441770 153196
rect 442920 153184 442948 153224
rect 441764 153156 442948 153184
rect 441764 153144 441770 153156
rect 442994 153144 443000 153196
rect 443052 153184 443058 153196
rect 444190 153184 444196 153196
rect 443052 153156 444196 153184
rect 443052 153144 443058 153156
rect 444190 153144 444196 153156
rect 444248 153144 444254 153196
rect 444300 153184 444328 153224
rect 449250 153184 449256 153196
rect 444300 153156 449256 153184
rect 449250 153144 449256 153156
rect 449308 153144 449314 153196
rect 453942 153144 453948 153196
rect 454000 153184 454006 153196
rect 459462 153184 459468 153196
rect 454000 153156 459468 153184
rect 454000 153144 454006 153156
rect 459462 153144 459468 153156
rect 459520 153144 459526 153196
rect 462222 153144 462228 153196
rect 462280 153184 462286 153196
rect 465902 153184 465908 153196
rect 462280 153156 465908 153184
rect 462280 153144 462286 153156
rect 465902 153144 465908 153156
rect 465960 153144 465966 153196
rect 466454 153144 466460 153196
rect 466512 153184 466518 153196
rect 469766 153184 469772 153196
rect 466512 153156 469772 153184
rect 466512 153144 466518 153156
rect 469766 153144 469772 153156
rect 469824 153144 469830 153196
rect 471330 153144 471336 153196
rect 471388 153184 471394 153196
rect 472986 153184 472992 153196
rect 471388 153156 472992 153184
rect 471388 153144 471394 153156
rect 472986 153144 472992 153156
rect 473044 153144 473050 153196
rect 473354 153144 473360 153196
rect 473412 153184 473418 153196
rect 475562 153184 475568 153196
rect 473412 153156 475568 153184
rect 473412 153144 473418 153156
rect 475562 153144 475568 153156
rect 475620 153144 475626 153196
rect 476114 153144 476120 153196
rect 476172 153184 476178 153196
rect 478138 153184 478144 153196
rect 476172 153156 478144 153184
rect 476172 153144 476178 153156
rect 478138 153144 478144 153156
rect 478196 153144 478202 153196
rect 484026 153144 484032 153196
rect 484084 153184 484090 153196
rect 488442 153184 488448 153196
rect 484084 153156 488448 153184
rect 484084 153144 484090 153156
rect 488442 153144 488448 153156
rect 488500 153144 488506 153196
rect 489914 153144 489920 153196
rect 489972 153184 489978 153196
rect 492858 153184 492864 153196
rect 489972 153156 492864 153184
rect 489972 153144 489978 153156
rect 492858 153144 492864 153156
rect 492916 153144 492922 153196
rect 494054 153144 494060 153196
rect 494112 153184 494118 153196
rect 496078 153184 496084 153196
rect 494112 153156 496084 153184
rect 494112 153144 494118 153156
rect 496078 153144 496084 153156
rect 496136 153144 496142 153196
rect 496630 153144 496636 153196
rect 496688 153184 496694 153196
rect 498010 153184 498016 153196
rect 496688 153156 498016 153184
rect 496688 153144 496694 153156
rect 498010 153144 498016 153156
rect 498068 153144 498074 153196
rect 512270 153144 512276 153196
rect 512328 153184 512334 153196
rect 514846 153184 514852 153196
rect 512328 153156 514852 153184
rect 512328 153144 512334 153156
rect 514846 153144 514852 153156
rect 514904 153144 514910 153196
rect 80054 153076 80060 153128
rect 80112 153116 80118 153128
rect 175090 153116 175096 153128
rect 80112 153088 175096 153116
rect 80112 153076 80118 153088
rect 175090 153076 175096 153088
rect 175148 153076 175154 153128
rect 180794 153076 180800 153128
rect 180852 153116 180858 153128
rect 257246 153116 257252 153128
rect 180852 153088 257252 153116
rect 180852 153076 180858 153088
rect 257246 153076 257252 153088
rect 257304 153076 257310 153128
rect 264974 153076 264980 153128
rect 265032 153116 265038 153128
rect 321462 153116 321468 153128
rect 265032 153088 321468 153116
rect 265032 153076 265038 153088
rect 321462 153076 321468 153088
rect 321520 153076 321526 153128
rect 324314 153076 324320 153128
rect 324372 153116 324378 153128
rect 367002 153116 367008 153128
rect 324372 153088 367008 153116
rect 324372 153076 324378 153088
rect 367002 153076 367008 153088
rect 367060 153076 367066 153128
rect 367186 153076 367192 153128
rect 367244 153116 367250 153128
rect 368934 153116 368940 153128
rect 367244 153088 368940 153116
rect 367244 153076 367250 153088
rect 368934 153076 368940 153088
rect 368992 153076 368998 153128
rect 375466 153076 375472 153128
rect 375524 153116 375530 153128
rect 405550 153116 405556 153128
rect 375524 153088 405556 153116
rect 375524 153076 375530 153088
rect 405550 153076 405556 153088
rect 405608 153076 405614 153128
rect 405826 153076 405832 153128
rect 405884 153116 405890 153128
rect 408770 153116 408776 153128
rect 405884 153088 408776 153116
rect 405884 153076 405890 153088
rect 408770 153076 408776 153088
rect 408828 153076 408834 153128
rect 410794 153076 410800 153128
rect 410852 153116 410858 153128
rect 410852 153088 429332 153116
rect 410852 153076 410858 153088
rect 103514 153008 103520 153060
rect 103572 153048 103578 153060
rect 198182 153048 198188 153060
rect 103572 153020 198188 153048
rect 103572 153008 103578 153020
rect 198182 153008 198188 153020
rect 198240 153008 198246 153060
rect 203702 153008 203708 153060
rect 203760 153048 203766 153060
rect 267550 153048 267556 153060
rect 203760 153020 267556 153048
rect 203760 153008 203766 153020
rect 267550 153008 267556 153020
rect 267608 153008 267614 153060
rect 272150 153008 272156 153060
rect 272208 153048 272214 153060
rect 326614 153048 326620 153060
rect 272208 153020 326620 153048
rect 272208 153008 272214 153020
rect 326614 153008 326620 153020
rect 326672 153008 326678 153060
rect 330938 153008 330944 153060
rect 330996 153048 331002 153060
rect 371510 153048 371516 153060
rect 330996 153020 371516 153048
rect 330996 153008 331002 153020
rect 371510 153008 371516 153020
rect 371568 153008 371574 153060
rect 372614 153008 372620 153060
rect 372672 153048 372678 153060
rect 403526 153048 403532 153060
rect 372672 153020 403532 153048
rect 372672 153008 372678 153020
rect 403526 153008 403532 153020
rect 403584 153008 403590 153060
rect 406654 153008 406660 153060
rect 406712 153048 406718 153060
rect 429194 153048 429200 153060
rect 406712 153020 429200 153048
rect 406712 153008 406718 153020
rect 429194 153008 429200 153020
rect 429252 153008 429258 153060
rect 429304 153048 429332 153088
rect 430666 153076 430672 153128
rect 430724 153116 430730 153128
rect 447962 153116 447968 153128
rect 430724 153088 447968 153116
rect 430724 153076 430730 153088
rect 447962 153076 447968 153088
rect 448020 153076 448026 153128
rect 456978 153076 456984 153128
rect 457036 153116 457042 153128
rect 460750 153116 460756 153128
rect 457036 153088 460756 153116
rect 457036 153076 457042 153088
rect 460750 153076 460756 153088
rect 460808 153076 460814 153128
rect 463510 153076 463516 153128
rect 463568 153116 463574 153128
rect 466546 153116 466552 153128
rect 463568 153088 466552 153116
rect 463568 153076 463574 153088
rect 466546 153076 466552 153088
rect 466604 153076 466610 153128
rect 466638 153076 466644 153128
rect 466696 153116 466702 153128
rect 470410 153116 470416 153128
rect 466696 153088 470416 153116
rect 466696 153076 466702 153088
rect 470410 153076 470416 153088
rect 470468 153076 470474 153128
rect 471422 153076 471428 153128
rect 471480 153116 471486 153128
rect 473630 153116 473636 153128
rect 471480 153088 473636 153116
rect 471480 153076 471486 153088
rect 473630 153076 473636 153088
rect 473688 153076 473694 153128
rect 474826 153076 474832 153128
rect 474884 153116 474890 153128
rect 476850 153116 476856 153128
rect 474884 153088 476856 153116
rect 474884 153076 474890 153088
rect 476850 153076 476856 153088
rect 476908 153076 476914 153128
rect 484946 153076 484952 153128
rect 485004 153116 485010 153128
rect 489638 153116 489644 153128
rect 485004 153088 489644 153116
rect 485004 153076 485010 153088
rect 489638 153076 489644 153088
rect 489696 153076 489702 153128
rect 491662 153076 491668 153128
rect 491720 153116 491726 153128
rect 494790 153116 494796 153128
rect 491720 153088 494796 153116
rect 491720 153076 491726 153088
rect 494790 153076 494796 153088
rect 494848 153076 494854 153128
rect 494974 153076 494980 153128
rect 495032 153116 495038 153128
rect 496722 153116 496728 153128
rect 495032 153088 496728 153116
rect 495032 153076 495038 153088
rect 496722 153076 496728 153088
rect 496780 153076 496786 153128
rect 496814 153076 496820 153128
rect 496872 153116 496878 153128
rect 498654 153116 498660 153128
rect 496872 153088 498660 153116
rect 496872 153076 496878 153088
rect 498654 153076 498660 153088
rect 498712 153076 498718 153128
rect 510982 153076 510988 153128
rect 511040 153116 511046 153128
rect 513466 153116 513472 153128
rect 511040 153088 513472 153116
rect 511040 153076 511046 153088
rect 513466 153076 513472 153088
rect 513524 153076 513530 153128
rect 513558 153076 513564 153128
rect 513616 153116 513622 153128
rect 516134 153116 516140 153128
rect 513616 153088 516140 153116
rect 513616 153076 513622 153088
rect 516134 153076 516140 153088
rect 516192 153076 516198 153128
rect 431218 153048 431224 153060
rect 429304 153020 431224 153048
rect 431218 153008 431224 153020
rect 431276 153008 431282 153060
rect 431954 153008 431960 153060
rect 432012 153048 432018 153060
rect 441706 153048 441712 153060
rect 432012 153020 441712 153048
rect 432012 153008 432018 153020
rect 441706 153008 441712 153020
rect 441764 153008 441770 153060
rect 441798 153008 441804 153060
rect 441856 153048 441862 153060
rect 449894 153048 449900 153060
rect 441856 153020 449900 153048
rect 441856 153008 441862 153020
rect 449894 153008 449900 153020
rect 449952 153008 449958 153060
rect 463602 153008 463608 153060
rect 463660 153048 463666 153060
rect 467282 153048 467288 153060
rect 463660 153020 467288 153048
rect 463660 153008 463666 153020
rect 467282 153008 467288 153020
rect 467340 153008 467346 153060
rect 472434 153008 472440 153060
rect 472492 153048 472498 153060
rect 474918 153048 474924 153060
rect 472492 153020 474924 153048
rect 472492 153008 472498 153020
rect 474918 153008 474924 153020
rect 474976 153008 474982 153060
rect 484394 153008 484400 153060
rect 484452 153048 484458 153060
rect 488994 153048 489000 153060
rect 484452 153020 489000 153048
rect 484452 153008 484458 153020
rect 488994 153008 489000 153020
rect 489052 153008 489058 153060
rect 492674 153008 492680 153060
rect 492732 153048 492738 153060
rect 495434 153048 495440 153060
rect 492732 153020 495440 153048
rect 492732 153008 492738 153020
rect 495434 153008 495440 153020
rect 495492 153008 495498 153060
rect 495526 153008 495532 153060
rect 495584 153048 495590 153060
rect 497366 153048 497372 153060
rect 495584 153020 497372 153048
rect 495584 153008 495590 153020
rect 497366 153008 497372 153020
rect 497424 153008 497430 153060
rect 511626 153008 511632 153060
rect 511684 153048 511690 153060
rect 514294 153048 514300 153060
rect 511684 153020 514300 153048
rect 511684 153008 511690 153020
rect 514294 153008 514300 153020
rect 514352 153008 514358 153060
rect 92566 152940 92572 152992
rect 92624 152980 92630 152992
rect 187878 152980 187884 152992
rect 92624 152952 187884 152980
rect 92624 152940 92630 152952
rect 187878 152940 187884 152952
rect 187936 152940 187942 152992
rect 194594 152940 194600 152992
rect 194652 152980 194658 152992
rect 218698 152980 218704 152992
rect 194652 152952 218704 152980
rect 194652 152940 194658 152952
rect 218698 152940 218704 152952
rect 218756 152940 218762 152992
rect 220354 152940 220360 152992
rect 220412 152980 220418 152992
rect 284846 152980 284852 152992
rect 220412 152952 284852 152980
rect 220412 152940 220418 152952
rect 284846 152940 284852 152952
rect 284904 152940 284910 152992
rect 288066 152940 288072 152992
rect 288124 152980 288130 152992
rect 289998 152980 290004 152992
rect 288124 152952 290004 152980
rect 288124 152940 288130 152952
rect 289998 152940 290004 152952
rect 290056 152940 290062 152992
rect 291378 152940 291384 152992
rect 291436 152980 291442 152992
rect 341334 152980 341340 152992
rect 291436 152952 341340 152980
rect 291436 152940 291442 152952
rect 341334 152940 341340 152952
rect 341392 152940 341398 152992
rect 342254 152940 342260 152992
rect 342312 152980 342318 152992
rect 343910 152980 343916 152992
rect 342312 152952 343916 152980
rect 342312 152940 342318 152952
rect 343910 152940 343916 152952
rect 343968 152940 343974 152992
rect 345290 152940 345296 152992
rect 345348 152980 345354 152992
rect 382458 152980 382464 152992
rect 345348 152952 382464 152980
rect 345348 152940 345354 152952
rect 382458 152940 382464 152952
rect 382516 152940 382522 152992
rect 382550 152940 382556 152992
rect 382608 152980 382614 152992
rect 386966 152980 386972 152992
rect 382608 152952 386972 152980
rect 382608 152940 382614 152952
rect 386966 152940 386972 152952
rect 387024 152940 387030 152992
rect 390370 152940 390376 152992
rect 390428 152980 390434 152992
rect 415210 152980 415216 152992
rect 390428 152952 415216 152980
rect 390428 152940 390434 152952
rect 415210 152940 415216 152952
rect 415268 152940 415274 152992
rect 415394 152940 415400 152992
rect 415452 152980 415458 152992
rect 436370 152980 436376 152992
rect 415452 152952 436376 152980
rect 415452 152940 415458 152952
rect 436370 152940 436376 152952
rect 436428 152940 436434 152992
rect 438854 152940 438860 152992
rect 438912 152980 438918 152992
rect 454402 152980 454408 152992
rect 438912 152952 454408 152980
rect 438912 152940 438918 152952
rect 454402 152940 454408 152952
rect 454460 152940 454466 152992
rect 464706 152940 464712 152992
rect 464764 152980 464770 152992
rect 468386 152980 468392 152992
rect 464764 152952 468392 152980
rect 464764 152940 464770 152952
rect 468386 152940 468392 152952
rect 468444 152940 468450 152992
rect 472526 152940 472532 152992
rect 472584 152980 472590 152992
rect 474274 152980 474280 152992
rect 472584 152952 474280 152980
rect 472584 152940 472590 152952
rect 474274 152940 474280 152952
rect 474332 152940 474338 152992
rect 483106 152940 483112 152992
rect 483164 152980 483170 152992
rect 487798 152980 487804 152992
rect 483164 152952 487804 152980
rect 483164 152940 483170 152952
rect 487798 152940 487804 152952
rect 487856 152940 487862 152992
rect 491294 152940 491300 152992
rect 491352 152980 491358 152992
rect 494146 152980 494152 152992
rect 491352 152952 494152 152980
rect 491352 152940 491358 152952
rect 494146 152940 494152 152952
rect 494204 152940 494210 152992
rect 512914 152940 512920 152992
rect 512972 152980 512978 152992
rect 515950 152980 515956 152992
rect 512972 152952 515956 152980
rect 512972 152940 512978 152952
rect 515950 152940 515956 152952
rect 516008 152940 516014 152992
rect 71406 152872 71412 152924
rect 71464 152912 71470 152924
rect 92474 152912 92480 152924
rect 71464 152884 92480 152912
rect 71464 152872 71470 152884
rect 92474 152872 92480 152884
rect 92532 152872 92538 152924
rect 96614 152872 96620 152924
rect 96672 152912 96678 152924
rect 193030 152912 193036 152924
rect 96672 152884 193036 152912
rect 96672 152872 96678 152884
rect 193030 152872 193036 152884
rect 193088 152872 193094 152924
rect 212442 152872 212448 152924
rect 212500 152912 212506 152924
rect 277762 152912 277768 152924
rect 212500 152884 277768 152912
rect 212500 152872 212506 152884
rect 277762 152872 277768 152884
rect 277820 152872 277826 152924
rect 278774 152872 278780 152924
rect 278832 152912 278838 152924
rect 331766 152912 331772 152924
rect 278832 152884 331772 152912
rect 278832 152872 278838 152884
rect 331766 152872 331772 152884
rect 331824 152872 331830 152924
rect 332594 152872 332600 152924
rect 332652 152912 332658 152924
rect 372798 152912 372804 152924
rect 332652 152884 372804 152912
rect 332652 152872 332658 152884
rect 372798 152872 372804 152884
rect 372856 152872 372862 152924
rect 382182 152872 382188 152924
rect 382240 152912 382246 152924
rect 410702 152912 410708 152924
rect 382240 152884 410708 152912
rect 382240 152872 382246 152884
rect 410702 152872 410708 152884
rect 410760 152872 410766 152924
rect 411254 152872 411260 152924
rect 411312 152912 411318 152924
rect 433150 152912 433156 152924
rect 411312 152884 433156 152912
rect 411312 152872 411318 152884
rect 433150 152872 433156 152884
rect 433208 152872 433214 152924
rect 433518 152872 433524 152924
rect 433576 152912 433582 152924
rect 441706 152912 441712 152924
rect 433576 152884 441712 152912
rect 433576 152872 433582 152884
rect 441706 152872 441712 152884
rect 441764 152872 441770 152924
rect 441890 152872 441896 152924
rect 441948 152912 441954 152924
rect 446950 152912 446956 152924
rect 441948 152884 446956 152912
rect 441948 152872 441954 152884
rect 446950 152872 446956 152884
rect 447008 152872 447014 152924
rect 456794 152872 456800 152924
rect 456852 152912 456858 152924
rect 463326 152912 463332 152924
rect 456852 152884 463332 152912
rect 456852 152872 456858 152884
rect 463326 152872 463332 152884
rect 463384 152872 463390 152924
rect 465074 152872 465080 152924
rect 465132 152912 465138 152924
rect 469122 152912 469128 152924
rect 465132 152884 469128 152912
rect 465132 152872 465138 152884
rect 469122 152872 469128 152884
rect 469180 152872 469186 152924
rect 490006 152872 490012 152924
rect 490064 152912 490070 152924
rect 493502 152912 493508 152924
rect 490064 152884 493508 152912
rect 490064 152872 490070 152884
rect 493502 152872 493508 152884
rect 493560 152872 493566 152924
rect 514202 152872 514208 152924
rect 514260 152912 514266 152924
rect 517422 152912 517428 152924
rect 514260 152884 517428 152912
rect 514260 152872 514266 152884
rect 517422 152872 517428 152884
rect 517480 152872 517486 152924
rect 33134 152804 33140 152856
rect 33192 152844 33198 152856
rect 138014 152844 138020 152856
rect 33192 152816 138020 152844
rect 33192 152804 33198 152816
rect 138014 152804 138020 152816
rect 138072 152804 138078 152856
rect 138106 152804 138112 152856
rect 138164 152844 138170 152856
rect 141694 152844 141700 152856
rect 138164 152816 141700 152844
rect 138164 152804 138170 152816
rect 141694 152804 141700 152816
rect 141752 152804 141758 152856
rect 146478 152804 146484 152856
rect 146536 152844 146542 152856
rect 167362 152844 167368 152856
rect 146536 152816 167368 152844
rect 146536 152804 146542 152816
rect 167362 152804 167368 152816
rect 167420 152804 167426 152856
rect 173894 152804 173900 152856
rect 173952 152844 173958 152856
rect 252094 152844 252100 152856
rect 173952 152816 252100 152844
rect 173952 152804 173958 152816
rect 252094 152804 252100 152816
rect 252152 152804 252158 152856
rect 255406 152804 255412 152856
rect 255464 152844 255470 152856
rect 313090 152844 313096 152856
rect 255464 152816 313096 152844
rect 255464 152804 255470 152816
rect 313090 152804 313096 152816
rect 313148 152804 313154 152856
rect 317046 152804 317052 152856
rect 317104 152844 317110 152856
rect 318242 152844 318248 152856
rect 317104 152816 318248 152844
rect 317104 152804 317110 152816
rect 318242 152804 318248 152816
rect 318300 152804 318306 152856
rect 361298 152844 361304 152856
rect 318352 152816 361304 152844
rect 26418 152736 26424 152788
rect 26476 152776 26482 152788
rect 139118 152776 139124 152788
rect 26476 152748 139124 152776
rect 26476 152736 26482 152748
rect 139118 152736 139124 152748
rect 139176 152736 139182 152788
rect 140774 152736 140780 152788
rect 140832 152776 140838 152788
rect 144270 152776 144276 152788
rect 140832 152748 144276 152776
rect 140832 152736 140838 152748
rect 144270 152736 144276 152748
rect 144328 152736 144334 152788
rect 144362 152736 144368 152788
rect 144420 152776 144426 152788
rect 162210 152776 162216 152788
rect 144420 152748 162216 152776
rect 144420 152736 144426 152748
rect 162210 152736 162216 152748
rect 162268 152736 162274 152788
rect 164418 152736 164424 152788
rect 164476 152776 164482 152788
rect 244366 152776 244372 152788
rect 164476 152748 244372 152776
rect 164476 152736 164482 152748
rect 244366 152736 244372 152748
rect 244424 152736 244430 152788
rect 257706 152736 257712 152788
rect 257764 152776 257770 152788
rect 315666 152776 315672 152788
rect 257764 152748 315672 152776
rect 257764 152736 257770 152748
rect 315666 152736 315672 152748
rect 315724 152736 315730 152788
rect 317414 152736 317420 152788
rect 317472 152776 317478 152788
rect 318352 152776 318380 152816
rect 361298 152804 361304 152816
rect 361356 152804 361362 152856
rect 361574 152804 361580 152856
rect 361632 152844 361638 152856
rect 395246 152844 395252 152856
rect 361632 152816 395252 152844
rect 361632 152804 361638 152816
rect 395246 152804 395252 152816
rect 395304 152804 395310 152856
rect 395522 152804 395528 152856
rect 395580 152844 395586 152856
rect 397822 152844 397828 152856
rect 395580 152816 397828 152844
rect 395580 152804 395586 152816
rect 397822 152804 397828 152816
rect 397880 152804 397886 152856
rect 402422 152804 402428 152856
rect 402480 152844 402486 152856
rect 426158 152844 426164 152856
rect 402480 152816 426164 152844
rect 402480 152804 402486 152816
rect 426158 152804 426164 152816
rect 426216 152804 426222 152856
rect 426434 152804 426440 152856
rect 426492 152844 426498 152856
rect 444742 152844 444748 152856
rect 426492 152816 444748 152844
rect 426492 152804 426498 152816
rect 444742 152804 444748 152816
rect 444800 152804 444806 152856
rect 446306 152804 446312 152856
rect 446364 152844 446370 152856
rect 460106 152844 460112 152856
rect 446364 152816 460112 152844
rect 446364 152804 446370 152816
rect 460106 152804 460112 152816
rect 460164 152804 460170 152856
rect 510338 152804 510344 152856
rect 510396 152844 510402 152856
rect 511994 152844 512000 152856
rect 510396 152816 512000 152844
rect 510396 152804 510402 152816
rect 511994 152804 512000 152816
rect 512052 152804 512058 152856
rect 317472 152748 318380 152776
rect 317472 152736 317478 152748
rect 320266 152736 320272 152788
rect 320324 152776 320330 152788
rect 323118 152776 323124 152788
rect 320324 152748 323124 152776
rect 320324 152736 320330 152748
rect 323118 152736 323124 152748
rect 323176 152736 323182 152788
rect 324222 152736 324228 152788
rect 324280 152776 324286 152788
rect 366358 152776 366364 152788
rect 324280 152748 366364 152776
rect 324280 152736 324286 152748
rect 366358 152736 366364 152748
rect 366416 152736 366422 152788
rect 368474 152736 368480 152788
rect 368532 152776 368538 152788
rect 400398 152776 400404 152788
rect 368532 152748 400404 152776
rect 368532 152736 368538 152748
rect 400398 152736 400404 152748
rect 400456 152736 400462 152788
rect 404354 152736 404360 152788
rect 404412 152776 404418 152788
rect 427998 152776 428004 152788
rect 404412 152748 428004 152776
rect 404412 152736 404418 152748
rect 427998 152736 428004 152748
rect 428056 152736 428062 152788
rect 429378 152736 429384 152788
rect 429436 152776 429442 152788
rect 447318 152776 447324 152788
rect 429436 152748 447324 152776
rect 429436 152736 429442 152748
rect 447318 152736 447324 152748
rect 447376 152736 447382 152788
rect 28166 152668 28172 152720
rect 28224 152708 28230 152720
rect 141050 152708 141056 152720
rect 28224 152680 141056 152708
rect 28224 152668 28230 152680
rect 141050 152668 141056 152680
rect 141108 152668 141114 152720
rect 142798 152668 142804 152720
rect 142856 152708 142862 152720
rect 149422 152708 149428 152720
rect 142856 152680 149428 152708
rect 142856 152668 142862 152680
rect 149422 152668 149428 152680
rect 149480 152668 149486 152720
rect 149514 152668 149520 152720
rect 149572 152708 149578 152720
rect 231578 152708 231584 152720
rect 149572 152680 231584 152708
rect 149572 152668 149578 152680
rect 231578 152668 231584 152680
rect 231636 152668 231642 152720
rect 240226 152668 240232 152720
rect 240284 152708 240290 152720
rect 241882 152708 241888 152720
rect 240284 152680 241888 152708
rect 240284 152668 240290 152680
rect 241882 152668 241888 152680
rect 241940 152668 241946 152720
rect 251174 152668 251180 152720
rect 251232 152708 251238 152720
rect 311158 152708 311164 152720
rect 251232 152680 311164 152708
rect 251232 152668 251238 152680
rect 311158 152668 311164 152680
rect 311216 152668 311222 152720
rect 312170 152668 312176 152720
rect 312228 152708 312234 152720
rect 356146 152708 356152 152720
rect 312228 152680 356152 152708
rect 312228 152668 312234 152680
rect 356146 152668 356152 152680
rect 356204 152668 356210 152720
rect 358814 152668 358820 152720
rect 358872 152708 358878 152720
rect 393406 152708 393412 152720
rect 358872 152680 393412 152708
rect 358872 152668 358878 152680
rect 393406 152668 393412 152680
rect 393464 152668 393470 152720
rect 394878 152668 394884 152720
rect 394936 152708 394942 152720
rect 420362 152708 420368 152720
rect 394936 152680 420368 152708
rect 394936 152668 394942 152680
rect 420362 152668 420368 152680
rect 420420 152668 420426 152720
rect 421006 152668 421012 152720
rect 421064 152708 421070 152720
rect 435358 152708 435364 152720
rect 421064 152680 435364 152708
rect 421064 152668 421070 152680
rect 435358 152668 435364 152680
rect 435416 152668 435422 152720
rect 438946 152708 438952 152720
rect 435560 152680 438952 152708
rect 22186 152600 22192 152652
rect 22244 152640 22250 152652
rect 135898 152640 135904 152652
rect 22244 152612 135904 152640
rect 22244 152600 22250 152612
rect 135898 152600 135904 152612
rect 135956 152600 135962 152652
rect 151906 152640 151912 152652
rect 137986 152612 151912 152640
rect 19334 152532 19340 152584
rect 19392 152572 19398 152584
rect 133966 152572 133972 152584
rect 19392 152544 133972 152572
rect 19392 152532 19398 152544
rect 133966 152532 133972 152544
rect 134024 152532 134030 152584
rect 136634 152532 136640 152584
rect 136692 152572 136698 152584
rect 137986 152572 138014 152612
rect 151906 152600 151912 152612
rect 151964 152600 151970 152652
rect 153562 152600 153568 152652
rect 153620 152640 153626 152652
rect 236730 152640 236736 152652
rect 153620 152612 236736 152640
rect 153620 152600 153626 152612
rect 236730 152600 236736 152612
rect 236788 152600 236794 152652
rect 247034 152600 247040 152652
rect 247092 152640 247098 152652
rect 307938 152640 307944 152652
rect 247092 152612 307944 152640
rect 247092 152600 247098 152612
rect 307938 152600 307944 152612
rect 307996 152600 308002 152652
rect 311526 152600 311532 152652
rect 311584 152640 311590 152652
rect 320634 152640 320640 152652
rect 311584 152612 320640 152640
rect 311584 152600 311590 152612
rect 320634 152600 320640 152612
rect 320692 152600 320698 152652
rect 320818 152600 320824 152652
rect 320876 152640 320882 152652
rect 361942 152640 361948 152652
rect 320876 152612 361948 152640
rect 320876 152600 320882 152612
rect 361942 152600 361948 152612
rect 362000 152600 362006 152652
rect 365714 152600 365720 152652
rect 365772 152640 365778 152652
rect 398466 152640 398472 152652
rect 365772 152612 398472 152640
rect 365772 152600 365778 152612
rect 398466 152600 398472 152612
rect 398524 152600 398530 152652
rect 399202 152600 399208 152652
rect 399260 152640 399266 152652
rect 417418 152640 417424 152652
rect 399260 152612 417424 152640
rect 399260 152600 399266 152612
rect 417418 152600 417424 152612
rect 417476 152600 417482 152652
rect 418614 152600 418620 152652
rect 418672 152640 418678 152652
rect 418672 152612 422294 152640
rect 418672 152600 418678 152612
rect 136692 152544 138014 152572
rect 136692 152532 136698 152544
rect 138106 152532 138112 152584
rect 138164 152572 138170 152584
rect 144270 152572 144276 152584
rect 138164 152544 144276 152572
rect 138164 152532 138170 152544
rect 144270 152532 144276 152544
rect 144328 152532 144334 152584
rect 144362 152532 144368 152584
rect 144420 152572 144426 152584
rect 226426 152572 226432 152584
rect 144420 152544 226432 152572
rect 144420 152532 144426 152544
rect 226426 152532 226432 152544
rect 226484 152532 226490 152584
rect 234154 152532 234160 152584
rect 234212 152572 234218 152584
rect 297726 152572 297732 152584
rect 234212 152544 297732 152572
rect 234212 152532 234218 152544
rect 297726 152532 297732 152544
rect 297784 152532 297790 152584
rect 303614 152532 303620 152584
rect 303672 152572 303678 152584
rect 350994 152572 351000 152584
rect 303672 152544 351000 152572
rect 303672 152532 303678 152544
rect 350994 152532 351000 152544
rect 351052 152532 351058 152584
rect 352006 152532 352012 152584
rect 352064 152572 352070 152584
rect 388254 152572 388260 152584
rect 352064 152544 388260 152572
rect 352064 152532 352070 152544
rect 388254 152532 388260 152544
rect 388312 152532 388318 152584
rect 393130 152532 393136 152584
rect 393188 152572 393194 152584
rect 419074 152572 419080 152584
rect 393188 152544 419080 152572
rect 393188 152532 393194 152544
rect 419074 152532 419080 152544
rect 419132 152532 419138 152584
rect 422266 152572 422294 152612
rect 423398 152600 423404 152652
rect 423456 152640 423462 152652
rect 427078 152640 427084 152652
rect 423456 152612 427084 152640
rect 423456 152600 423462 152612
rect 427078 152600 427084 152612
rect 427136 152600 427142 152652
rect 427814 152600 427820 152652
rect 427872 152640 427878 152652
rect 435450 152640 435456 152652
rect 427872 152612 435456 152640
rect 427872 152600 427878 152612
rect 435450 152600 435456 152612
rect 435508 152600 435514 152652
rect 435560 152572 435588 152680
rect 438946 152668 438952 152680
rect 439004 152668 439010 152720
rect 440234 152668 440240 152720
rect 440292 152708 440298 152720
rect 440510 152708 440516 152720
rect 440292 152680 440516 152708
rect 440292 152668 440298 152680
rect 440510 152668 440516 152680
rect 440568 152668 440574 152720
rect 441614 152668 441620 152720
rect 441672 152708 441678 152720
rect 445202 152708 445208 152720
rect 441672 152680 445208 152708
rect 441672 152668 441678 152680
rect 445202 152668 445208 152680
rect 445260 152668 445266 152720
rect 445294 152668 445300 152720
rect 445352 152708 445358 152720
rect 458910 152708 458916 152720
rect 445352 152680 458916 152708
rect 445352 152668 445358 152680
rect 458910 152668 458916 152680
rect 458968 152668 458974 152720
rect 459646 152668 459652 152720
rect 459704 152708 459710 152720
rect 464614 152708 464620 152720
rect 459704 152680 464620 152708
rect 459704 152668 459710 152680
rect 464614 152668 464620 152680
rect 464672 152668 464678 152720
rect 435634 152600 435640 152652
rect 435692 152640 435698 152652
rect 446030 152640 446036 152652
rect 435692 152612 446036 152640
rect 435692 152600 435698 152612
rect 446030 152600 446036 152612
rect 446088 152600 446094 152652
rect 422266 152544 435588 152572
rect 436186 152532 436192 152584
rect 436244 152572 436250 152584
rect 452470 152572 452476 152584
rect 436244 152544 452476 152572
rect 436244 152532 436250 152544
rect 452470 152532 452476 152544
rect 452528 152532 452534 152584
rect 459554 152532 459560 152584
rect 459612 152572 459618 152584
rect 465258 152572 465264 152584
rect 459612 152544 465264 152572
rect 459612 152532 459618 152544
rect 465258 152532 465264 152544
rect 465316 152532 465322 152584
rect 2866 152464 2872 152516
rect 2924 152504 2930 152516
rect 121086 152504 121092 152516
rect 2924 152476 121092 152504
rect 2924 152464 2930 152476
rect 121086 152464 121092 152476
rect 121144 152464 121150 152516
rect 126974 152464 126980 152516
rect 127032 152504 127038 152516
rect 216122 152504 216128 152516
rect 127032 152476 216128 152504
rect 127032 152464 127038 152476
rect 216122 152464 216128 152476
rect 216180 152464 216186 152516
rect 227714 152464 227720 152516
rect 227772 152504 227778 152516
rect 293218 152504 293224 152516
rect 227772 152476 293224 152504
rect 227772 152464 227778 152476
rect 293218 152464 293224 152476
rect 293276 152464 293282 152516
rect 298646 152464 298652 152516
rect 298704 152504 298710 152516
rect 347130 152504 347136 152516
rect 298704 152476 347136 152504
rect 298704 152464 298710 152476
rect 347130 152464 347136 152476
rect 347188 152464 347194 152516
rect 348142 152464 348148 152516
rect 348200 152504 348206 152516
rect 385034 152504 385040 152516
rect 348200 152476 385040 152504
rect 348200 152464 348206 152476
rect 385034 152464 385040 152476
rect 385092 152464 385098 152516
rect 385494 152464 385500 152516
rect 385552 152504 385558 152516
rect 387610 152504 387616 152516
rect 385552 152476 387616 152504
rect 385552 152464 385558 152476
rect 387610 152464 387616 152476
rect 387668 152464 387674 152516
rect 387702 152464 387708 152516
rect 387760 152504 387766 152516
rect 413922 152504 413928 152516
rect 387760 152476 413928 152504
rect 387760 152464 387766 152476
rect 413922 152464 413928 152476
rect 413980 152464 413986 152516
rect 414290 152464 414296 152516
rect 414348 152504 414354 152516
rect 435726 152504 435732 152516
rect 414348 152476 435732 152504
rect 414348 152464 414354 152476
rect 435726 152464 435732 152476
rect 435784 152464 435790 152516
rect 438302 152504 438308 152516
rect 435836 152476 438308 152504
rect 66622 152396 66628 152448
rect 66680 152436 66686 152448
rect 159634 152436 159640 152448
rect 66680 152408 159640 152436
rect 66680 152396 66686 152408
rect 159634 152396 159640 152408
rect 159692 152396 159698 152448
rect 173250 152396 173256 152448
rect 173308 152436 173314 152448
rect 249518 152436 249524 152448
rect 173308 152408 249524 152436
rect 173308 152396 173314 152408
rect 249518 152396 249524 152408
rect 249576 152396 249582 152448
rect 260926 152396 260932 152448
rect 260984 152436 260990 152448
rect 316310 152436 316316 152448
rect 260984 152408 316316 152436
rect 260984 152396 260990 152408
rect 316310 152396 316316 152408
rect 316368 152396 316374 152448
rect 317506 152396 317512 152448
rect 317564 152436 317570 152448
rect 320726 152436 320732 152448
rect 317564 152408 320732 152436
rect 317564 152396 317570 152408
rect 320726 152396 320732 152408
rect 320784 152396 320790 152448
rect 320818 152396 320824 152448
rect 320876 152436 320882 152448
rect 325970 152436 325976 152448
rect 320876 152408 325976 152436
rect 320876 152396 320882 152408
rect 325970 152396 325976 152408
rect 326028 152396 326034 152448
rect 326062 152396 326068 152448
rect 326120 152436 326126 152448
rect 367646 152436 367652 152448
rect 326120 152408 367652 152436
rect 326120 152396 326126 152408
rect 367646 152396 367652 152408
rect 367704 152396 367710 152448
rect 371326 152396 371332 152448
rect 371384 152436 371390 152448
rect 402330 152436 402336 152448
rect 371384 152408 402336 152436
rect 371384 152396 371390 152408
rect 402330 152396 402336 152408
rect 402388 152396 402394 152448
rect 403894 152396 403900 152448
rect 403952 152436 403958 152448
rect 415854 152436 415860 152448
rect 403952 152408 415860 152436
rect 403952 152396 403958 152408
rect 415854 152396 415860 152408
rect 415912 152396 415918 152448
rect 418154 152396 418160 152448
rect 418212 152436 418218 152448
rect 435836 152436 435864 152476
rect 438302 152464 438308 152476
rect 438360 152464 438366 152516
rect 438394 152464 438400 152516
rect 438452 152504 438458 152516
rect 440878 152504 440884 152516
rect 438452 152476 440884 152504
rect 438452 152464 438458 152476
rect 440878 152464 440884 152476
rect 440936 152464 440942 152516
rect 442074 152464 442080 152516
rect 442132 152504 442138 152516
rect 446674 152504 446680 152516
rect 442132 152476 446680 152504
rect 442132 152464 442138 152476
rect 446674 152464 446680 152476
rect 446732 152464 446738 152516
rect 446766 152464 446772 152516
rect 446824 152504 446830 152516
rect 456978 152504 456984 152516
rect 446824 152476 456984 152504
rect 446824 152464 446830 152476
rect 456978 152464 456984 152476
rect 457036 152464 457042 152516
rect 458174 152464 458180 152516
rect 458232 152504 458238 152516
rect 463970 152504 463976 152516
rect 458232 152476 463976 152504
rect 458232 152464 458238 152476
rect 463970 152464 463976 152476
rect 464028 152464 464034 152516
rect 418212 152408 435864 152436
rect 418212 152396 418218 152408
rect 436094 152396 436100 152448
rect 436152 152436 436158 152448
rect 437106 152436 437112 152448
rect 436152 152408 437112 152436
rect 436152 152396 436158 152408
rect 437106 152396 437112 152408
rect 437164 152396 437170 152448
rect 437750 152396 437756 152448
rect 437808 152436 437814 152448
rect 453114 152436 453120 152448
rect 437808 152408 453120 152436
rect 437808 152396 437814 152408
rect 453114 152396 453120 152408
rect 453172 152396 453178 152448
rect 33594 152328 33600 152380
rect 33652 152368 33658 152380
rect 109678 152368 109684 152380
rect 33652 152340 109684 152368
rect 33652 152328 33658 152340
rect 109678 152328 109684 152340
rect 109736 152328 109742 152380
rect 109770 152328 109776 152380
rect 109828 152368 109834 152380
rect 110506 152368 110512 152380
rect 109828 152340 110512 152368
rect 109828 152328 109834 152340
rect 110506 152328 110512 152340
rect 110564 152328 110570 152380
rect 120074 152328 120080 152380
rect 120132 152368 120138 152380
rect 211062 152368 211068 152380
rect 120132 152340 211068 152368
rect 120132 152328 120138 152340
rect 211062 152328 211068 152340
rect 211120 152328 211126 152380
rect 224402 152328 224408 152380
rect 224460 152368 224466 152380
rect 288066 152368 288072 152380
rect 224460 152340 288072 152368
rect 224460 152328 224466 152340
rect 288066 152328 288072 152340
rect 288124 152328 288130 152380
rect 292206 152328 292212 152380
rect 292264 152368 292270 152380
rect 341978 152368 341984 152380
rect 292264 152340 341984 152368
rect 292264 152328 292270 152340
rect 341978 152328 341984 152340
rect 342036 152328 342042 152380
rect 343818 152328 343824 152380
rect 343876 152368 343882 152380
rect 349798 152368 349804 152380
rect 343876 152340 349804 152368
rect 343876 152328 343882 152340
rect 349798 152328 349804 152340
rect 349856 152328 349862 152380
rect 349890 152328 349896 152380
rect 349948 152368 349954 152380
rect 385678 152368 385684 152380
rect 349948 152340 385684 152368
rect 349948 152328 349954 152340
rect 385678 152328 385684 152340
rect 385736 152328 385742 152380
rect 386414 152328 386420 152380
rect 386472 152368 386478 152380
rect 387702 152368 387708 152380
rect 386472 152340 387708 152368
rect 386472 152328 386478 152340
rect 387702 152328 387708 152340
rect 387760 152328 387766 152380
rect 389174 152328 389180 152380
rect 389232 152368 389238 152380
rect 412634 152368 412640 152380
rect 389232 152340 412640 152368
rect 389232 152328 389238 152340
rect 412634 152328 412640 152340
rect 412692 152328 412698 152380
rect 413830 152328 413836 152380
rect 413888 152368 413894 152380
rect 416498 152368 416504 152380
rect 413888 152340 416504 152368
rect 413888 152328 413894 152340
rect 416498 152328 416504 152340
rect 416556 152328 416562 152380
rect 416590 152328 416596 152380
rect 416648 152368 416654 152380
rect 416648 152340 422294 152368
rect 416648 152328 416654 152340
rect 9490 152260 9496 152312
rect 9548 152300 9554 152312
rect 82814 152300 82820 152312
rect 9548 152272 82820 152300
rect 9548 152260 9554 152272
rect 82814 152260 82820 152272
rect 82872 152260 82878 152312
rect 91094 152260 91100 152312
rect 91152 152300 91158 152312
rect 180242 152300 180248 152312
rect 91152 152272 180248 152300
rect 91152 152260 91158 152272
rect 180242 152260 180248 152272
rect 180300 152260 180306 152312
rect 187970 152260 187976 152312
rect 188028 152300 188034 152312
rect 262398 152300 262404 152312
rect 188028 152272 262404 152300
rect 188028 152260 188034 152272
rect 262398 152260 262404 152272
rect 262456 152260 262462 152312
rect 266354 152260 266360 152312
rect 266412 152300 266418 152312
rect 320910 152300 320916 152312
rect 266412 152272 320916 152300
rect 266412 152260 266418 152272
rect 320910 152260 320916 152272
rect 320968 152260 320974 152312
rect 331214 152260 331220 152312
rect 331272 152300 331278 152312
rect 372154 152300 372160 152312
rect 331272 152272 372160 152300
rect 331272 152260 331278 152272
rect 372154 152260 372160 152272
rect 372212 152260 372218 152312
rect 384942 152260 384948 152312
rect 385000 152300 385006 152312
rect 392118 152300 392124 152312
rect 385000 152272 392124 152300
rect 385000 152260 385006 152272
rect 392118 152260 392124 152272
rect 392176 152260 392182 152312
rect 393682 152260 393688 152312
rect 393740 152300 393746 152312
rect 417786 152300 417792 152312
rect 393740 152272 417792 152300
rect 393740 152260 393746 152272
rect 417786 152260 417792 152272
rect 417844 152260 417850 152312
rect 417878 152260 417884 152312
rect 417936 152300 417942 152312
rect 421742 152300 421748 152312
rect 417936 152272 421748 152300
rect 417936 152260 417942 152272
rect 421742 152260 421748 152272
rect 421800 152260 421806 152312
rect 422266 152300 422294 152340
rect 425974 152328 425980 152380
rect 426032 152368 426038 152380
rect 426032 152340 427032 152368
rect 426032 152328 426038 152340
rect 426802 152300 426808 152312
rect 422266 152272 426808 152300
rect 426802 152260 426808 152272
rect 426860 152260 426866 152312
rect 427004 152300 427032 152340
rect 427078 152328 427084 152380
rect 427136 152368 427142 152380
rect 442166 152368 442172 152380
rect 427136 152340 442172 152368
rect 427136 152328 427142 152340
rect 442166 152328 442172 152340
rect 442224 152328 442230 152380
rect 442810 152328 442816 152380
rect 442868 152368 442874 152380
rect 446766 152368 446772 152380
rect 442868 152340 446772 152368
rect 442868 152328 442874 152340
rect 446766 152328 446772 152340
rect 446824 152328 446830 152380
rect 457622 152368 457628 152380
rect 446876 152340 457628 152368
rect 444098 152300 444104 152312
rect 427004 152272 444104 152300
rect 444098 152260 444104 152272
rect 444156 152260 444162 152312
rect 444190 152260 444196 152312
rect 444248 152300 444254 152312
rect 446876 152300 446904 152340
rect 457622 152328 457628 152340
rect 457680 152328 457686 152380
rect 444248 152272 446904 152300
rect 444248 152260 444254 152272
rect 446950 152260 446956 152312
rect 447008 152300 447014 152312
rect 456334 152300 456340 152312
rect 447008 152272 456340 152300
rect 447008 152260 447014 152272
rect 456334 152260 456340 152272
rect 456392 152260 456398 152312
rect 19794 152192 19800 152244
rect 19852 152232 19858 152244
rect 97902 152232 97908 152244
rect 19852 152204 97908 152232
rect 19852 152192 19858 152204
rect 97902 152192 97908 152204
rect 97960 152192 97966 152244
rect 109034 152192 109040 152244
rect 109092 152232 109098 152244
rect 130746 152232 130752 152244
rect 109092 152204 130752 152232
rect 109092 152192 109098 152204
rect 130746 152192 130752 152204
rect 130804 152192 130810 152244
rect 134058 152192 134064 152244
rect 134116 152232 134122 152244
rect 221274 152232 221280 152244
rect 134116 152204 221280 152232
rect 134116 152192 134122 152204
rect 221274 152192 221280 152204
rect 221332 152192 221338 152244
rect 222102 152192 222108 152244
rect 222160 152232 222166 152244
rect 282914 152232 282920 152244
rect 222160 152204 282920 152232
rect 222160 152192 222166 152204
rect 282914 152192 282920 152204
rect 282972 152192 282978 152244
rect 285766 152192 285772 152244
rect 285824 152232 285830 152244
rect 336182 152232 336188 152244
rect 285824 152204 336188 152232
rect 285824 152192 285830 152204
rect 336182 152192 336188 152204
rect 336240 152192 336246 152244
rect 342438 152192 342444 152244
rect 342496 152232 342502 152244
rect 344554 152232 344560 152244
rect 342496 152204 344560 152232
rect 342496 152192 342502 152204
rect 344554 152192 344560 152204
rect 344612 152192 344618 152244
rect 349154 152192 349160 152244
rect 349212 152232 349218 152244
rect 349890 152232 349896 152244
rect 349212 152204 349896 152232
rect 349212 152192 349218 152204
rect 349890 152192 349896 152204
rect 349948 152192 349954 152244
rect 351914 152192 351920 152244
rect 351972 152232 351978 152244
rect 353478 152232 353484 152244
rect 351972 152204 353484 152232
rect 351972 152192 351978 152204
rect 353478 152192 353484 152204
rect 353536 152192 353542 152244
rect 354490 152192 354496 152244
rect 354548 152232 354554 152244
rect 389542 152232 389548 152244
rect 354548 152204 389548 152232
rect 354548 152192 354554 152204
rect 389542 152192 389548 152204
rect 389600 152192 389606 152244
rect 398098 152192 398104 152244
rect 398156 152232 398162 152244
rect 408126 152232 408132 152244
rect 398156 152204 408132 152232
rect 398156 152192 398162 152204
rect 408126 152192 408132 152204
rect 408184 152192 408190 152244
rect 409230 152192 409236 152244
rect 409288 152232 409294 152244
rect 428642 152232 428648 152244
rect 409288 152204 428648 152232
rect 409288 152192 409294 152204
rect 428642 152192 428648 152204
rect 428700 152192 428706 152244
rect 429286 152192 429292 152244
rect 429344 152232 429350 152244
rect 442074 152232 442080 152244
rect 429344 152204 442080 152232
rect 429344 152192 429350 152204
rect 442074 152192 442080 152204
rect 442132 152192 442138 152244
rect 443454 152232 443460 152244
rect 442276 152204 443460 152232
rect 82906 152124 82912 152176
rect 82964 152164 82970 152176
rect 169938 152164 169944 152176
rect 82964 152136 169944 152164
rect 82964 152124 82970 152136
rect 169938 152124 169944 152136
rect 169996 152124 170002 152176
rect 172146 152124 172152 152176
rect 172204 152164 172210 152176
rect 190454 152164 190460 152176
rect 172204 152136 190460 152164
rect 172204 152124 172210 152136
rect 190454 152124 190460 152136
rect 190512 152124 190518 152176
rect 194134 152124 194140 152176
rect 194192 152164 194198 152176
rect 213546 152164 213552 152176
rect 194192 152136 213552 152164
rect 194192 152124 194198 152136
rect 213546 152124 213552 152136
rect 213604 152124 213610 152176
rect 225322 152124 225328 152176
rect 225380 152164 225386 152176
rect 229002 152164 229008 152176
rect 225380 152136 229008 152164
rect 225380 152124 225386 152136
rect 229002 152124 229008 152136
rect 229060 152124 229066 152176
rect 244458 152124 244464 152176
rect 244516 152164 244522 152176
rect 306006 152164 306012 152176
rect 244516 152136 306012 152164
rect 244516 152124 244522 152136
rect 306006 152124 306012 152136
rect 306064 152124 306070 152176
rect 320634 152124 320640 152176
rect 320692 152164 320698 152176
rect 356790 152164 356796 152176
rect 320692 152136 356796 152164
rect 320692 152124 320698 152136
rect 356790 152124 356796 152136
rect 356848 152124 356854 152176
rect 357526 152124 357532 152176
rect 357584 152164 357590 152176
rect 359366 152164 359372 152176
rect 357584 152136 359372 152164
rect 357584 152124 357590 152136
rect 359366 152124 359372 152136
rect 359424 152124 359430 152176
rect 364518 152124 364524 152176
rect 364576 152164 364582 152176
rect 397178 152164 397184 152176
rect 364576 152136 397184 152164
rect 364576 152124 364582 152136
rect 397178 152124 397184 152136
rect 397236 152124 397242 152176
rect 404630 152124 404636 152176
rect 404688 152164 404694 152176
rect 421006 152164 421012 152176
rect 404688 152136 421012 152164
rect 404688 152124 404694 152136
rect 421006 152124 421012 152136
rect 421064 152124 421070 152176
rect 422570 152124 422576 152176
rect 422628 152164 422634 152176
rect 441522 152164 441528 152176
rect 422628 152136 441528 152164
rect 422628 152124 422634 152136
rect 441522 152124 441528 152136
rect 441580 152124 441586 152176
rect 78766 152056 78772 152108
rect 78824 152096 78830 152108
rect 164786 152096 164792 152108
rect 78824 152068 164792 152096
rect 78824 152056 78830 152068
rect 164786 152056 164792 152068
rect 164844 152056 164850 152108
rect 166994 152056 167000 152108
rect 167052 152096 167058 152108
rect 182726 152096 182732 152108
rect 167052 152068 182732 152096
rect 167052 152056 167058 152068
rect 182726 152056 182732 152068
rect 182784 152056 182790 152108
rect 183462 152056 183468 152108
rect 183520 152096 183526 152108
rect 200758 152096 200764 152108
rect 183520 152068 200764 152096
rect 183520 152056 183526 152068
rect 200758 152056 200764 152068
rect 200816 152056 200822 152108
rect 212718 152056 212724 152108
rect 212776 152096 212782 152108
rect 274542 152096 274548 152108
rect 212776 152068 274548 152096
rect 212776 152056 212782 152068
rect 274542 152056 274548 152068
rect 274600 152056 274606 152108
rect 277394 152056 277400 152108
rect 277452 152096 277458 152108
rect 331122 152096 331128 152108
rect 277452 152068 331128 152096
rect 277452 152056 277458 152068
rect 331122 152056 331128 152068
rect 331180 152056 331186 152108
rect 335354 152056 335360 152108
rect 335412 152096 335418 152108
rect 375374 152096 375380 152108
rect 335412 152068 375380 152096
rect 335412 152056 335418 152068
rect 375374 152056 375380 152068
rect 375432 152056 375438 152108
rect 388438 152056 388444 152108
rect 388496 152096 388502 152108
rect 407482 152096 407488 152108
rect 388496 152068 407488 152096
rect 388496 152056 388502 152068
rect 407482 152056 407488 152068
rect 407540 152056 407546 152108
rect 408494 152056 408500 152108
rect 408552 152096 408558 152108
rect 423582 152096 423588 152108
rect 408552 152068 423588 152096
rect 408552 152056 408558 152068
rect 423582 152056 423588 152068
rect 423640 152056 423646 152108
rect 425146 152056 425152 152108
rect 425204 152096 425210 152108
rect 442276 152096 442304 152204
rect 443454 152192 443460 152204
rect 443512 152192 443518 152244
rect 445202 152192 445208 152244
rect 445260 152232 445266 152244
rect 450538 152232 450544 152244
rect 445260 152204 450544 152232
rect 445260 152192 445266 152204
rect 450538 152192 450544 152204
rect 450596 152192 450602 152244
rect 455690 152164 455696 152176
rect 425204 152068 442304 152096
rect 442368 152136 455696 152164
rect 425204 152056 425210 152068
rect 68922 151988 68928 152040
rect 68980 152028 68986 152040
rect 142798 152028 142804 152040
rect 68980 152000 142804 152028
rect 68980 151988 68986 152000
rect 142798 151988 142804 152000
rect 142856 151988 142862 152040
rect 143258 151988 143264 152040
rect 143316 152028 143322 152040
rect 146938 152028 146944 152040
rect 143316 152000 146944 152028
rect 143316 151988 143322 152000
rect 146938 151988 146944 152000
rect 146996 151988 147002 152040
rect 156782 151988 156788 152040
rect 156840 152028 156846 152040
rect 172514 152028 172520 152040
rect 156840 152000 172520 152028
rect 156840 151988 156846 152000
rect 172514 151988 172520 152000
rect 172572 151988 172578 152040
rect 191466 151988 191472 152040
rect 191524 152028 191530 152040
rect 208486 152028 208492 152040
rect 191524 152000 208492 152028
rect 191524 151988 191530 152000
rect 208486 151988 208492 152000
rect 208544 151988 208550 152040
rect 212626 151988 212632 152040
rect 212684 152028 212690 152040
rect 272702 152028 272708 152040
rect 212684 152000 272708 152028
rect 212684 151988 212690 152000
rect 272702 151988 272708 152000
rect 272760 151988 272766 152040
rect 272794 151988 272800 152040
rect 272852 152028 272858 152040
rect 320818 152028 320824 152040
rect 272852 152000 320824 152028
rect 272852 151988 272858 152000
rect 320818 151988 320824 152000
rect 320876 151988 320882 152040
rect 321554 151988 321560 152040
rect 321612 152028 321618 152040
rect 362586 152028 362592 152040
rect 321612 152000 362592 152028
rect 321612 151988 321618 152000
rect 362586 151988 362592 152000
rect 362644 151988 362650 152040
rect 378778 151988 378784 152040
rect 378836 152028 378842 152040
rect 384390 152028 384396 152040
rect 378836 152000 384396 152028
rect 378836 151988 378842 152000
rect 384390 151988 384396 152000
rect 384448 151988 384454 152040
rect 388346 151988 388352 152040
rect 388404 152028 388410 152040
rect 404906 152028 404912 152040
rect 388404 152000 404912 152028
rect 388404 151988 388410 152000
rect 404906 151988 404912 152000
rect 404964 151988 404970 152040
rect 413738 151988 413744 152040
rect 413796 152028 413802 152040
rect 413796 152000 418568 152028
rect 413796 151988 413802 152000
rect 75086 151920 75092 151972
rect 75144 151960 75150 151972
rect 154482 151960 154488 151972
rect 75144 151932 154488 151960
rect 75144 151920 75150 151932
rect 154482 151920 154488 151932
rect 154540 151920 154546 151972
rect 162486 151920 162492 151972
rect 162544 151960 162550 151972
rect 177666 151960 177672 151972
rect 162544 151932 177672 151960
rect 162544 151920 162550 151932
rect 177666 151920 177672 151932
rect 177724 151920 177730 151972
rect 184382 151920 184388 151972
rect 184440 151960 184446 151972
rect 195606 151960 195612 151972
rect 184440 151932 195612 151960
rect 184440 151920 184446 151932
rect 195606 151920 195612 151932
rect 195664 151920 195670 151972
rect 243354 151920 243360 151972
rect 243412 151960 243418 151972
rect 302878 151960 302884 151972
rect 243412 151932 302884 151960
rect 243412 151920 243418 151932
rect 302878 151920 302884 151932
rect 302936 151920 302942 151972
rect 304166 151920 304172 151972
rect 304224 151960 304230 151972
rect 351638 151960 351644 151972
rect 304224 151932 351644 151960
rect 304224 151920 304230 151932
rect 351638 151920 351644 151932
rect 351696 151920 351702 151972
rect 354674 151920 354680 151972
rect 354732 151960 354738 151972
rect 390186 151960 390192 151972
rect 354732 151932 390192 151960
rect 354732 151920 354738 151932
rect 390186 151920 390192 151932
rect 390244 151920 390250 151972
rect 396166 151920 396172 151972
rect 396224 151960 396230 151972
rect 402974 151960 402980 151972
rect 396224 151932 402980 151960
rect 396224 151920 396230 151932
rect 402974 151920 402980 151932
rect 403032 151920 403038 151972
rect 404262 151920 404268 151972
rect 404320 151960 404326 151972
rect 418430 151960 418436 151972
rect 404320 151932 418436 151960
rect 404320 151920 404326 151932
rect 418430 151920 418436 151932
rect 418488 151920 418494 151972
rect 418540 151960 418568 152000
rect 419534 151988 419540 152040
rect 419592 152028 419598 152040
rect 437014 152028 437020 152040
rect 419592 152000 437020 152028
rect 419592 151988 419598 152000
rect 437014 151988 437020 152000
rect 437072 151988 437078 152040
rect 437106 151988 437112 152040
rect 437164 152028 437170 152040
rect 440234 152028 440240 152040
rect 437164 152000 440240 152028
rect 437164 151988 437170 152000
rect 440234 151988 440240 152000
rect 440292 151988 440298 152040
rect 440326 151988 440332 152040
rect 440384 152028 440390 152040
rect 442368 152028 442396 152136
rect 455690 152124 455696 152136
rect 455748 152124 455754 152176
rect 440384 152000 442396 152028
rect 443380 152068 443684 152096
rect 440384 151988 440390 152000
rect 421650 151960 421656 151972
rect 418540 151932 421656 151960
rect 421650 151920 421656 151932
rect 421708 151920 421714 151972
rect 421742 151920 421748 151972
rect 421800 151960 421806 151972
rect 422846 151960 422852 151972
rect 421800 151932 422852 151960
rect 421800 151920 421806 151932
rect 422846 151920 422852 151932
rect 422904 151920 422910 151972
rect 423490 151920 423496 151972
rect 423548 151960 423554 151972
rect 439590 151960 439596 151972
rect 423548 151932 439596 151960
rect 423548 151920 423554 151932
rect 439590 151920 439596 151932
rect 439648 151920 439654 151972
rect 440510 151920 440516 151972
rect 440568 151960 440574 151972
rect 443380 151960 443408 152068
rect 440568 151932 443408 151960
rect 443656 151960 443684 152068
rect 444466 152056 444472 152108
rect 444524 152096 444530 152108
rect 458174 152096 458180 152108
rect 444524 152068 458180 152096
rect 444524 152056 444530 152068
rect 458174 152056 458180 152068
rect 458232 152056 458238 152108
rect 516686 152056 516692 152108
rect 516744 152096 516750 152108
rect 520274 152096 520280 152108
rect 516744 152068 520280 152096
rect 516744 152056 516750 152068
rect 520274 152056 520280 152068
rect 520332 152056 520338 152108
rect 443730 151988 443736 152040
rect 443788 152028 443794 152040
rect 453758 152028 453764 152040
rect 443788 152000 453764 152028
rect 443788 151988 443794 152000
rect 453758 151988 453764 152000
rect 453816 151988 453822 152040
rect 456886 151988 456892 152040
rect 456944 152028 456950 152040
rect 462682 152028 462688 152040
rect 456944 152000 462688 152028
rect 456944 151988 456950 152000
rect 462682 151988 462688 152000
rect 462740 151988 462746 152040
rect 485774 151988 485780 152040
rect 485832 152028 485838 152040
rect 490282 152028 490288 152040
rect 485832 152000 490288 152028
rect 485832 151988 485838 152000
rect 490282 151988 490288 152000
rect 490340 151988 490346 152040
rect 455046 151960 455052 151972
rect 443656 151932 455052 151960
rect 440568 151920 440574 151932
rect 455046 151920 455052 151932
rect 455104 151920 455110 151972
rect 456058 151920 456064 151972
rect 456116 151960 456122 151972
rect 461394 151960 461400 151972
rect 456116 151932 461400 151960
rect 456116 151920 456122 151932
rect 461394 151920 461400 151932
rect 461452 151920 461458 151972
rect 469214 151920 469220 151972
rect 469272 151960 469278 151972
rect 472342 151960 472348 151972
rect 469272 151932 472348 151960
rect 469272 151920 469278 151932
rect 472342 151920 472348 151932
rect 472400 151920 472406 151972
rect 487338 151920 487344 151972
rect 487396 151960 487402 151972
rect 490926 151960 490932 151972
rect 487396 151932 490932 151960
rect 487396 151920 487402 151932
rect 490926 151920 490932 151932
rect 490984 151920 490990 151972
rect 509050 151920 509056 151972
rect 509108 151960 509114 151972
rect 510890 151960 510896 151972
rect 509108 151932 510896 151960
rect 509108 151920 509114 151932
rect 510890 151920 510896 151932
rect 510948 151920 510954 151972
rect 517422 151920 517428 151972
rect 517480 151960 517486 151972
rect 521562 151960 521568 151972
rect 517480 151932 521568 151960
rect 517480 151920 517486 151932
rect 521562 151920 521568 151932
rect 521620 151920 521626 151972
rect 30190 151852 30196 151904
rect 30248 151892 30254 151904
rect 110322 151892 110328 151904
rect 30248 151864 110328 151892
rect 30248 151852 30254 151864
rect 110322 151852 110328 151864
rect 110380 151852 110386 151904
rect 110506 151852 110512 151904
rect 110564 151892 110570 151904
rect 138474 151892 138480 151904
rect 110564 151864 138480 151892
rect 110564 151852 110570 151864
rect 138474 151852 138480 151864
rect 138532 151852 138538 151904
rect 139302 151852 139308 151904
rect 139360 151892 139366 151904
rect 203334 151892 203340 151904
rect 139360 151864 203340 151892
rect 139360 151852 139366 151864
rect 203334 151852 203340 151864
rect 203392 151852 203398 151904
rect 241606 151852 241612 151904
rect 241664 151892 241670 151904
rect 300946 151892 300952 151904
rect 241664 151864 300952 151892
rect 241664 151852 241670 151864
rect 300946 151852 300952 151864
rect 301004 151852 301010 151904
rect 307386 151852 307392 151904
rect 307444 151892 307450 151904
rect 352282 151892 352288 151904
rect 307444 151864 352288 151892
rect 307444 151852 307450 151864
rect 352282 151852 352288 151864
rect 352340 151852 352346 151904
rect 363138 151852 363144 151904
rect 363196 151892 363202 151904
rect 364518 151892 364524 151904
rect 363196 151864 364524 151892
rect 363196 151852 363202 151864
rect 364518 151852 364524 151864
rect 364576 151852 364582 151904
rect 386138 151852 386144 151904
rect 386196 151892 386202 151904
rect 399754 151892 399760 151904
rect 386196 151864 399760 151892
rect 386196 151852 386202 151864
rect 399754 151852 399760 151864
rect 399812 151852 399818 151904
rect 417418 151852 417424 151904
rect 417476 151892 417482 151904
rect 424134 151892 424140 151904
rect 417476 151864 424140 151892
rect 417476 151852 417482 151864
rect 424134 151852 424140 151864
rect 424192 151852 424198 151904
rect 434438 151892 434444 151904
rect 424244 151864 434444 151892
rect 74810 151784 74816 151836
rect 74868 151824 74874 151836
rect 81342 151824 81348 151836
rect 74868 151796 81348 151824
rect 74868 151784 74874 151796
rect 81342 151784 81348 151796
rect 81400 151784 81406 151836
rect 105814 151784 105820 151836
rect 105872 151824 105878 151836
rect 110230 151824 110236 151836
rect 105872 151796 110236 151824
rect 105872 151784 105878 151796
rect 110230 151784 110236 151796
rect 110288 151784 110294 151836
rect 110414 151784 110420 151836
rect 110472 151824 110478 151836
rect 128170 151824 128176 151836
rect 110472 151796 128176 151824
rect 110472 151784 110478 151796
rect 128170 151784 128176 151796
rect 128228 151784 128234 151836
rect 129734 151784 129740 151836
rect 129792 151824 129798 151836
rect 146846 151824 146852 151836
rect 129792 151796 146852 151824
rect 129792 151784 129798 151796
rect 146846 151784 146852 151796
rect 146904 151784 146910 151836
rect 146938 151784 146944 151836
rect 146996 151824 147002 151836
rect 157058 151824 157064 151836
rect 146996 151796 157064 151824
rect 146996 151784 147002 151796
rect 157058 151784 157064 151796
rect 157116 151784 157122 151836
rect 169754 151784 169760 151836
rect 169812 151824 169818 151836
rect 185302 151824 185308 151836
rect 169812 151796 185308 151824
rect 169812 151784 169818 151796
rect 185302 151784 185308 151796
rect 185360 151784 185366 151836
rect 283190 151784 283196 151836
rect 283248 151824 283254 151836
rect 287422 151824 287428 151836
rect 283248 151796 287428 151824
rect 283248 151784 283254 151796
rect 287422 151784 287428 151796
rect 287480 151784 287486 151836
rect 300394 151784 300400 151836
rect 300452 151824 300458 151836
rect 346486 151824 346492 151836
rect 300452 151796 342852 151824
rect 300452 151784 300458 151796
rect 102318 151716 102324 151768
rect 102376 151756 102382 151768
rect 116118 151756 116124 151768
rect 102376 151728 116124 151756
rect 102376 151716 102382 151728
rect 116118 151716 116124 151728
rect 116176 151716 116182 151768
rect 342824 151756 342852 151796
rect 344020 151796 346492 151824
rect 344020 151756 344048 151796
rect 346486 151784 346492 151796
rect 346544 151784 346550 151836
rect 349798 151784 349804 151836
rect 349856 151824 349862 151836
rect 380526 151824 380532 151836
rect 349856 151796 380532 151824
rect 349856 151784 349862 151796
rect 380526 151784 380532 151796
rect 380584 151784 380590 151836
rect 386230 151784 386236 151836
rect 386288 151824 386294 151836
rect 394694 151824 394700 151836
rect 386288 151796 394700 151824
rect 386288 151784 386294 151796
rect 394694 151784 394700 151796
rect 394752 151784 394758 151836
rect 398834 151784 398840 151836
rect 398892 151824 398898 151836
rect 413278 151824 413284 151836
rect 398892 151796 413284 151824
rect 398892 151784 398898 151796
rect 413278 151784 413284 151796
rect 413336 151784 413342 151836
rect 419626 151784 419632 151836
rect 419684 151824 419690 151836
rect 424244 151824 424272 151864
rect 434438 151852 434444 151864
rect 434496 151852 434502 151904
rect 435358 151852 435364 151904
rect 435416 151892 435422 151904
rect 438394 151892 438400 151904
rect 435416 151864 438400 151892
rect 435416 151852 435422 151864
rect 438394 151852 438400 151864
rect 438452 151852 438458 151904
rect 438578 151852 438584 151904
rect 438636 151892 438642 151904
rect 443546 151892 443552 151904
rect 438636 151864 443552 151892
rect 438636 151852 438642 151864
rect 443546 151852 443552 151864
rect 443604 151852 443610 151904
rect 451826 151892 451832 151904
rect 443656 151864 451832 151892
rect 431770 151824 431776 151836
rect 419684 151796 424272 151824
rect 424336 151796 431776 151824
rect 419684 151784 419690 151796
rect 342824 151728 344048 151756
rect 422846 151716 422852 151768
rect 422904 151756 422910 151768
rect 424336 151756 424364 151796
rect 431770 151784 431776 151796
rect 431828 151784 431834 151836
rect 434714 151784 434720 151836
rect 434772 151824 434778 151836
rect 440050 151824 440056 151836
rect 434772 151796 440056 151824
rect 434772 151784 434778 151796
rect 440050 151784 440056 151796
rect 440108 151784 440114 151836
rect 440234 151784 440240 151836
rect 440292 151824 440298 151836
rect 443656 151824 443684 151864
rect 451826 151852 451832 151864
rect 451884 151852 451890 151904
rect 467834 151852 467840 151904
rect 467892 151892 467898 151904
rect 471054 151892 471060 151904
rect 467892 151864 471060 151892
rect 467892 151852 467898 151864
rect 471054 151852 471060 151864
rect 471112 151852 471118 151904
rect 488534 151852 488540 151904
rect 488592 151892 488598 151904
rect 492214 151892 492220 151904
rect 488592 151864 492220 151892
rect 488592 151852 488598 151864
rect 492214 151852 492220 151864
rect 492272 151852 492278 151904
rect 507762 151852 507768 151904
rect 507820 151892 507826 151904
rect 509510 151892 509516 151904
rect 507820 151864 509516 151892
rect 507820 151852 507826 151864
rect 509510 151852 509516 151864
rect 509568 151852 509574 151904
rect 516042 151852 516048 151904
rect 516100 151892 516106 151904
rect 519446 151892 519452 151904
rect 516100 151864 519452 151892
rect 516100 151852 516106 151864
rect 519446 151852 519452 151864
rect 519504 151852 519510 151904
rect 451090 151824 451096 151836
rect 440292 151796 443684 151824
rect 443748 151796 451096 151824
rect 440292 151784 440298 151796
rect 443748 151756 443776 151796
rect 451090 151784 451096 151796
rect 451148 151784 451154 151836
rect 456150 151784 456156 151836
rect 456208 151824 456214 151836
rect 462038 151824 462044 151836
rect 456208 151796 462044 151824
rect 456208 151784 456214 151796
rect 462038 151784 462044 151796
rect 462096 151784 462102 151836
rect 463878 151784 463884 151836
rect 463936 151824 463942 151836
rect 467742 151824 467748 151836
rect 463936 151796 467748 151824
rect 463936 151784 463942 151796
rect 467742 151784 467748 151796
rect 467800 151784 467806 151836
rect 467926 151784 467932 151836
rect 467984 151824 467990 151836
rect 471698 151824 471704 151836
rect 467984 151796 471704 151824
rect 467984 151784 467990 151796
rect 471698 151784 471704 151796
rect 471756 151784 471762 151836
rect 488166 151784 488172 151836
rect 488224 151824 488230 151836
rect 491570 151824 491576 151836
rect 488224 151796 491576 151824
rect 488224 151784 488230 151796
rect 491570 151784 491576 151796
rect 491628 151784 491634 151836
rect 499114 151784 499120 151836
rect 499172 151824 499178 151836
rect 499942 151824 499948 151836
rect 499172 151796 499948 151824
rect 499172 151784 499178 151796
rect 499942 151784 499948 151796
rect 500000 151784 500006 151836
rect 515490 151784 515496 151836
rect 515548 151824 515554 151836
rect 518894 151824 518900 151836
rect 515548 151796 518900 151824
rect 515548 151784 515554 151796
rect 518894 151784 518900 151796
rect 518952 151784 518958 151836
rect 422904 151728 424364 151756
rect 441586 151728 443776 151756
rect 422904 151716 422910 151728
rect 98914 151648 98920 151700
rect 98972 151688 98978 151700
rect 116026 151688 116032 151700
rect 98972 151660 116032 151688
rect 98972 151648 98978 151660
rect 116026 151648 116032 151660
rect 116084 151648 116090 151700
rect 440142 151648 440148 151700
rect 440200 151688 440206 151700
rect 441586 151688 441614 151728
rect 440200 151660 441614 151688
rect 440200 151648 440206 151660
rect 40494 151580 40500 151632
rect 40552 151620 40558 151632
rect 110966 151620 110972 151632
rect 40552 151592 110972 151620
rect 40552 151580 40558 151592
rect 110966 151580 110972 151592
rect 111024 151580 111030 151632
rect 92014 151512 92020 151564
rect 92072 151552 92078 151564
rect 113082 151552 113088 151564
rect 92072 151524 113088 151552
rect 92072 151512 92078 151524
rect 113082 151512 113088 151524
rect 113140 151512 113146 151564
rect 26694 151444 26700 151496
rect 26752 151484 26758 151496
rect 116946 151484 116952 151496
rect 26752 151456 116952 151484
rect 26752 151444 26758 151456
rect 116946 151444 116952 151456
rect 117004 151444 117010 151496
rect 16390 151376 16396 151428
rect 16448 151416 16454 151428
rect 116762 151416 116768 151428
rect 16448 151388 116768 151416
rect 16448 151376 16454 151388
rect 116762 151376 116768 151388
rect 116820 151376 116826 151428
rect 12986 151308 12992 151360
rect 13044 151348 13050 151360
rect 116670 151348 116676 151360
rect 13044 151320 116676 151348
rect 13044 151308 13050 151320
rect 116670 151308 116676 151320
rect 116728 151308 116734 151360
rect 68002 151240 68008 151292
rect 68060 151280 68066 151292
rect 112714 151280 112720 151292
rect 68060 151252 112720 151280
rect 68060 151240 68066 151252
rect 112714 151240 112720 151252
rect 112772 151240 112778 151292
rect 64506 151172 64512 151224
rect 64564 151212 64570 151224
rect 112622 151212 112628 151224
rect 64564 151184 112628 151212
rect 64564 151172 64570 151184
rect 112622 151172 112628 151184
rect 112680 151172 112686 151224
rect 61102 151104 61108 151156
rect 61160 151144 61166 151156
rect 112530 151144 112536 151156
rect 61160 151116 112536 151144
rect 61160 151104 61166 151116
rect 112530 151104 112536 151116
rect 112588 151104 112594 151156
rect 57698 151036 57704 151088
rect 57756 151076 57762 151088
rect 111702 151076 111708 151088
rect 57756 151048 111708 151076
rect 57756 151036 57762 151048
rect 111702 151036 111708 151048
rect 111760 151036 111766 151088
rect 54202 150968 54208 151020
rect 54260 151008 54266 151020
rect 112438 151008 112444 151020
rect 54260 150980 112444 151008
rect 54260 150968 54266 150980
rect 112438 150968 112444 150980
rect 112496 150968 112502 151020
rect 50798 150900 50804 150952
rect 50856 150940 50862 150952
rect 111610 150940 111616 150952
rect 50856 150912 111616 150940
rect 50856 150900 50862 150912
rect 111610 150900 111616 150912
rect 111668 150900 111674 150952
rect 47302 150832 47308 150884
rect 47360 150872 47366 150884
rect 111518 150872 111524 150884
rect 47360 150844 111524 150872
rect 47360 150832 47366 150844
rect 111518 150832 111524 150844
rect 111576 150832 111582 150884
rect 43898 150764 43904 150816
rect 43956 150804 43962 150816
rect 111426 150804 111432 150816
rect 43956 150776 111432 150804
rect 43956 150764 43962 150776
rect 111426 150764 111432 150776
rect 111484 150764 111490 150816
rect 95510 150696 95516 150748
rect 95568 150736 95574 150748
rect 115290 150736 115296 150748
rect 95568 150708 115296 150736
rect 95568 150696 95574 150708
rect 115290 150696 115296 150708
rect 115348 150696 115354 150748
rect 36998 150628 37004 150680
rect 37056 150668 37062 150680
rect 111242 150668 111248 150680
rect 37056 150640 111248 150668
rect 37056 150628 37062 150640
rect 111242 150628 111248 150640
rect 111300 150628 111306 150680
rect 88610 150560 88616 150612
rect 88668 150600 88674 150612
rect 112990 150600 112996 150612
rect 88668 150572 112996 150600
rect 88668 150560 88674 150572
rect 112990 150560 112996 150572
rect 113048 150560 113054 150612
rect 85206 150492 85212 150544
rect 85264 150532 85270 150544
rect 115198 150532 115204 150544
rect 85264 150504 115204 150532
rect 85264 150492 85270 150504
rect 115198 150492 115204 150504
rect 115256 150492 115262 150544
rect 81710 150424 81716 150476
rect 81768 150464 81774 150476
rect 112898 150464 112904 150476
rect 81768 150436 112904 150464
rect 81768 150424 81774 150436
rect 112898 150424 112904 150436
rect 112956 150424 112962 150476
rect 78306 150288 78312 150340
rect 78364 150328 78370 150340
rect 112806 150328 112812 150340
rect 78364 150300 112812 150328
rect 78364 150288 78370 150300
rect 112806 150288 112812 150300
rect 112864 150288 112870 150340
rect 263686 150288 263692 150340
rect 263744 150328 263750 150340
rect 263744 150300 264422 150328
rect 263744 150288 263750 150300
rect 110322 150220 110328 150272
rect 110380 150260 110386 150272
rect 117130 150260 117136 150272
rect 110380 150232 117136 150260
rect 110380 150220 110386 150232
rect 117130 150220 117136 150232
rect 117188 150220 117194 150272
rect 264394 150204 264422 150300
rect 97902 150152 97908 150204
rect 97960 150192 97966 150204
rect 116854 150192 116860 150204
rect 97960 150164 116860 150192
rect 97960 150152 97966 150164
rect 116854 150152 116860 150164
rect 116912 150152 116918 150204
rect 122834 150152 122840 150204
rect 122892 150192 122898 150204
rect 123708 150192 123714 150204
rect 122892 150164 123714 150192
rect 122892 150152 122898 150164
rect 123708 150152 123714 150164
rect 123766 150152 123772 150204
rect 136910 150152 136916 150204
rect 136968 150192 136974 150204
rect 139808 150192 139814 150204
rect 136968 150164 139814 150192
rect 136968 150152 136974 150164
rect 139808 150152 139814 150164
rect 139866 150152 139872 150204
rect 146386 150152 146392 150204
rect 146444 150192 146450 150204
rect 147536 150192 147542 150204
rect 146444 150164 147542 150192
rect 146444 150152 146450 150164
rect 147536 150152 147542 150164
rect 147594 150152 147600 150204
rect 147674 150152 147680 150204
rect 147732 150192 147738 150204
rect 148824 150192 148830 150204
rect 147732 150164 148830 150192
rect 147732 150152 147738 150164
rect 148824 150152 148830 150164
rect 148882 150152 148888 150204
rect 164326 150152 164332 150204
rect 164384 150192 164390 150204
rect 165476 150192 165482 150204
rect 164384 150164 165482 150192
rect 164384 150152 164390 150164
rect 165476 150152 165482 150164
rect 165534 150152 165540 150204
rect 168466 150152 168472 150204
rect 168524 150192 168530 150204
rect 169340 150192 169346 150204
rect 168524 150164 169346 150192
rect 168524 150152 168530 150164
rect 169340 150152 169346 150164
rect 169398 150152 169404 150204
rect 171134 150152 171140 150204
rect 171192 150192 171198 150204
rect 171916 150192 171922 150204
rect 171192 150164 171922 150192
rect 171192 150152 171198 150164
rect 171916 150152 171922 150164
rect 171974 150152 171980 150204
rect 172698 150152 172704 150204
rect 172756 150192 172762 150204
rect 173848 150192 173854 150204
rect 172756 150164 173854 150192
rect 172756 150152 172762 150164
rect 173848 150152 173854 150164
rect 173906 150152 173912 150204
rect 182266 150152 182272 150204
rect 182324 150192 182330 150204
rect 183416 150192 183422 150204
rect 182324 150164 183422 150192
rect 182324 150152 182330 150164
rect 183416 150152 183422 150164
rect 183474 150152 183480 150204
rect 196526 150152 196532 150204
rect 196584 150192 196590 150204
rect 199516 150192 199522 150204
rect 196584 150164 199522 150192
rect 196584 150152 196590 150164
rect 199516 150152 199522 150164
rect 199574 150152 199580 150204
rect 225046 150152 225052 150204
rect 225104 150192 225110 150204
rect 225828 150192 225834 150204
rect 225104 150164 225834 150192
rect 225104 150152 225110 150164
rect 225828 150152 225834 150164
rect 225886 150152 225892 150204
rect 229186 150152 229192 150204
rect 229244 150192 229250 150204
rect 230336 150192 230342 150204
rect 229244 150164 230342 150192
rect 229244 150152 229250 150164
rect 230336 150152 230342 150164
rect 230394 150152 230400 150204
rect 233234 150152 233240 150204
rect 233292 150192 233298 150204
rect 234200 150192 234206 150204
rect 233292 150164 234206 150192
rect 233292 150152 233298 150164
rect 234200 150152 234206 150164
rect 234258 150152 234264 150204
rect 238938 150152 238944 150204
rect 238996 150192 239002 150204
rect 239996 150192 240002 150204
rect 238996 150164 240002 150192
rect 238996 150152 239002 150164
rect 239996 150152 240002 150164
rect 240054 150152 240060 150204
rect 253934 150152 253940 150204
rect 253992 150192 253998 150204
rect 254716 150192 254722 150204
rect 253992 150164 254722 150192
rect 253992 150152 253998 150164
rect 254716 150152 254722 150164
rect 254774 150152 254780 150204
rect 256786 150152 256792 150204
rect 256844 150192 256850 150204
rect 257936 150192 257942 150204
rect 256844 150164 257942 150192
rect 256844 150152 256850 150164
rect 257936 150152 257942 150164
rect 257994 150152 258000 150204
rect 264376 150152 264382 150204
rect 264434 150152 264440 150204
rect 269114 150152 269120 150204
rect 269172 150192 269178 150204
rect 270172 150192 270178 150204
rect 269172 150164 270178 150192
rect 269172 150152 269178 150164
rect 270172 150152 270178 150164
rect 270230 150152 270236 150204
rect 283098 150152 283104 150204
rect 283156 150192 283162 150204
rect 284248 150192 284254 150204
rect 283156 150164 284254 150192
rect 283156 150152 283162 150164
rect 284248 150152 284254 150164
rect 284306 150152 284312 150204
rect 284386 150152 284392 150204
rect 284444 150192 284450 150204
rect 285536 150192 285542 150204
rect 284444 150164 285542 150192
rect 284444 150152 284450 150164
rect 285536 150152 285542 150164
rect 285594 150152 285600 150204
rect 299474 150152 299480 150204
rect 299532 150192 299538 150204
rect 300348 150192 300354 150204
rect 299532 150164 300354 150192
rect 299532 150152 299538 150164
rect 300348 150152 300354 150164
rect 300406 150152 300412 150204
rect 328454 150152 328460 150204
rect 328512 150192 328518 150204
rect 329236 150192 329242 150204
rect 328512 150164 329242 150192
rect 328512 150152 328518 150164
rect 329236 150152 329242 150164
rect 329294 150152 329300 150204
rect 332686 150152 332692 150204
rect 332744 150192 332750 150204
rect 333744 150192 333750 150204
rect 332744 150164 333750 150192
rect 332744 150152 332750 150164
rect 333744 150152 333750 150164
rect 333802 150152 333808 150204
rect 338390 150152 338396 150204
rect 338448 150192 338454 150204
rect 339448 150192 339454 150204
rect 338448 150164 339454 150192
rect 338448 150152 338454 150164
rect 339448 150152 339454 150164
rect 339506 150152 339512 150204
rect 345106 150152 345112 150204
rect 345164 150192 345170 150204
rect 345888 150192 345894 150204
rect 345164 150164 345894 150192
rect 345164 150152 345170 150164
rect 345888 150152 345894 150164
rect 345946 150152 345952 150204
rect 358906 150152 358912 150204
rect 358964 150192 358970 150204
rect 360056 150192 360062 150204
rect 358964 150164 360062 150192
rect 358964 150152 358970 150164
rect 360056 150152 360062 150164
rect 360114 150152 360120 150204
rect 362954 150152 362960 150204
rect 363012 150192 363018 150204
rect 363920 150192 363926 150204
rect 363012 150164 363926 150192
rect 363012 150152 363018 150164
rect 363920 150152 363926 150164
rect 363978 150152 363984 150204
rect 375558 150152 375564 150204
rect 375616 150192 375622 150204
rect 376708 150192 376714 150204
rect 375616 150164 376714 150192
rect 375616 150152 375622 150164
rect 376708 150152 376714 150164
rect 376766 150152 376772 150204
rect 378134 150152 378140 150204
rect 378192 150192 378198 150204
rect 379284 150192 379290 150204
rect 378192 150164 379290 150192
rect 378192 150152 378198 150164
rect 379284 150152 379290 150164
rect 379342 150152 379348 150204
rect 394970 150152 394976 150204
rect 395028 150192 395034 150204
rect 396028 150192 396034 150204
rect 395028 150164 396034 150192
rect 395028 150152 395034 150164
rect 396028 150152 396034 150164
rect 396086 150152 396092 150204
rect 403158 150152 403164 150204
rect 403216 150192 403222 150204
rect 404308 150192 404314 150204
rect 403216 150164 404314 150192
rect 403216 150152 403222 150164
rect 404308 150152 404314 150164
rect 404366 150152 404372 150204
rect 477678 150152 477684 150204
rect 477736 150192 477742 150204
rect 478828 150192 478834 150204
rect 477736 150164 478834 150192
rect 477736 150152 477742 150164
rect 478828 150152 478834 150164
rect 478886 150152 478892 150204
rect 478966 150152 478972 150204
rect 479024 150192 479030 150204
rect 480116 150192 480122 150204
rect 479024 150164 480122 150192
rect 479024 150152 479030 150164
rect 480116 150152 480122 150164
rect 480174 150152 480180 150204
rect 480254 150152 480260 150204
rect 480312 150192 480318 150204
rect 481404 150192 481410 150204
rect 480312 150164 481410 150192
rect 480312 150152 480318 150164
rect 481404 150152 481410 150164
rect 481462 150152 481468 150204
rect 483198 150152 483204 150204
rect 483256 150192 483262 150204
rect 483980 150192 483986 150204
rect 483256 150164 483986 150192
rect 483256 150152 483262 150164
rect 483980 150152 483986 150164
rect 484038 150152 484044 150204
rect 502334 150152 502340 150204
rect 502392 150192 502398 150204
rect 503208 150192 503214 150204
rect 502392 150164 503214 150192
rect 502392 150152 502398 150164
rect 503208 150152 503214 150164
rect 503266 150152 503272 150204
rect 518020 150152 518026 150204
rect 518078 150192 518084 150204
rect 518802 150192 518808 150204
rect 518078 150164 518808 150192
rect 518078 150152 518084 150164
rect 518802 150152 518808 150164
rect 518860 150152 518866 150204
rect 81342 150084 81348 150136
rect 81400 150124 81406 150136
rect 81400 150096 84194 150124
rect 81400 150084 81406 150096
rect 84166 150056 84194 150096
rect 92474 150084 92480 150136
rect 92532 150124 92538 150136
rect 117222 150124 117228 150136
rect 92532 150096 117228 150124
rect 92532 150084 92538 150096
rect 117222 150084 117228 150096
rect 117280 150084 117286 150136
rect 116486 150056 116492 150068
rect 84166 150028 116492 150056
rect 116486 150016 116492 150028
rect 116544 150016 116550 150068
rect 111150 148316 111156 148368
rect 111208 148356 111214 148368
rect 117038 148356 117044 148368
rect 111208 148328 117044 148356
rect 111208 148316 111214 148328
rect 117038 148316 117044 148328
rect 117096 148316 117102 148368
rect 113082 140700 113088 140752
rect 113140 140740 113146 140752
rect 116118 140740 116124 140752
rect 113140 140712 116124 140740
rect 113140 140700 113146 140712
rect 116118 140700 116124 140712
rect 116176 140700 116182 140752
rect 112990 137912 112996 137964
rect 113048 137952 113054 137964
rect 116118 137952 116124 137964
rect 113048 137924 116124 137952
rect 113048 137912 113054 137924
rect 116118 137912 116124 137924
rect 116176 137912 116182 137964
rect 112898 133832 112904 133884
rect 112956 133872 112962 133884
rect 116026 133872 116032 133884
rect 112956 133844 116032 133872
rect 112956 133832 112962 133844
rect 116026 133832 116032 133844
rect 116084 133832 116090 133884
rect 114186 132608 114192 132660
rect 114244 132648 114250 132660
rect 115198 132648 115204 132660
rect 114244 132620 115204 132648
rect 114244 132608 114250 132620
rect 115198 132608 115204 132620
rect 115256 132608 115262 132660
rect 112806 132404 112812 132456
rect 112864 132444 112870 132456
rect 116118 132444 116124 132456
rect 112864 132416 116124 132444
rect 112864 132404 112870 132416
rect 116118 132404 116124 132416
rect 116176 132404 116182 132456
rect 112714 126896 112720 126948
rect 112772 126936 112778 126948
rect 116118 126936 116124 126948
rect 112772 126908 116124 126936
rect 112772 126896 112778 126908
rect 116118 126896 116124 126908
rect 116176 126896 116182 126948
rect 112622 124108 112628 124160
rect 112680 124148 112686 124160
rect 116118 124148 116124 124160
rect 112680 124120 116124 124148
rect 112680 124108 112686 124120
rect 116118 124108 116124 124120
rect 116176 124108 116182 124160
rect 112530 122748 112536 122800
rect 112588 122788 112594 122800
rect 115934 122788 115940 122800
rect 112588 122760 115940 122788
rect 112588 122748 112594 122760
rect 115934 122748 115940 122760
rect 115992 122748 115998 122800
rect 111702 121388 111708 121440
rect 111760 121428 111766 121440
rect 116118 121428 116124 121440
rect 111760 121400 116124 121428
rect 111760 121388 111766 121400
rect 116118 121388 116124 121400
rect 116176 121388 116182 121440
rect 112438 118600 112444 118652
rect 112496 118640 112502 118652
rect 116118 118640 116124 118652
rect 112496 118612 116124 118640
rect 112496 118600 112502 118612
rect 116118 118600 116124 118612
rect 116176 118600 116182 118652
rect 111610 117240 111616 117292
rect 111668 117280 111674 117292
rect 116118 117280 116124 117292
rect 111668 117252 116124 117280
rect 111668 117240 111674 117252
rect 116118 117240 116124 117252
rect 116176 117240 116182 117292
rect 111518 114452 111524 114504
rect 111576 114492 111582 114504
rect 116118 114492 116124 114504
rect 111576 114464 116124 114492
rect 111576 114452 111582 114464
rect 116118 114452 116124 114464
rect 116176 114452 116182 114504
rect 111426 113092 111432 113144
rect 111484 113132 111490 113144
rect 115934 113132 115940 113144
rect 111484 113104 115940 113132
rect 111484 113092 111490 113104
rect 115934 113092 115940 113104
rect 115992 113092 115998 113144
rect 111334 111732 111340 111784
rect 111392 111772 111398 111784
rect 116118 111772 116124 111784
rect 111392 111744 116124 111772
rect 111392 111732 111398 111744
rect 116118 111732 116124 111744
rect 116176 111732 116182 111784
rect 111150 108944 111156 108996
rect 111208 108984 111214 108996
rect 116118 108984 116124 108996
rect 111208 108956 116124 108984
rect 111208 108944 111214 108956
rect 116118 108944 116124 108956
rect 116176 108944 116182 108996
rect 111242 92420 111248 92472
rect 111300 92460 111306 92472
rect 116118 92460 116124 92472
rect 111300 92432 116124 92460
rect 111300 92420 111306 92432
rect 116118 92420 116124 92432
rect 116176 92420 116182 92472
rect 111058 89632 111064 89684
rect 111116 89672 111122 89684
rect 116118 89672 116124 89684
rect 111116 89644 116124 89672
rect 111116 89632 111122 89644
rect 116118 89632 116124 89644
rect 116176 89632 116182 89684
rect 113818 88272 113824 88324
rect 113876 88312 113882 88324
rect 116026 88312 116032 88324
rect 113876 88284 116032 88312
rect 113876 88272 113882 88284
rect 116026 88272 116032 88284
rect 116084 88272 116090 88324
rect 113910 83920 113916 83972
rect 113968 83960 113974 83972
rect 116578 83960 116584 83972
rect 113968 83932 116584 83960
rect 113968 83920 113974 83932
rect 116578 83920 116584 83932
rect 116636 83920 116642 83972
rect 114002 82764 114008 82816
rect 114060 82804 114066 82816
rect 116210 82804 116216 82816
rect 114060 82776 116216 82804
rect 114060 82764 114066 82776
rect 116210 82764 116216 82776
rect 116268 82764 116274 82816
rect 114094 79976 114100 80028
rect 114152 80016 114158 80028
rect 115934 80016 115940 80028
rect 114152 79988 115940 80016
rect 114152 79976 114158 79988
rect 115934 79976 115940 79988
rect 115992 79976 115998 80028
rect 114186 78616 114192 78668
rect 114244 78656 114250 78668
rect 116118 78656 116124 78668
rect 114244 78628 116124 78656
rect 114244 78616 114250 78628
rect 116118 78616 116124 78628
rect 116176 78616 116182 78668
rect 114186 71748 114192 71800
rect 114244 71788 114250 71800
rect 116578 71788 116584 71800
rect 114244 71760 116584 71788
rect 114244 71748 114250 71760
rect 116578 71748 116584 71760
rect 116636 71748 116642 71800
rect 114094 69028 114100 69080
rect 114152 69068 114158 69080
rect 116302 69068 116308 69080
rect 114152 69040 116308 69068
rect 114152 69028 114158 69040
rect 116302 69028 116308 69040
rect 116360 69028 116366 69080
rect 114002 67600 114008 67652
rect 114060 67640 114066 67652
rect 116118 67640 116124 67652
rect 114060 67612 116124 67640
rect 114060 67600 114066 67612
rect 116118 67600 116124 67612
rect 116176 67600 116182 67652
rect 113910 66240 113916 66292
rect 113968 66280 113974 66292
rect 116578 66280 116584 66292
rect 113968 66252 116584 66280
rect 113968 66240 113974 66252
rect 116578 66240 116584 66252
rect 116636 66240 116642 66292
rect 113358 64676 113364 64728
rect 113416 64716 113422 64728
rect 116578 64716 116584 64728
rect 113416 64688 116584 64716
rect 113416 64676 113422 64688
rect 116578 64676 116584 64688
rect 116636 64676 116642 64728
rect 113818 63520 113824 63572
rect 113876 63560 113882 63572
rect 116210 63560 116216 63572
rect 113876 63532 116216 63560
rect 113876 63520 113882 63532
rect 116210 63520 116216 63532
rect 116268 63520 116274 63572
rect 112438 62092 112444 62144
rect 112496 62132 112502 62144
rect 116118 62132 116124 62144
rect 112496 62104 116124 62132
rect 112496 62092 112502 62104
rect 116118 62092 116124 62104
rect 116176 62092 116182 62144
rect 112530 42780 112536 42832
rect 112588 42820 112594 42832
rect 116118 42820 116124 42832
rect 112588 42792 116124 42820
rect 112588 42780 112594 42792
rect 116118 42780 116124 42792
rect 116176 42780 116182 42832
rect 116670 7896 116676 7948
rect 116728 7896 116734 7948
rect 116854 7896 116860 7948
rect 116912 7896 116918 7948
rect 116688 7596 116716 7896
rect 116872 7744 116900 7896
rect 117038 7760 117044 7812
rect 117096 7800 117102 7812
rect 117314 7800 117320 7812
rect 117096 7772 117320 7800
rect 117096 7760 117102 7772
rect 117314 7760 117320 7772
rect 117372 7760 117378 7812
rect 116854 7692 116860 7744
rect 116912 7692 116918 7744
rect 116762 7624 116768 7676
rect 116820 7664 116826 7676
rect 117222 7664 117228 7676
rect 116820 7636 117228 7664
rect 116820 7624 116826 7636
rect 117222 7624 117228 7636
rect 117280 7624 117286 7676
rect 116688 7568 116992 7596
rect 116964 7460 116992 7568
rect 117038 7460 117044 7472
rect 116964 7432 117044 7460
rect 117038 7420 117044 7432
rect 117096 7420 117102 7472
rect 170140 3012 179414 3040
rect 111702 2864 111708 2916
rect 111760 2904 111766 2916
rect 111760 2876 170076 2904
rect 111760 2864 111766 2876
rect 111794 2796 111800 2848
rect 111852 2836 111858 2848
rect 111852 2808 168374 2836
rect 111852 2796 111858 2808
rect 168346 2360 168374 2808
rect 170048 2774 170076 2876
rect 169956 2746 170076 2774
rect 169956 2700 169984 2746
rect 169680 2672 169984 2700
rect 170140 2700 170168 3012
rect 179386 2972 179414 3012
rect 180766 3012 183554 3040
rect 180766 2972 180794 3012
rect 179386 2944 180794 2972
rect 183526 2972 183554 3012
rect 183526 2944 200114 2972
rect 183526 2876 186452 2904
rect 183526 2768 183554 2876
rect 186424 2836 186452 2876
rect 200086 2836 200114 2944
rect 186424 2808 193444 2836
rect 200086 2808 293954 2836
rect 182146 2740 183554 2768
rect 182146 2700 182174 2740
rect 170140 2672 170352 2700
rect 169680 2428 169708 2672
rect 170324 2508 170352 2672
rect 178006 2672 182174 2700
rect 178006 2632 178034 2672
rect 176626 2604 178034 2632
rect 170306 2456 170312 2508
rect 170364 2456 170370 2508
rect 176626 2428 176654 2604
rect 193416 2496 193444 2808
rect 193582 2496 193588 2508
rect 193416 2468 193588 2496
rect 193582 2456 193588 2468
rect 193640 2456 193646 2508
rect 293926 2496 293954 2808
rect 425808 2808 443684 2836
rect 425808 2508 425836 2808
rect 443656 2508 443684 2808
rect 294782 2496 294788 2508
rect 293926 2468 294788 2496
rect 294782 2456 294788 2468
rect 294840 2456 294846 2508
rect 425790 2456 425796 2508
rect 425848 2456 425854 2508
rect 443638 2456 443644 2508
rect 443696 2456 443702 2508
rect 169680 2400 176654 2428
rect 170306 2360 170312 2372
rect 168346 2332 170312 2360
rect 170306 2320 170312 2332
rect 170364 2320 170370 2372
rect 111058 1952 111064 1964
rect 99346 1924 104480 1952
rect 62390 1844 62396 1896
rect 62448 1884 62454 1896
rect 65334 1884 65340 1896
rect 62448 1856 65340 1884
rect 62448 1844 62454 1856
rect 65334 1844 65340 1856
rect 65392 1844 65398 1896
rect 68002 1844 68008 1896
rect 68060 1884 68066 1896
rect 77110 1884 77116 1896
rect 68060 1856 77116 1884
rect 68060 1844 68066 1856
rect 77110 1844 77116 1856
rect 77168 1844 77174 1896
rect 77754 1844 77760 1896
rect 77812 1884 77818 1896
rect 89254 1884 89260 1896
rect 77812 1856 89260 1884
rect 77812 1844 77818 1856
rect 89254 1844 89260 1856
rect 89312 1844 89318 1896
rect 89346 1844 89352 1896
rect 89404 1884 89410 1896
rect 99346 1884 99374 1924
rect 89404 1856 99374 1884
rect 89404 1844 89410 1856
rect 99650 1844 99656 1896
rect 99708 1884 99714 1896
rect 104342 1884 104348 1896
rect 99708 1856 104348 1884
rect 99708 1844 99714 1856
rect 104342 1844 104348 1856
rect 104400 1844 104406 1896
rect 64138 1776 64144 1828
rect 64196 1816 64202 1828
rect 69382 1816 69388 1828
rect 64196 1788 69388 1816
rect 64196 1776 64202 1788
rect 69382 1776 69388 1788
rect 69440 1776 69446 1828
rect 77018 1776 77024 1828
rect 77076 1816 77082 1828
rect 85942 1816 85948 1828
rect 77076 1788 85948 1816
rect 77076 1776 77082 1788
rect 85942 1776 85948 1788
rect 86000 1776 86006 1828
rect 86034 1776 86040 1828
rect 86092 1816 86098 1828
rect 104452 1816 104480 1924
rect 105832 1924 111064 1952
rect 105832 1896 105860 1924
rect 111058 1912 111064 1924
rect 111116 1912 111122 1964
rect 104526 1844 104532 1896
rect 104584 1884 104590 1896
rect 105722 1884 105728 1896
rect 104584 1856 105728 1884
rect 104584 1844 104590 1856
rect 105722 1844 105728 1856
rect 105780 1844 105786 1896
rect 105814 1844 105820 1896
rect 105872 1844 105878 1896
rect 105906 1844 105912 1896
rect 105964 1884 105970 1896
rect 109218 1884 109224 1896
rect 105964 1856 109224 1884
rect 105964 1844 105970 1856
rect 109218 1844 109224 1856
rect 109276 1844 109282 1896
rect 109310 1844 109316 1896
rect 109368 1884 109374 1896
rect 109368 1856 110184 1884
rect 109368 1844 109374 1856
rect 109586 1816 109592 1828
rect 86092 1788 104204 1816
rect 104452 1788 109592 1816
rect 86092 1776 86098 1788
rect 62666 1708 62672 1760
rect 62724 1748 62730 1760
rect 68830 1748 68836 1760
rect 62724 1720 68836 1748
rect 62724 1708 62730 1720
rect 68830 1708 68836 1720
rect 68888 1708 68894 1760
rect 79962 1708 79968 1760
rect 80020 1748 80026 1760
rect 80790 1748 80796 1760
rect 80020 1720 80796 1748
rect 80020 1708 80026 1720
rect 80790 1708 80796 1720
rect 80848 1708 80854 1760
rect 82630 1708 82636 1760
rect 82688 1748 82694 1760
rect 104066 1748 104072 1760
rect 82688 1720 104072 1748
rect 82688 1708 82694 1720
rect 104066 1708 104072 1720
rect 104124 1708 104130 1760
rect 104176 1748 104204 1788
rect 109586 1776 109592 1788
rect 109644 1776 109650 1828
rect 109954 1748 109960 1760
rect 104176 1720 109960 1748
rect 109954 1708 109960 1720
rect 110012 1708 110018 1760
rect 110156 1748 110184 1856
rect 112438 1748 112444 1760
rect 110156 1720 112444 1748
rect 112438 1708 112444 1720
rect 112496 1708 112502 1760
rect 69290 1640 69296 1692
rect 69348 1680 69354 1692
rect 102594 1680 102600 1692
rect 69348 1652 102600 1680
rect 69348 1640 69354 1652
rect 102594 1640 102600 1652
rect 102652 1640 102658 1692
rect 102686 1640 102692 1692
rect 102744 1680 102750 1692
rect 105814 1680 105820 1692
rect 102744 1652 105820 1680
rect 102744 1640 102750 1652
rect 105814 1640 105820 1652
rect 105872 1640 105878 1692
rect 106182 1640 106188 1692
rect 106240 1680 106246 1692
rect 116578 1680 116584 1692
rect 106240 1652 116584 1680
rect 106240 1640 106246 1652
rect 116578 1640 116584 1652
rect 116636 1640 116642 1692
rect 59354 1572 59360 1624
rect 59412 1612 59418 1624
rect 68462 1612 68468 1624
rect 59412 1584 68468 1612
rect 59412 1572 59418 1584
rect 68462 1572 68468 1584
rect 68520 1572 68526 1624
rect 79318 1572 79324 1624
rect 79376 1612 79382 1624
rect 99466 1612 99472 1624
rect 79376 1584 99472 1612
rect 79376 1572 79382 1584
rect 99466 1572 99472 1584
rect 99524 1572 99530 1624
rect 99558 1572 99564 1624
rect 99616 1612 99622 1624
rect 105906 1612 105912 1624
rect 99616 1584 105912 1612
rect 99616 1572 99622 1584
rect 105906 1572 105912 1584
rect 105964 1572 105970 1624
rect 105998 1572 106004 1624
rect 106056 1612 106062 1624
rect 110138 1612 110144 1624
rect 106056 1584 110144 1612
rect 106056 1572 106062 1584
rect 110138 1572 110144 1584
rect 110196 1572 110202 1624
rect 72694 1504 72700 1556
rect 72752 1544 72758 1556
rect 110506 1544 110512 1556
rect 72752 1516 99374 1544
rect 72752 1504 72758 1516
rect 42610 1436 42616 1488
rect 42668 1476 42674 1488
rect 80422 1476 80428 1488
rect 42668 1448 80428 1476
rect 42668 1436 42674 1448
rect 80422 1436 80428 1448
rect 80480 1436 80486 1488
rect 94130 1436 94136 1488
rect 94188 1476 94194 1488
rect 96614 1476 96620 1488
rect 94188 1448 96620 1476
rect 94188 1436 94194 1448
rect 96614 1436 96620 1448
rect 96672 1436 96678 1488
rect 99346 1476 99374 1516
rect 99576 1516 110512 1544
rect 99576 1476 99604 1516
rect 110506 1504 110512 1516
rect 110564 1504 110570 1556
rect 99346 1448 99604 1476
rect 99650 1436 99656 1488
rect 99708 1476 99714 1488
rect 108206 1476 108212 1488
rect 99708 1448 108212 1476
rect 99708 1436 99714 1448
rect 108206 1436 108212 1448
rect 108264 1436 108270 1488
rect 108298 1436 108304 1488
rect 108356 1476 108362 1488
rect 143626 1476 143632 1488
rect 108356 1448 143632 1476
rect 108356 1436 108362 1448
rect 143626 1436 143632 1448
rect 143684 1436 143690 1488
rect 46014 1368 46020 1420
rect 46072 1408 46078 1420
rect 116486 1408 116492 1420
rect 46072 1380 116492 1408
rect 46072 1368 46078 1380
rect 116486 1368 116492 1380
rect 116544 1368 116550 1420
rect 294782 1368 294788 1420
rect 294840 1408 294846 1420
rect 343634 1408 343640 1420
rect 294840 1380 343640 1408
rect 294840 1368 294846 1380
rect 343634 1368 343640 1380
rect 343692 1368 343698 1420
rect 491294 1368 491300 1420
rect 491352 1408 491358 1420
rect 493594 1408 493600 1420
rect 491352 1380 493600 1408
rect 491352 1368 491358 1380
rect 493594 1368 493600 1380
rect 493652 1368 493658 1420
rect 2682 1300 2688 1352
rect 2740 1340 2746 1352
rect 116302 1340 116308 1352
rect 2740 1312 116308 1340
rect 2740 1300 2746 1312
rect 116302 1300 116308 1312
rect 116360 1300 116366 1352
rect 39298 1232 39304 1284
rect 39356 1272 39362 1284
rect 116394 1272 116400 1284
rect 39356 1244 116400 1272
rect 39356 1232 39362 1244
rect 116394 1232 116400 1244
rect 116452 1232 116458 1284
rect 49326 1164 49332 1216
rect 49384 1204 49390 1216
rect 116762 1204 116768 1216
rect 49384 1176 116768 1204
rect 49384 1164 49390 1176
rect 116762 1164 116768 1176
rect 116820 1164 116826 1216
rect 52638 1096 52644 1148
rect 52696 1136 52702 1148
rect 117222 1136 117228 1148
rect 52696 1108 117228 1136
rect 52696 1096 52702 1108
rect 117222 1096 117228 1108
rect 117280 1096 117286 1148
rect 55950 1028 55956 1080
rect 56008 1068 56014 1080
rect 111794 1068 111800 1080
rect 56008 1040 111800 1068
rect 56008 1028 56014 1040
rect 111794 1028 111800 1040
rect 111852 1028 111858 1080
rect 65978 960 65984 1012
rect 66036 1000 66042 1012
rect 116854 1000 116860 1012
rect 66036 972 116860 1000
rect 66036 960 66042 972
rect 116854 960 116860 972
rect 116912 960 116918 1012
rect 76006 892 76012 944
rect 76064 932 76070 944
rect 112530 932 112536 944
rect 76064 904 112536 932
rect 76064 892 76070 904
rect 112530 892 112536 904
rect 112588 892 112594 944
rect 94682 824 94688 876
rect 94740 864 94746 876
rect 100110 864 100116 876
rect 94740 836 100116 864
rect 94740 824 94746 836
rect 100110 824 100116 836
rect 100168 824 100174 876
rect 96338 756 96344 808
rect 96396 796 96402 808
rect 101858 796 101864 808
rect 96396 768 101864 796
rect 96396 756 96402 768
rect 101858 756 101864 768
rect 101916 756 101922 808
<< via1 >>
rect 213184 160216 213236 160268
rect 221188 160216 221240 160268
rect 126520 160080 126572 160132
rect 134156 160080 134208 160132
rect 63408 160012 63460 160064
rect 146484 160012 146536 160064
rect 146944 160012 146996 160064
rect 154488 160012 154540 160064
rect 156788 160012 156840 160064
rect 191748 160012 191800 160064
rect 197176 160012 197228 160064
rect 207020 160012 207072 160064
rect 211436 160012 211488 160064
rect 280344 160012 280396 160064
rect 281264 160012 281316 160064
rect 332692 160012 332744 160064
rect 334256 160012 334308 160064
rect 374092 160012 374144 160064
rect 378876 160012 378928 160064
rect 398104 160012 398156 160064
rect 409972 160012 410024 160064
rect 417884 160012 417936 160064
rect 25596 159944 25648 159996
rect 109776 159944 109828 159996
rect 117228 159944 117280 159996
rect 191472 159944 191524 159996
rect 198004 159944 198056 159996
rect 269120 159944 269172 159996
rect 271236 159944 271288 159996
rect 272800 159944 272852 159996
rect 275376 159944 275428 159996
rect 328460 159944 328512 159996
rect 329196 159944 329248 159996
rect 369952 159944 370004 159996
rect 374644 159944 374696 159996
rect 388352 159944 388404 159996
rect 389824 159944 389876 159996
rect 413836 159944 413888 159996
rect 449532 159944 449584 159996
rect 456156 159944 456208 159996
rect 457076 159944 457128 159996
rect 463884 159944 463936 159996
rect 469680 159944 469732 159996
rect 477408 159944 477460 159996
rect 76932 159876 76984 159928
rect 162492 159876 162544 159928
rect 166908 159876 166960 159928
rect 186412 159876 186464 159928
rect 191288 159876 191340 159928
rect 264888 159876 264940 159928
rect 268660 159876 268712 159928
rect 324044 159876 324096 159928
rect 328368 159876 328420 159928
rect 369492 159876 369544 159928
rect 372160 159876 372212 159928
rect 396172 159876 396224 159928
rect 403256 159876 403308 159928
rect 416596 159876 416648 159928
rect 480628 159876 480680 159928
rect 485964 159876 486016 159928
rect 70124 159808 70176 159860
rect 153384 159808 153436 159860
rect 153476 159808 153528 159860
rect 179420 159808 179472 159860
rect 184572 159808 184624 159860
rect 259552 159808 259604 159860
rect 261944 159808 261996 159860
rect 312360 159808 312412 159860
rect 312452 159808 312504 159860
rect 313372 159808 313424 159860
rect 322480 159808 322532 159860
rect 365168 159808 365220 159860
rect 376300 159808 376352 159860
rect 406200 159808 406252 159860
rect 424324 159808 424376 159860
rect 442724 159808 442776 159860
rect 450360 159808 450412 159860
rect 456892 159808 456944 159860
rect 458732 159808 458784 159860
rect 465080 159808 465132 159860
rect 468024 159808 468076 159860
rect 476028 159808 476080 159860
rect 479800 159808 479852 159860
rect 485228 159808 485280 159860
rect 56692 159740 56744 159792
rect 131212 159740 131264 159792
rect 18880 159672 18932 159724
rect 109132 159672 109184 159724
rect 113088 159672 113140 159724
rect 126428 159672 126480 159724
rect 49976 159604 50028 159656
rect 143264 159740 143316 159792
rect 143356 159740 143408 159792
rect 160100 159740 160152 159792
rect 171140 159740 171192 159792
rect 173256 159740 173308 159792
rect 177856 159740 177908 159792
rect 253940 159740 253992 159792
rect 255228 159740 255280 159792
rect 313464 159740 313516 159792
rect 314108 159740 314160 159792
rect 357992 159740 358044 159792
rect 365444 159740 365496 159792
rect 395528 159740 395580 159792
rect 396540 159740 396592 159792
rect 413744 159740 413796 159792
rect 420920 159740 420972 159792
rect 440424 159740 440476 159792
rect 134156 159672 134208 159724
rect 156512 159672 156564 159724
rect 131672 159604 131724 159656
rect 136548 159604 136600 159656
rect 136640 159604 136692 159656
rect 139400 159604 139452 159656
rect 139952 159604 140004 159656
rect 163780 159672 163832 159724
rect 167736 159672 167788 159724
rect 246948 159672 247000 159724
rect 248512 159672 248564 159724
rect 161020 159604 161072 159656
rect 240232 159604 240284 159656
rect 244280 159604 244332 159656
rect 305368 159604 305420 159656
rect 308220 159672 308272 159724
rect 342628 159672 342680 159724
rect 342720 159672 342772 159724
rect 343824 159672 343876 159724
rect 347780 159672 347832 159724
rect 378784 159672 378836 159724
rect 379704 159672 379756 159724
rect 405832 159672 405884 159724
rect 417516 159672 417568 159724
rect 437664 159672 437716 159724
rect 308588 159604 308640 159656
rect 309048 159604 309100 159656
rect 341616 159604 341668 159656
rect 43260 159536 43312 159588
rect 32312 159468 32364 159520
rect 36544 159400 36596 159452
rect 126244 159400 126296 159452
rect 126428 159468 126480 159520
rect 127808 159468 127860 159520
rect 129924 159536 129976 159588
rect 146944 159536 146996 159588
rect 153384 159536 153436 159588
rect 156788 159536 156840 159588
rect 157616 159536 157668 159588
rect 239312 159536 239364 159588
rect 250996 159536 251048 159588
rect 310612 159536 310664 159588
rect 315764 159536 315816 159588
rect 342812 159604 342864 159656
rect 354220 159604 354272 159656
rect 357440 159604 357492 159656
rect 363144 159604 363196 159656
rect 369584 159604 369636 159656
rect 401048 159604 401100 159656
rect 407488 159604 407540 159656
rect 429936 159604 429988 159656
rect 478972 159604 479024 159656
rect 484584 159604 484636 159656
rect 358912 159536 358964 159588
rect 362868 159536 362920 159588
rect 394976 159536 395028 159588
rect 399024 159536 399076 159588
rect 408500 159536 408552 159588
rect 410800 159536 410852 159588
rect 432512 159536 432564 159588
rect 467196 159536 467248 159588
rect 473360 159536 473412 159588
rect 131120 159468 131172 159520
rect 131212 159468 131264 159520
rect 144092 159468 144144 159520
rect 144184 159468 144236 159520
rect 225328 159468 225380 159520
rect 230848 159468 230900 159520
rect 293960 159468 294012 159520
rect 294788 159468 294840 159520
rect 126796 159400 126848 159452
rect 6276 159332 6328 159384
rect 122840 159332 122892 159384
rect 123116 159332 123168 159384
rect 147496 159400 147548 159452
rect 147588 159400 147640 159452
rect 149520 159400 149572 159452
rect 150900 159400 150952 159452
rect 233240 159400 233292 159452
rect 234988 159400 235040 159452
rect 298008 159400 298060 159452
rect 301504 159400 301556 159452
rect 341432 159400 341484 159452
rect 341616 159468 341668 159520
rect 354864 159468 354916 159520
rect 356152 159468 356204 159520
rect 390560 159468 390612 159520
rect 400772 159468 400824 159520
rect 424876 159468 424928 159520
rect 448704 159468 448756 159520
rect 456064 159468 456116 159520
rect 457904 159468 457956 159520
rect 464712 159468 464764 159520
rect 342260 159400 342312 159452
rect 342352 159400 342404 159452
rect 349344 159400 349396 159452
rect 358636 159400 358688 159452
rect 392768 159400 392820 159452
rect 404084 159400 404136 159452
rect 427360 159400 427412 159452
rect 427636 159400 427688 159452
rect 445392 159400 445444 159452
rect 451188 159400 451240 159452
rect 456800 159400 456852 159452
rect 459652 159400 459704 159452
rect 466460 159400 466512 159452
rect 468852 159400 468904 159452
rect 474832 159400 474884 159452
rect 477316 159400 477368 159452
rect 483296 159400 483348 159452
rect 518808 159400 518860 159452
rect 522672 159400 522724 159452
rect 129924 159332 129976 159384
rect 137100 159332 137152 159384
rect 137468 159332 137520 159384
rect 223580 159332 223632 159384
rect 231676 159332 231728 159384
rect 295524 159332 295576 159384
rect 295616 159332 295668 159384
rect 342444 159332 342496 159384
rect 346032 159332 346084 159384
rect 382832 159332 382884 159384
rect 383108 159332 383160 159384
rect 411352 159332 411404 159384
rect 414204 159332 414256 159384
rect 435088 159332 435140 159384
rect 447876 159332 447928 159384
rect 456984 159332 457036 159384
rect 470508 159332 470560 159384
rect 476120 159332 476172 159384
rect 478144 159332 478196 159384
rect 483204 159332 483256 159384
rect 518716 159332 518768 159384
rect 523500 159332 523552 159384
rect 73528 159264 73580 159316
rect 80060 159264 80112 159316
rect 83648 159264 83700 159316
rect 167000 159264 167052 159316
rect 170220 159264 170272 159316
rect 198924 159264 198976 159316
rect 201408 159264 201460 159316
rect 212632 159264 212684 159316
rect 214012 159264 214064 159316
rect 281540 159264 281592 159316
rect 282092 159264 282144 159316
rect 334348 159264 334400 159316
rect 335084 159264 335136 159316
rect 374736 159264 374788 159316
rect 388996 159264 389048 159316
rect 403900 159264 403952 159316
rect 460480 159264 460532 159316
rect 466644 159264 466696 159316
rect 80244 159196 80296 159248
rect 91100 159196 91152 159248
rect 100484 159196 100536 159248
rect 184388 159196 184440 159248
rect 187056 159196 187108 159248
rect 214656 159196 214708 159248
rect 218244 159196 218296 159248
rect 284392 159196 284444 159248
rect 287980 159196 288032 159248
rect 338764 159196 338816 159248
rect 339316 159196 339368 159248
rect 377956 159196 378008 159248
rect 86960 159128 87012 159180
rect 93676 159060 93728 159112
rect 162860 159060 162912 159112
rect 163044 159128 163096 159180
rect 172152 159128 172204 159180
rect 193772 159128 193824 159180
rect 218060 159128 218112 159180
rect 224960 159128 225012 159180
rect 290648 159128 290700 159180
rect 293960 159128 294012 159180
rect 295156 159128 295208 159180
rect 302332 159128 302384 159180
rect 169760 159060 169812 159112
rect 173624 159060 173676 159112
rect 197360 159060 197412 159112
rect 203892 159060 203944 159112
rect 212724 159060 212776 159112
rect 220728 159060 220780 159112
rect 283196 159060 283248 159112
rect 284668 159060 284720 159112
rect 285772 159060 285824 159112
rect 107200 158992 107252 159044
rect 183468 158992 183520 159044
rect 183744 158992 183796 159044
rect 201408 158992 201460 159044
rect 214840 158992 214892 159044
rect 222108 158992 222160 159044
rect 224132 158992 224184 159044
rect 288072 159060 288124 159112
rect 288900 159060 288952 159112
rect 338396 159060 338448 159112
rect 338488 159060 338540 159112
rect 339684 159060 339736 159112
rect 341432 159128 341484 159180
rect 345664 159128 345716 159180
rect 345756 159128 345808 159180
rect 351828 159128 351880 159180
rect 351920 159128 351972 159180
rect 385500 159196 385552 159248
rect 385592 159196 385644 159248
rect 398840 159196 398892 159248
rect 349252 159060 349304 159112
rect 349344 159060 349396 159112
rect 376944 159060 376996 159112
rect 378048 159060 378100 159112
rect 388444 159128 388496 159180
rect 392308 159128 392360 159180
rect 404268 159128 404320 159180
rect 461308 159128 461360 159180
rect 467840 159128 467892 159180
rect 472256 159128 472308 159180
rect 479432 159128 479484 159180
rect 395712 159060 395764 159112
rect 404636 159060 404688 159112
rect 452016 159060 452068 159112
rect 458180 159060 458232 159112
rect 462136 159060 462188 159112
rect 467932 159060 467984 159112
rect 471428 159060 471480 159112
rect 477684 159060 477736 159112
rect 298100 158992 298152 159044
rect 300400 158992 300452 159044
rect 307392 158992 307444 159044
rect 345572 158992 345624 159044
rect 345848 158992 345900 159044
rect 349068 158992 349120 159044
rect 351092 158992 351144 159044
rect 382556 158992 382608 159044
rect 455420 158992 455472 159044
rect 463516 158992 463568 159044
rect 465540 158992 465592 159044
rect 472532 158992 472584 159044
rect 473912 158992 473964 159044
rect 480720 158992 480772 159044
rect 96252 158924 96304 158976
rect 121920 158924 121972 158976
rect 124036 158924 124088 158976
rect 194140 158924 194192 158976
rect 200580 158924 200632 158976
rect 224960 158924 225012 158976
rect 237564 158924 237616 158976
rect 299480 158924 299532 158976
rect 314936 158924 314988 158976
rect 357532 158924 357584 158976
rect 357808 158924 357860 158976
rect 384948 158924 385000 158976
rect 420092 158924 420144 158976
rect 423496 158924 423548 158976
rect 446128 158924 446180 158976
rect 453948 158924 454000 158976
rect 456248 158924 456300 158976
rect 463608 158924 463660 158976
rect 464620 158924 464672 158976
rect 471428 158924 471480 158976
rect 475568 158924 475620 158976
rect 481640 158924 481692 158976
rect 102968 158856 103020 158908
rect 125508 158856 125560 158908
rect 126244 158856 126296 158908
rect 129740 158856 129792 158908
rect 130752 158856 130804 158908
rect 194600 158856 194652 158908
rect 194692 158856 194744 158908
rect 203708 158856 203760 158908
rect 208124 158856 208176 158908
rect 212448 158856 212500 158908
rect 109684 158788 109736 158840
rect 129924 158788 129976 158840
rect 133236 158788 133288 158840
rect 158720 158788 158772 158840
rect 163504 158788 163556 158840
rect 195980 158788 196032 158840
rect 207296 158788 207348 158840
rect 230756 158856 230808 158908
rect 241796 158856 241848 158908
rect 303528 158856 303580 158908
rect 305644 158856 305696 158908
rect 307392 158856 307444 158908
rect 310704 158856 310756 158908
rect 312176 158856 312228 158908
rect 312360 158856 312412 158908
rect 318892 158856 318944 158908
rect 320824 158856 320876 158908
rect 217324 158788 217376 158840
rect 220360 158788 220412 158840
rect 238392 158788 238444 158840
rect 241612 158788 241664 158840
rect 261116 158788 261168 158840
rect 317052 158788 317104 158840
rect 319168 158788 319220 158840
rect 90364 158720 90416 158772
rect 92572 158720 92624 158772
rect 92848 158720 92900 158772
rect 114468 158720 114520 158772
rect 119804 158720 119856 158772
rect 146576 158720 146628 158772
rect 146668 158720 146720 158772
rect 176660 158720 176712 158772
rect 180340 158720 180392 158772
rect 204904 158720 204956 158772
rect 210608 158720 210660 158772
rect 215392 158720 215444 158772
rect 221556 158720 221608 158772
rect 224408 158720 224460 158772
rect 240876 158720 240928 158772
rect 243360 158720 243412 158772
rect 254400 158720 254452 158772
rect 255412 158720 255464 158772
rect 258540 158720 258592 158772
rect 260932 158720 260984 158772
rect 264428 158720 264480 158772
rect 266360 158720 266412 158772
rect 267832 158720 267884 158772
rect 320272 158720 320324 158772
rect 321652 158788 321704 158840
rect 357440 158788 357492 158840
rect 361212 158856 361264 158908
rect 376760 158856 376812 158908
rect 376944 158856 376996 158908
rect 378232 158856 378284 158908
rect 362960 158788 363012 158840
rect 367928 158788 367980 158840
rect 386144 158856 386196 158908
rect 391480 158856 391532 158908
rect 393688 158856 393740 158908
rect 412548 158856 412600 158908
rect 412916 158856 412968 158908
rect 454592 158856 454644 158908
rect 462228 158856 462280 158908
rect 466368 158856 466420 158908
rect 472440 158856 472492 158908
rect 476396 158856 476448 158908
rect 482652 158856 482704 158908
rect 508320 158856 508372 158908
rect 510068 158856 510120 158908
rect 327540 158720 327592 158772
rect 367192 158720 367244 158772
rect 81072 158652 81124 158704
rect 180892 158652 180944 158704
rect 181996 158652 182048 158704
rect 256792 158652 256844 158704
rect 321560 158652 321612 158704
rect 386236 158788 386288 158840
rect 388076 158788 388128 158840
rect 390376 158788 390428 158840
rect 409144 158788 409196 158840
rect 410800 158788 410852 158840
rect 416688 158788 416740 158840
rect 419540 158788 419592 158840
rect 452844 158788 452896 158840
rect 459652 158788 459704 158840
rect 463792 158788 463844 158840
rect 471336 158788 471388 158840
rect 474740 158788 474792 158840
rect 480260 158788 480312 158840
rect 482284 158788 482336 158840
rect 487252 158788 487304 158840
rect 506388 158788 506440 158840
rect 507584 158788 507636 158840
rect 67640 158584 67692 158636
rect 170312 158584 170364 158636
rect 171968 158584 172020 158636
rect 250076 158584 250128 158636
rect 376760 158584 376812 158636
rect 384764 158720 384816 158772
rect 389180 158720 389232 158772
rect 405740 158720 405792 158772
rect 409236 158720 409288 158772
rect 413376 158720 413428 158772
rect 419632 158720 419684 158772
rect 453764 158720 453816 158772
rect 459560 158720 459612 158772
rect 462964 158720 463016 158772
rect 469220 158720 469272 158772
rect 473084 158720 473136 158772
rect 478972 158720 479024 158772
rect 481456 158720 481508 158772
rect 486516 158720 486568 158772
rect 505284 158720 505336 158772
rect 506756 158720 506808 158772
rect 507032 158720 507084 158772
rect 508412 158720 508464 158772
rect 509424 158720 509476 158772
rect 511724 158720 511776 158772
rect 514944 158720 514996 158772
rect 518532 158720 518584 158772
rect 74356 158516 74408 158568
rect 175188 158516 175240 158568
rect 175280 158516 175332 158568
rect 252744 158516 252796 158568
rect 71044 158448 71096 158500
rect 64236 158380 64288 158432
rect 167552 158380 167604 158432
rect 168564 158380 168616 158432
rect 169668 158380 169720 158432
rect 171784 158448 171836 158500
rect 178040 158448 178092 158500
rect 178684 158448 178736 158500
rect 255596 158448 255648 158500
rect 173072 158380 173124 158432
rect 173164 158380 173216 158432
rect 247132 158380 247184 158432
rect 60924 158312 60976 158364
rect 164332 158312 164384 158364
rect 165252 158312 165304 158364
rect 245016 158312 245068 158364
rect 54208 158244 54260 158296
rect 160284 158244 160336 158296
rect 161848 158244 161900 158296
rect 242072 158244 242124 158296
rect 50804 158176 50856 158228
rect 157708 158176 157760 158228
rect 158444 158176 158496 158228
rect 238944 158176 238996 158228
rect 256884 158176 256936 158228
rect 315028 158176 315080 158228
rect 47492 158108 47544 158160
rect 155040 158108 155092 158160
rect 155132 158108 155184 158160
rect 237380 158108 237432 158160
rect 246764 158108 246816 158160
rect 306932 158108 306984 158160
rect 37372 158040 37424 158092
rect 146392 158040 146444 158092
rect 148416 158040 148468 158092
rect 231952 158040 232004 158092
rect 243452 158040 243504 158092
rect 304724 158040 304776 158092
rect 388 157972 440 158024
rect 118884 157972 118936 158024
rect 131764 157972 131816 158024
rect 219348 157972 219400 158024
rect 236736 157972 236788 158024
rect 299664 157972 299716 158024
rect 77760 157904 77812 157956
rect 171784 157904 171836 157956
rect 171876 157904 171928 157956
rect 182272 157904 182324 157956
rect 87788 157836 87840 157888
rect 84476 157768 84528 157820
rect 171784 157768 171836 157820
rect 185124 157836 185176 157888
rect 179420 157768 179472 157820
rect 185308 157904 185360 157956
rect 185400 157904 185452 157956
rect 260472 157904 260524 157956
rect 188804 157836 188856 157888
rect 263048 157836 263100 157888
rect 91192 157700 91244 157752
rect 185308 157700 185360 157752
rect 94596 157632 94648 157684
rect 190644 157768 190696 157820
rect 195520 157768 195572 157820
rect 267740 157768 267792 157820
rect 185676 157700 185728 157752
rect 188528 157700 188580 157752
rect 190460 157700 190512 157752
rect 263692 157700 263744 157752
rect 185584 157632 185636 157684
rect 236092 157632 236144 157684
rect 97908 157564 97960 157616
rect 193220 157564 193272 157616
rect 197360 157564 197412 157616
rect 251456 157564 251508 157616
rect 111340 157496 111392 157548
rect 203432 157496 203484 157548
rect 204904 157496 204956 157548
rect 255872 157496 255924 157548
rect 114744 157428 114796 157480
rect 206560 157428 206612 157480
rect 214564 157428 214616 157480
rect 141700 157360 141752 157412
rect 49148 157292 49200 157344
rect 156420 157292 156472 157344
rect 158720 157292 158772 157344
rect 210516 157292 210568 157344
rect 227076 157360 227128 157412
rect 214380 157292 214432 157344
rect 221188 157292 221240 157344
rect 45744 157224 45796 157276
rect 153752 157224 153804 157276
rect 163780 157224 163832 157276
rect 166448 157224 166500 157276
rect 192116 157224 192168 157276
rect 265164 157224 265216 157276
rect 42432 157156 42484 157208
rect 151268 157156 151320 157208
rect 156512 157156 156564 157208
rect 159088 157156 159140 157208
rect 160100 157156 160152 157208
rect 166172 157156 166224 157208
rect 166264 157156 166316 157208
rect 171140 157156 171192 157208
rect 177028 157156 177080 157208
rect 254032 157156 254084 157208
rect 283840 157224 283892 157276
rect 335544 157224 335596 157276
rect 281632 157156 281684 157208
rect 300676 157156 300728 157208
rect 348056 157156 348108 157208
rect 39028 157088 39080 157140
rect 147680 157088 147732 157140
rect 150072 157088 150124 157140
rect 233516 157088 233568 157140
rect 287152 157088 287204 157140
rect 338120 157088 338172 157140
rect 35716 157020 35768 157072
rect 146208 157020 146260 157072
rect 151728 157020 151780 157072
rect 234804 157020 234856 157072
rect 280436 157020 280488 157072
rect 333060 157020 333112 157072
rect 24768 156952 24820 157004
rect 137376 156952 137428 157004
rect 138296 156952 138348 157004
rect 224132 156952 224184 157004
rect 273720 156952 273772 157004
rect 327908 156952 327960 157004
rect 21364 156884 21416 156936
rect 135260 156884 135312 156936
rect 135812 156884 135864 156936
rect 222568 156884 222620 156936
rect 224960 156884 225012 156936
rect 272064 156884 272116 156936
rect 277124 156884 277176 156936
rect 330484 156884 330536 156936
rect 18052 156816 18104 156868
rect 132500 156816 132552 156868
rect 134892 156816 134944 156868
rect 210424 156816 210476 156868
rect 210608 156816 210660 156868
rect 214196 156816 214248 156868
rect 219716 156816 219768 156868
rect 14648 156748 14700 156800
rect 130108 156748 130160 156800
rect 139124 156748 139176 156800
rect 225144 156748 225196 156800
rect 226616 156816 226668 156868
rect 291936 156816 291988 156868
rect 293868 156816 293920 156868
rect 342536 156816 342588 156868
rect 228364 156748 228416 156800
rect 230020 156748 230072 156800
rect 294052 156748 294104 156800
rect 297272 156748 297324 156800
rect 345112 156748 345164 156800
rect 11244 156680 11296 156732
rect 127532 156680 127584 156732
rect 128176 156680 128228 156732
rect 216772 156680 216824 156732
rect 223212 156680 223264 156732
rect 289360 156680 289412 156732
rect 290556 156680 290608 156732
rect 340052 156680 340104 156732
rect 2044 156612 2096 156664
rect 120448 156612 120500 156664
rect 124864 156612 124916 156664
rect 209780 156612 209832 156664
rect 209964 156612 210016 156664
rect 211620 156612 211672 156664
rect 216496 156612 216548 156664
rect 283104 156612 283156 156664
rect 498292 156612 498344 156664
rect 499304 156612 499356 156664
rect 502340 156612 502392 156664
rect 503352 156612 503404 156664
rect 52460 156544 52512 156596
rect 158996 156544 159048 156596
rect 159088 156544 159140 156596
rect 200764 156544 200816 156596
rect 200948 156544 201000 156596
rect 270500 156544 270552 156596
rect 59268 156476 59320 156528
rect 164148 156476 164200 156528
rect 166172 156476 166224 156528
rect 69296 156408 69348 156460
rect 166264 156408 166316 156460
rect 166448 156476 166500 156528
rect 225052 156476 225104 156528
rect 219716 156408 219768 156460
rect 219808 156408 219860 156460
rect 221372 156408 221424 156460
rect 82820 156340 82872 156392
rect 182088 156340 182140 156392
rect 198832 156340 198884 156392
rect 200948 156340 201000 156392
rect 209872 156340 209924 156392
rect 279056 156340 279108 156392
rect 99564 156272 99616 156324
rect 194968 156272 195020 156324
rect 195980 156272 196032 156324
rect 196992 156272 197044 156324
rect 200764 156272 200816 156324
rect 101312 156204 101364 156256
rect 196256 156204 196308 156256
rect 198004 156204 198056 156256
rect 209964 156204 210016 156256
rect 108028 156136 108080 156188
rect 200672 156136 200724 156188
rect 118148 156068 118200 156120
rect 209136 156136 209188 156188
rect 210424 156272 210476 156324
rect 219808 156272 219860 156324
rect 219900 156272 219952 156324
rect 286232 156272 286284 156324
rect 210516 156204 210568 156256
rect 219992 156204 220044 156256
rect 215484 156136 215536 156188
rect 218060 156136 218112 156188
rect 266912 156204 266964 156256
rect 230756 156136 230808 156188
rect 277124 156136 277176 156188
rect 203064 156068 203116 156120
rect 273904 156068 273956 156120
rect 121460 156000 121512 156052
rect 198004 156000 198056 156052
rect 202236 156000 202288 156052
rect 273260 156000 273312 156052
rect 145012 155932 145064 155984
rect 229652 155932 229704 155984
rect 66812 155864 66864 155916
rect 82912 155864 82964 155916
rect 88708 155864 88760 155916
rect 186872 155864 186924 155916
rect 192944 155864 192996 155916
rect 266268 155864 266320 155916
rect 296444 155864 296496 155916
rect 345204 155864 345256 155916
rect 60096 155796 60148 155848
rect 78772 155796 78824 155848
rect 89536 155796 89588 155848
rect 186320 155796 186372 155848
rect 186412 155796 186464 155848
rect 189540 155796 189592 155848
rect 189632 155796 189684 155848
rect 263784 155796 263836 155848
rect 293040 155796 293092 155848
rect 342352 155796 342404 155848
rect 12164 155728 12216 155780
rect 110328 155728 110380 155780
rect 112260 155728 112312 155780
rect 204628 155728 204680 155780
rect 206468 155728 206520 155780
rect 276480 155728 276532 155780
rect 289728 155728 289780 155780
rect 339592 155728 339644 155780
rect 46572 155660 46624 155712
rect 75092 155660 75144 155712
rect 81900 155660 81952 155712
rect 180984 155660 181036 155712
rect 186228 155660 186280 155712
rect 260840 155660 260892 155712
rect 270316 155660 270368 155712
rect 325332 155660 325384 155712
rect 344376 155660 344428 155712
rect 381820 155660 381872 155712
rect 53380 155592 53432 155644
rect 66628 155592 66680 155644
rect 71872 155592 71924 155644
rect 172704 155592 172756 155644
rect 176108 155592 176160 155644
rect 253388 155592 253440 155644
rect 267004 155592 267056 155644
rect 322112 155592 322164 155644
rect 340972 155592 341024 155644
rect 378140 155592 378192 155644
rect 39856 155524 39908 155576
rect 68928 155524 68980 155576
rect 75184 155524 75236 155576
rect 176384 155524 176436 155576
rect 179512 155524 179564 155576
rect 255688 155524 255740 155576
rect 263600 155524 263652 155576
rect 320180 155524 320232 155576
rect 337660 155524 337712 155576
rect 375564 155524 375616 155576
rect 65156 155456 65208 155508
rect 168656 155456 168708 155508
rect 169392 155456 169444 155508
rect 248236 155456 248288 155508
rect 260288 155456 260340 155508
rect 317604 155456 317656 155508
rect 333428 155456 333480 155508
rect 373448 155456 373500 155508
rect 7932 155388 7984 155440
rect 124680 155388 124732 155440
rect 149244 155388 149296 155440
rect 232872 155388 232924 155440
rect 253572 155388 253624 155440
rect 312452 155388 312504 155440
rect 330116 155388 330168 155440
rect 370872 155388 370924 155440
rect 8760 155320 8812 155372
rect 125692 155320 125744 155372
rect 145840 155320 145892 155372
rect 229192 155320 229244 155372
rect 250168 155320 250220 155372
rect 309876 155320 309928 155372
rect 319996 155320 320048 155372
rect 363236 155320 363288 155372
rect 4528 155252 4580 155304
rect 122012 155252 122064 155304
rect 142528 155252 142580 155304
rect 227812 155252 227864 155304
rect 233332 155252 233384 155304
rect 297088 155252 297140 155304
rect 299756 155252 299808 155304
rect 347872 155252 347924 155304
rect 373816 155252 373868 155304
rect 403164 155252 403216 155304
rect 5356 155184 5408 155236
rect 123024 155184 123076 155236
rect 129004 155184 129056 155236
rect 217416 155184 217468 155236
rect 240048 155184 240100 155236
rect 302516 155184 302568 155236
rect 306564 155184 306616 155236
rect 352472 155184 352524 155236
rect 370412 155184 370464 155236
rect 401784 155184 401836 155236
rect 92020 155116 92072 155168
rect 189172 155116 189224 155168
rect 189540 155116 189592 155168
rect 194324 155116 194376 155168
rect 196348 155116 196400 155168
rect 268844 155116 268896 155168
rect 95424 155048 95476 155100
rect 98736 154980 98788 155032
rect 186320 154980 186372 155032
rect 186780 155048 186832 155100
rect 191748 154980 191800 155032
rect 199660 155048 199712 155100
rect 271420 155048 271472 155100
rect 303160 155048 303212 155100
rect 350356 155048 350408 155100
rect 200120 154980 200172 155032
rect 207020 154980 207072 155032
rect 269488 154980 269540 155032
rect 15476 154912 15528 154964
rect 109040 154912 109092 154964
rect 122288 154912 122340 154964
rect 212264 154912 212316 154964
rect 214656 154912 214708 154964
rect 261392 154912 261444 154964
rect 106372 154844 106424 154896
rect 186412 154844 186464 154896
rect 186688 154844 186740 154896
rect 245844 154844 245896 154896
rect 125784 154776 125836 154828
rect 214840 154776 214892 154828
rect 110512 154708 110564 154760
rect 139308 154708 139360 154760
rect 155960 154708 156012 154760
rect 238024 154708 238076 154760
rect 109132 154640 109184 154692
rect 133052 154640 133104 154692
rect 159364 154640 159416 154692
rect 240600 154640 240652 154692
rect 114468 154572 114520 154624
rect 119988 154572 120040 154624
rect 137100 154572 137152 154624
rect 138204 154572 138256 154624
rect 154488 154572 154540 154624
rect 51080 154504 51132 154556
rect 155040 154504 155092 154556
rect 156696 154572 156748 154624
rect 162676 154572 162728 154624
rect 243084 154572 243136 154624
rect 156604 154504 156656 154556
rect 212908 154504 212960 154556
rect 215300 154504 215352 154556
rect 275468 154776 275520 154828
rect 275468 154640 275520 154692
rect 44180 154436 44232 154488
rect 142528 154436 142580 154488
rect 142804 154436 142856 154488
rect 188436 154436 188488 154488
rect 115940 154368 115992 154420
rect 119896 154368 119948 154420
rect 119988 154368 120040 154420
rect 185400 154368 185452 154420
rect 34520 154300 34572 154352
rect 142620 154300 142672 154352
rect 142712 154300 142764 154352
rect 185860 154368 185912 154420
rect 202696 154436 202748 154488
rect 218336 154436 218388 154488
rect 283012 154504 283064 154556
rect 283748 154504 283800 154556
rect 283656 154436 283708 154488
rect 283932 154504 283984 154556
rect 334900 154504 334952 154556
rect 353668 154504 353720 154556
rect 388904 154504 388956 154556
rect 285588 154436 285640 154488
rect 285680 154436 285732 154488
rect 337476 154436 337528 154488
rect 349528 154436 349580 154488
rect 386328 154436 386380 154488
rect 390652 154436 390704 154488
rect 417148 154436 417200 154488
rect 191012 154368 191064 154420
rect 202052 154368 202104 154420
rect 204996 154368 205048 154420
rect 275284 154368 275336 154420
rect 276204 154368 276256 154420
rect 329932 154368 329984 154420
rect 346400 154368 346452 154420
rect 383752 154368 383804 154420
rect 393320 154368 393372 154420
rect 419724 154368 419776 154420
rect 205272 154300 205324 154352
rect 208400 154300 208452 154352
rect 278412 154300 278464 154352
rect 278872 154300 278924 154352
rect 332416 154300 332468 154352
rect 336832 154300 336884 154352
rect 376024 154300 376076 154352
rect 397368 154300 397420 154352
rect 422484 154300 422536 154352
rect 37924 154232 37976 154284
rect 27252 154164 27304 154216
rect 136916 154164 136968 154216
rect 23480 154096 23532 154148
rect 137008 154096 137060 154148
rect 13820 154028 13872 154080
rect 129464 154028 129516 154080
rect 142804 154164 142856 154216
rect 9680 153960 9732 154012
rect 126888 153960 126940 154012
rect 142436 154096 142488 154148
rect 143172 154232 143224 154284
rect 185308 154232 185360 154284
rect 185768 154232 185820 154284
rect 186872 154232 186924 154284
rect 186964 154232 187016 154284
rect 258540 154232 258592 154284
rect 262220 154232 262272 154284
rect 319536 154232 319588 154284
rect 339500 154232 339552 154284
rect 378600 154232 378652 154284
rect 386512 154232 386564 154284
rect 414572 154232 414624 154284
rect 147588 154164 147640 154216
rect 147772 154164 147824 154216
rect 156604 154164 156656 154216
rect 172520 154164 172572 154216
rect 250812 154164 250864 154216
rect 255320 154164 255372 154216
rect 314384 154164 314436 154216
rect 343548 154164 343600 154216
rect 381176 154164 381228 154216
rect 383660 154164 383712 154216
rect 411996 154164 412048 154216
rect 143448 154096 143500 154148
rect 145564 154096 145616 154148
rect 147128 154096 147180 154148
rect 138388 154028 138440 154080
rect 143172 154028 143224 154080
rect 143356 154028 143408 154080
rect 150624 154028 150676 154080
rect 151820 154028 151872 154080
rect 155868 154028 155920 154080
rect 156512 154096 156564 154148
rect 163504 154096 163556 154148
rect 165620 154096 165672 154148
rect 245660 154096 245712 154148
rect 245936 154096 245988 154148
rect 306656 154096 306708 154148
rect 326712 154096 326764 154148
rect 368296 154096 368348 154148
rect 376852 154096 376904 154148
rect 406844 154096 406896 154148
rect 156604 154028 156656 154080
rect 156696 154028 156748 154080
rect 158536 154028 158588 154080
rect 160192 154028 160244 154080
rect 241244 154028 241296 154080
rect 248604 154028 248656 154080
rect 309232 154028 309284 154080
rect 323308 154028 323360 154080
rect 365812 154028 365864 154080
rect 380164 154028 380216 154080
rect 409420 154028 409472 154080
rect 7104 153892 7156 153944
rect 124312 153892 124364 153944
rect 125508 153892 125560 153944
rect 480 153824 532 153876
rect 119804 153824 119856 153876
rect 119896 153824 119948 153876
rect 127716 153892 127768 153944
rect 127808 153892 127860 153944
rect 132408 153892 132460 153944
rect 219900 153960 219952 154012
rect 222384 153960 222436 154012
rect 288716 153960 288768 154012
rect 313280 153960 313332 154012
rect 357900 153960 357952 154012
rect 367100 153960 367152 154012
rect 399116 153960 399168 154012
rect 139860 153892 139912 153944
rect 142436 153892 142488 153944
rect 142528 153892 142580 153944
rect 127624 153824 127676 153876
rect 142804 153824 142856 153876
rect 142988 153892 143040 153944
rect 223212 153892 223264 153944
rect 225236 153892 225288 153944
rect 291292 153892 291344 153944
rect 316040 153892 316092 153944
rect 360660 153892 360712 153944
rect 363052 153892 363104 153944
rect 396540 153892 396592 153944
rect 401600 153892 401652 153944
rect 425520 153892 425572 153944
rect 153292 153824 153344 153876
rect 155040 153824 155092 153876
rect 158352 153824 158404 153876
rect 48320 153756 48372 153808
rect 155776 153756 155828 153808
rect 155868 153756 155920 153808
rect 235448 153824 235500 153876
rect 241888 153824 241940 153876
rect 304080 153824 304132 153876
rect 309140 153824 309192 153876
rect 355508 153824 355560 153876
rect 356244 153824 356296 153876
rect 391480 153824 391532 153876
rect 397460 153824 397512 153876
rect 423036 153824 423088 153876
rect 158536 153756 158588 153808
rect 218060 153756 218112 153808
rect 231860 153756 231912 153808
rect 296444 153756 296496 153808
rect 360384 153756 360436 153808
rect 394056 153756 394108 153808
rect 61108 153688 61160 153740
rect 166080 153688 166132 153740
rect 57980 153620 58032 153672
rect 156512 153620 156564 153672
rect 156604 153620 156656 153672
rect 210424 153688 210476 153740
rect 229100 153688 229152 153740
rect 293868 153688 293920 153740
rect 176660 153620 176712 153672
rect 78680 153552 78732 153604
rect 179604 153552 179656 153604
rect 182180 153620 182232 153672
rect 186964 153620 187016 153672
rect 188436 153620 188488 153672
rect 195980 153620 196032 153672
rect 196072 153620 196124 153672
rect 230940 153552 230992 153604
rect 235080 153620 235132 153672
rect 299020 153620 299072 153672
rect 238668 153552 238720 153604
rect 238852 153552 238904 153604
rect 301596 153552 301648 153604
rect 102140 153484 102192 153536
rect 196900 153484 196952 153536
rect 198924 153484 198976 153536
rect 248880 153484 248932 153536
rect 252652 153484 252704 153536
rect 311808 153484 311860 153536
rect 104900 153416 104952 153468
rect 196532 153416 196584 153468
rect 196992 153416 197044 153468
rect 108304 153348 108356 153400
rect 191012 153348 191064 153400
rect 191656 153348 191708 153400
rect 195888 153348 195940 153400
rect 195980 153348 196032 153400
rect 197544 153348 197596 153400
rect 201408 153416 201460 153468
rect 259184 153416 259236 153468
rect 265440 153416 265492 153468
rect 322020 153416 322072 153468
rect 243728 153348 243780 153400
rect 259460 153348 259512 153400
rect 316960 153348 317012 153400
rect 41604 153280 41656 153332
rect 142712 153280 142764 153332
rect 142804 153280 142856 153332
rect 209780 153280 209832 153332
rect 269212 153280 269264 153332
rect 324688 153280 324740 153332
rect 118700 153212 118752 153264
rect 127624 153212 127676 153264
rect 127716 153212 127768 153264
rect 207848 153212 207900 153264
rect 272892 153212 272944 153264
rect 327264 153212 327316 153264
rect 23296 153144 23348 153196
rect 110972 153144 111024 153196
rect 113180 153144 113232 153196
rect 205916 153144 205968 153196
rect 215392 153144 215444 153196
rect 279700 153144 279752 153196
rect 285496 153144 285548 153196
rect 336832 153144 336884 153196
rect 339684 153144 339736 153196
rect 377312 153144 377364 153196
rect 378232 153144 378284 153196
rect 379888 153144 379940 153196
rect 380992 153144 381044 153196
rect 410064 153144 410116 153196
rect 412916 153144 412968 153196
rect 433800 153144 433852 153196
rect 434352 153144 434404 153196
rect 441620 153144 441672 153196
rect 441712 153144 441764 153196
rect 443000 153144 443052 153196
rect 444196 153144 444248 153196
rect 449256 153144 449308 153196
rect 453948 153144 454000 153196
rect 459468 153144 459520 153196
rect 462228 153144 462280 153196
rect 465908 153144 465960 153196
rect 466460 153144 466512 153196
rect 469772 153144 469824 153196
rect 471336 153144 471388 153196
rect 472992 153144 473044 153196
rect 473360 153144 473412 153196
rect 475568 153144 475620 153196
rect 476120 153144 476172 153196
rect 478144 153144 478196 153196
rect 484032 153144 484084 153196
rect 488448 153144 488500 153196
rect 489920 153144 489972 153196
rect 492864 153144 492916 153196
rect 494060 153144 494112 153196
rect 496084 153144 496136 153196
rect 496636 153144 496688 153196
rect 498016 153144 498068 153196
rect 512276 153144 512328 153196
rect 514852 153144 514904 153196
rect 80060 153076 80112 153128
rect 175096 153076 175148 153128
rect 180800 153076 180852 153128
rect 257252 153076 257304 153128
rect 264980 153076 265032 153128
rect 321468 153076 321520 153128
rect 324320 153076 324372 153128
rect 367008 153076 367060 153128
rect 367192 153076 367244 153128
rect 368940 153076 368992 153128
rect 375472 153076 375524 153128
rect 405556 153076 405608 153128
rect 405832 153076 405884 153128
rect 408776 153076 408828 153128
rect 410800 153076 410852 153128
rect 103520 153008 103572 153060
rect 198188 153008 198240 153060
rect 203708 153008 203760 153060
rect 267556 153008 267608 153060
rect 272156 153008 272208 153060
rect 326620 153008 326672 153060
rect 330944 153008 330996 153060
rect 371516 153008 371568 153060
rect 372620 153008 372672 153060
rect 403532 153008 403584 153060
rect 406660 153008 406712 153060
rect 429200 153008 429252 153060
rect 430672 153076 430724 153128
rect 447968 153076 448020 153128
rect 456984 153076 457036 153128
rect 460756 153076 460808 153128
rect 463516 153076 463568 153128
rect 466552 153076 466604 153128
rect 466644 153076 466696 153128
rect 470416 153076 470468 153128
rect 471428 153076 471480 153128
rect 473636 153076 473688 153128
rect 474832 153076 474884 153128
rect 476856 153076 476908 153128
rect 484952 153076 485004 153128
rect 489644 153076 489696 153128
rect 491668 153076 491720 153128
rect 494796 153076 494848 153128
rect 494980 153076 495032 153128
rect 496728 153076 496780 153128
rect 496820 153076 496872 153128
rect 498660 153076 498712 153128
rect 510988 153076 511040 153128
rect 513472 153076 513524 153128
rect 513564 153076 513616 153128
rect 516140 153076 516192 153128
rect 431224 153008 431276 153060
rect 431960 153008 432012 153060
rect 441712 153008 441764 153060
rect 441804 153008 441856 153060
rect 449900 153008 449952 153060
rect 463608 153008 463660 153060
rect 467288 153008 467340 153060
rect 472440 153008 472492 153060
rect 474924 153008 474976 153060
rect 484400 153008 484452 153060
rect 489000 153008 489052 153060
rect 492680 153008 492732 153060
rect 495440 153008 495492 153060
rect 495532 153008 495584 153060
rect 497372 153008 497424 153060
rect 511632 153008 511684 153060
rect 514300 153008 514352 153060
rect 92572 152940 92624 152992
rect 187884 152940 187936 152992
rect 194600 152940 194652 152992
rect 218704 152940 218756 152992
rect 220360 152940 220412 152992
rect 284852 152940 284904 152992
rect 288072 152940 288124 152992
rect 290004 152940 290056 152992
rect 291384 152940 291436 152992
rect 341340 152940 341392 152992
rect 342260 152940 342312 152992
rect 343916 152940 343968 152992
rect 345296 152940 345348 152992
rect 382464 152940 382516 152992
rect 382556 152940 382608 152992
rect 386972 152940 387024 152992
rect 390376 152940 390428 152992
rect 415216 152940 415268 152992
rect 415400 152940 415452 152992
rect 436376 152940 436428 152992
rect 438860 152940 438912 152992
rect 454408 152940 454460 152992
rect 464712 152940 464764 152992
rect 468392 152940 468444 152992
rect 472532 152940 472584 152992
rect 474280 152940 474332 152992
rect 483112 152940 483164 152992
rect 487804 152940 487856 152992
rect 491300 152940 491352 152992
rect 494152 152940 494204 152992
rect 512920 152940 512972 152992
rect 515956 152940 516008 152992
rect 71412 152872 71464 152924
rect 92480 152872 92532 152924
rect 96620 152872 96672 152924
rect 193036 152872 193088 152924
rect 212448 152872 212500 152924
rect 277768 152872 277820 152924
rect 278780 152872 278832 152924
rect 331772 152872 331824 152924
rect 332600 152872 332652 152924
rect 372804 152872 372856 152924
rect 382188 152872 382240 152924
rect 410708 152872 410760 152924
rect 411260 152872 411312 152924
rect 433156 152872 433208 152924
rect 433524 152872 433576 152924
rect 441712 152872 441764 152924
rect 441896 152872 441948 152924
rect 446956 152872 447008 152924
rect 456800 152872 456852 152924
rect 463332 152872 463384 152924
rect 465080 152872 465132 152924
rect 469128 152872 469180 152924
rect 490012 152872 490064 152924
rect 493508 152872 493560 152924
rect 514208 152872 514260 152924
rect 517428 152872 517480 152924
rect 33140 152804 33192 152856
rect 138020 152804 138072 152856
rect 138112 152804 138164 152856
rect 141700 152804 141752 152856
rect 146484 152804 146536 152856
rect 167368 152804 167420 152856
rect 173900 152804 173952 152856
rect 252100 152804 252152 152856
rect 255412 152804 255464 152856
rect 313096 152804 313148 152856
rect 317052 152804 317104 152856
rect 318248 152804 318300 152856
rect 26424 152736 26476 152788
rect 139124 152736 139176 152788
rect 140780 152736 140832 152788
rect 144276 152736 144328 152788
rect 144368 152736 144420 152788
rect 162216 152736 162268 152788
rect 164424 152736 164476 152788
rect 244372 152736 244424 152788
rect 257712 152736 257764 152788
rect 315672 152736 315724 152788
rect 317420 152736 317472 152788
rect 361304 152804 361356 152856
rect 361580 152804 361632 152856
rect 395252 152804 395304 152856
rect 395528 152804 395580 152856
rect 397828 152804 397880 152856
rect 402428 152804 402480 152856
rect 426164 152804 426216 152856
rect 426440 152804 426492 152856
rect 444748 152804 444800 152856
rect 446312 152804 446364 152856
rect 460112 152804 460164 152856
rect 510344 152804 510396 152856
rect 512000 152804 512052 152856
rect 320272 152736 320324 152788
rect 323124 152736 323176 152788
rect 324228 152736 324280 152788
rect 366364 152736 366416 152788
rect 368480 152736 368532 152788
rect 400404 152736 400456 152788
rect 404360 152736 404412 152788
rect 428004 152736 428056 152788
rect 429384 152736 429436 152788
rect 447324 152736 447376 152788
rect 28172 152668 28224 152720
rect 141056 152668 141108 152720
rect 142804 152668 142856 152720
rect 149428 152668 149480 152720
rect 149520 152668 149572 152720
rect 231584 152668 231636 152720
rect 240232 152668 240284 152720
rect 241888 152668 241940 152720
rect 251180 152668 251232 152720
rect 311164 152668 311216 152720
rect 312176 152668 312228 152720
rect 356152 152668 356204 152720
rect 358820 152668 358872 152720
rect 393412 152668 393464 152720
rect 394884 152668 394936 152720
rect 420368 152668 420420 152720
rect 421012 152668 421064 152720
rect 435364 152668 435416 152720
rect 22192 152600 22244 152652
rect 135904 152600 135956 152652
rect 19340 152532 19392 152584
rect 133972 152532 134024 152584
rect 136640 152532 136692 152584
rect 151912 152600 151964 152652
rect 153568 152600 153620 152652
rect 236736 152600 236788 152652
rect 247040 152600 247092 152652
rect 307944 152600 307996 152652
rect 311532 152600 311584 152652
rect 320640 152600 320692 152652
rect 320824 152600 320876 152652
rect 361948 152600 362000 152652
rect 365720 152600 365772 152652
rect 398472 152600 398524 152652
rect 399208 152600 399260 152652
rect 417424 152600 417476 152652
rect 418620 152600 418672 152652
rect 138112 152532 138164 152584
rect 144276 152532 144328 152584
rect 144368 152532 144420 152584
rect 226432 152532 226484 152584
rect 234160 152532 234212 152584
rect 297732 152532 297784 152584
rect 303620 152532 303672 152584
rect 351000 152532 351052 152584
rect 352012 152532 352064 152584
rect 388260 152532 388312 152584
rect 393136 152532 393188 152584
rect 419080 152532 419132 152584
rect 423404 152600 423456 152652
rect 427084 152600 427136 152652
rect 427820 152600 427872 152652
rect 435456 152600 435508 152652
rect 438952 152668 439004 152720
rect 440240 152668 440292 152720
rect 440516 152668 440568 152720
rect 441620 152668 441672 152720
rect 445208 152668 445260 152720
rect 445300 152668 445352 152720
rect 458916 152668 458968 152720
rect 459652 152668 459704 152720
rect 464620 152668 464672 152720
rect 435640 152600 435692 152652
rect 446036 152600 446088 152652
rect 436192 152532 436244 152584
rect 452476 152532 452528 152584
rect 459560 152532 459612 152584
rect 465264 152532 465316 152584
rect 2872 152464 2924 152516
rect 121092 152464 121144 152516
rect 126980 152464 127032 152516
rect 216128 152464 216180 152516
rect 227720 152464 227772 152516
rect 293224 152464 293276 152516
rect 298652 152464 298704 152516
rect 347136 152464 347188 152516
rect 348148 152464 348200 152516
rect 385040 152464 385092 152516
rect 385500 152464 385552 152516
rect 387616 152464 387668 152516
rect 387708 152464 387760 152516
rect 413928 152464 413980 152516
rect 414296 152464 414348 152516
rect 435732 152464 435784 152516
rect 66628 152396 66680 152448
rect 159640 152396 159692 152448
rect 173256 152396 173308 152448
rect 249524 152396 249576 152448
rect 260932 152396 260984 152448
rect 316316 152396 316368 152448
rect 317512 152396 317564 152448
rect 320732 152396 320784 152448
rect 320824 152396 320876 152448
rect 325976 152396 326028 152448
rect 326068 152396 326120 152448
rect 367652 152396 367704 152448
rect 371332 152396 371384 152448
rect 402336 152396 402388 152448
rect 403900 152396 403952 152448
rect 415860 152396 415912 152448
rect 418160 152396 418212 152448
rect 438308 152464 438360 152516
rect 438400 152464 438452 152516
rect 440884 152464 440936 152516
rect 442080 152464 442132 152516
rect 446680 152464 446732 152516
rect 446772 152464 446824 152516
rect 456984 152464 457036 152516
rect 458180 152464 458232 152516
rect 463976 152464 464028 152516
rect 436100 152396 436152 152448
rect 437112 152396 437164 152448
rect 437756 152396 437808 152448
rect 453120 152396 453172 152448
rect 33600 152328 33652 152380
rect 109684 152328 109736 152380
rect 109776 152328 109828 152380
rect 110512 152328 110564 152380
rect 120080 152328 120132 152380
rect 211068 152328 211120 152380
rect 224408 152328 224460 152380
rect 288072 152328 288124 152380
rect 292212 152328 292264 152380
rect 341984 152328 342036 152380
rect 343824 152328 343876 152380
rect 349804 152328 349856 152380
rect 349896 152328 349948 152380
rect 385684 152328 385736 152380
rect 386420 152328 386472 152380
rect 387708 152328 387760 152380
rect 389180 152328 389232 152380
rect 412640 152328 412692 152380
rect 413836 152328 413888 152380
rect 416504 152328 416556 152380
rect 416596 152328 416648 152380
rect 9496 152260 9548 152312
rect 82820 152260 82872 152312
rect 91100 152260 91152 152312
rect 180248 152260 180300 152312
rect 187976 152260 188028 152312
rect 262404 152260 262456 152312
rect 266360 152260 266412 152312
rect 320916 152260 320968 152312
rect 331220 152260 331272 152312
rect 372160 152260 372212 152312
rect 384948 152260 385000 152312
rect 392124 152260 392176 152312
rect 393688 152260 393740 152312
rect 417792 152260 417844 152312
rect 417884 152260 417936 152312
rect 421748 152260 421800 152312
rect 425980 152328 426032 152380
rect 426808 152260 426860 152312
rect 427084 152328 427136 152380
rect 442172 152328 442224 152380
rect 442816 152328 442868 152380
rect 446772 152328 446824 152380
rect 444104 152260 444156 152312
rect 444196 152260 444248 152312
rect 457628 152328 457680 152380
rect 446956 152260 447008 152312
rect 456340 152260 456392 152312
rect 19800 152192 19852 152244
rect 97908 152192 97960 152244
rect 109040 152192 109092 152244
rect 130752 152192 130804 152244
rect 134064 152192 134116 152244
rect 221280 152192 221332 152244
rect 222108 152192 222160 152244
rect 282920 152192 282972 152244
rect 285772 152192 285824 152244
rect 336188 152192 336240 152244
rect 342444 152192 342496 152244
rect 344560 152192 344612 152244
rect 349160 152192 349212 152244
rect 349896 152192 349948 152244
rect 351920 152192 351972 152244
rect 353484 152192 353536 152244
rect 354496 152192 354548 152244
rect 389548 152192 389600 152244
rect 398104 152192 398156 152244
rect 408132 152192 408184 152244
rect 409236 152192 409288 152244
rect 428648 152192 428700 152244
rect 429292 152192 429344 152244
rect 442080 152192 442132 152244
rect 82912 152124 82964 152176
rect 169944 152124 169996 152176
rect 172152 152124 172204 152176
rect 190460 152124 190512 152176
rect 194140 152124 194192 152176
rect 213552 152124 213604 152176
rect 225328 152124 225380 152176
rect 229008 152124 229060 152176
rect 244464 152124 244516 152176
rect 306012 152124 306064 152176
rect 320640 152124 320692 152176
rect 356796 152124 356848 152176
rect 357532 152124 357584 152176
rect 359372 152124 359424 152176
rect 364524 152124 364576 152176
rect 397184 152124 397236 152176
rect 404636 152124 404688 152176
rect 421012 152124 421064 152176
rect 422576 152124 422628 152176
rect 441528 152124 441580 152176
rect 78772 152056 78824 152108
rect 164792 152056 164844 152108
rect 167000 152056 167052 152108
rect 182732 152056 182784 152108
rect 183468 152056 183520 152108
rect 200764 152056 200816 152108
rect 212724 152056 212776 152108
rect 274548 152056 274600 152108
rect 277400 152056 277452 152108
rect 331128 152056 331180 152108
rect 335360 152056 335412 152108
rect 375380 152056 375432 152108
rect 388444 152056 388496 152108
rect 407488 152056 407540 152108
rect 408500 152056 408552 152108
rect 423588 152056 423640 152108
rect 425152 152056 425204 152108
rect 443460 152192 443512 152244
rect 445208 152192 445260 152244
rect 450544 152192 450596 152244
rect 68928 151988 68980 152040
rect 142804 151988 142856 152040
rect 143264 151988 143316 152040
rect 146944 151988 146996 152040
rect 156788 151988 156840 152040
rect 172520 151988 172572 152040
rect 191472 151988 191524 152040
rect 208492 151988 208544 152040
rect 212632 151988 212684 152040
rect 272708 151988 272760 152040
rect 272800 151988 272852 152040
rect 320824 151988 320876 152040
rect 321560 151988 321612 152040
rect 362592 151988 362644 152040
rect 378784 151988 378836 152040
rect 384396 151988 384448 152040
rect 388352 151988 388404 152040
rect 404912 151988 404964 152040
rect 413744 151988 413796 152040
rect 75092 151920 75144 151972
rect 154488 151920 154540 151972
rect 162492 151920 162544 151972
rect 177672 151920 177724 151972
rect 184388 151920 184440 151972
rect 195612 151920 195664 151972
rect 243360 151920 243412 151972
rect 302884 151920 302936 151972
rect 304172 151920 304224 151972
rect 351644 151920 351696 151972
rect 354680 151920 354732 151972
rect 390192 151920 390244 151972
rect 396172 151920 396224 151972
rect 402980 151920 403032 151972
rect 404268 151920 404320 151972
rect 418436 151920 418488 151972
rect 419540 151988 419592 152040
rect 437020 151988 437072 152040
rect 437112 151988 437164 152040
rect 440240 151988 440292 152040
rect 440332 151988 440384 152040
rect 455696 152124 455748 152176
rect 421656 151920 421708 151972
rect 421748 151920 421800 151972
rect 422852 151920 422904 151972
rect 423496 151920 423548 151972
rect 439596 151920 439648 151972
rect 440516 151920 440568 151972
rect 444472 152056 444524 152108
rect 458180 152056 458232 152108
rect 516692 152056 516744 152108
rect 520280 152056 520332 152108
rect 443736 151988 443788 152040
rect 453764 151988 453816 152040
rect 456892 151988 456944 152040
rect 462688 151988 462740 152040
rect 485780 151988 485832 152040
rect 490288 151988 490340 152040
rect 455052 151920 455104 151972
rect 456064 151920 456116 151972
rect 461400 151920 461452 151972
rect 469220 151920 469272 151972
rect 472348 151920 472400 151972
rect 487344 151920 487396 151972
rect 490932 151920 490984 151972
rect 509056 151920 509108 151972
rect 510896 151920 510948 151972
rect 517428 151920 517480 151972
rect 521568 151920 521620 151972
rect 30196 151852 30248 151904
rect 110328 151852 110380 151904
rect 110512 151852 110564 151904
rect 138480 151852 138532 151904
rect 139308 151852 139360 151904
rect 203340 151852 203392 151904
rect 241612 151852 241664 151904
rect 300952 151852 301004 151904
rect 307392 151852 307444 151904
rect 352288 151852 352340 151904
rect 363144 151852 363196 151904
rect 364524 151852 364576 151904
rect 386144 151852 386196 151904
rect 399760 151852 399812 151904
rect 417424 151852 417476 151904
rect 424140 151852 424192 151904
rect 74816 151784 74868 151836
rect 81348 151784 81400 151836
rect 105820 151784 105872 151836
rect 110236 151784 110288 151836
rect 110420 151784 110472 151836
rect 128176 151784 128228 151836
rect 129740 151784 129792 151836
rect 146852 151784 146904 151836
rect 146944 151784 146996 151836
rect 157064 151784 157116 151836
rect 169760 151784 169812 151836
rect 185308 151784 185360 151836
rect 283196 151784 283248 151836
rect 287428 151784 287480 151836
rect 300400 151784 300452 151836
rect 102324 151716 102376 151768
rect 116124 151716 116176 151768
rect 346492 151784 346544 151836
rect 349804 151784 349856 151836
rect 380532 151784 380584 151836
rect 386236 151784 386288 151836
rect 394700 151784 394752 151836
rect 398840 151784 398892 151836
rect 413284 151784 413336 151836
rect 419632 151784 419684 151836
rect 434444 151852 434496 151904
rect 435364 151852 435416 151904
rect 438400 151852 438452 151904
rect 438584 151852 438636 151904
rect 443552 151852 443604 151904
rect 422852 151716 422904 151768
rect 431776 151784 431828 151836
rect 434720 151784 434772 151836
rect 440056 151784 440108 151836
rect 440240 151784 440292 151836
rect 451832 151852 451884 151904
rect 467840 151852 467892 151904
rect 471060 151852 471112 151904
rect 488540 151852 488592 151904
rect 492220 151852 492272 151904
rect 507768 151852 507820 151904
rect 509516 151852 509568 151904
rect 516048 151852 516100 151904
rect 519452 151852 519504 151904
rect 451096 151784 451148 151836
rect 456156 151784 456208 151836
rect 462044 151784 462096 151836
rect 463884 151784 463936 151836
rect 467748 151784 467800 151836
rect 467932 151784 467984 151836
rect 471704 151784 471756 151836
rect 488172 151784 488224 151836
rect 491576 151784 491628 151836
rect 499120 151784 499172 151836
rect 499948 151784 500000 151836
rect 515496 151784 515548 151836
rect 518900 151784 518952 151836
rect 98920 151648 98972 151700
rect 116032 151648 116084 151700
rect 440148 151648 440200 151700
rect 40500 151580 40552 151632
rect 110972 151580 111024 151632
rect 92020 151512 92072 151564
rect 113088 151512 113140 151564
rect 26700 151444 26752 151496
rect 116952 151444 117004 151496
rect 16396 151376 16448 151428
rect 116768 151376 116820 151428
rect 12992 151308 13044 151360
rect 116676 151308 116728 151360
rect 68008 151240 68060 151292
rect 112720 151240 112772 151292
rect 64512 151172 64564 151224
rect 112628 151172 112680 151224
rect 61108 151104 61160 151156
rect 112536 151104 112588 151156
rect 57704 151036 57756 151088
rect 111708 151036 111760 151088
rect 54208 150968 54260 151020
rect 112444 150968 112496 151020
rect 50804 150900 50856 150952
rect 111616 150900 111668 150952
rect 47308 150832 47360 150884
rect 111524 150832 111576 150884
rect 43904 150764 43956 150816
rect 111432 150764 111484 150816
rect 95516 150696 95568 150748
rect 115296 150696 115348 150748
rect 37004 150628 37056 150680
rect 111248 150628 111300 150680
rect 88616 150560 88668 150612
rect 112996 150560 113048 150612
rect 85212 150492 85264 150544
rect 115204 150492 115256 150544
rect 81716 150424 81768 150476
rect 112904 150424 112956 150476
rect 78312 150288 78364 150340
rect 112812 150288 112864 150340
rect 263692 150288 263744 150340
rect 110328 150220 110380 150272
rect 117136 150220 117188 150272
rect 97908 150152 97960 150204
rect 116860 150152 116912 150204
rect 122840 150152 122892 150204
rect 123714 150152 123766 150204
rect 136916 150152 136968 150204
rect 139814 150152 139866 150204
rect 146392 150152 146444 150204
rect 147542 150152 147594 150204
rect 147680 150152 147732 150204
rect 148830 150152 148882 150204
rect 164332 150152 164384 150204
rect 165482 150152 165534 150204
rect 168472 150152 168524 150204
rect 169346 150152 169398 150204
rect 171140 150152 171192 150204
rect 171922 150152 171974 150204
rect 172704 150152 172756 150204
rect 173854 150152 173906 150204
rect 182272 150152 182324 150204
rect 183422 150152 183474 150204
rect 196532 150152 196584 150204
rect 199522 150152 199574 150204
rect 225052 150152 225104 150204
rect 225834 150152 225886 150204
rect 229192 150152 229244 150204
rect 230342 150152 230394 150204
rect 233240 150152 233292 150204
rect 234206 150152 234258 150204
rect 238944 150152 238996 150204
rect 240002 150152 240054 150204
rect 253940 150152 253992 150204
rect 254722 150152 254774 150204
rect 256792 150152 256844 150204
rect 257942 150152 257994 150204
rect 264382 150152 264434 150204
rect 269120 150152 269172 150204
rect 270178 150152 270230 150204
rect 283104 150152 283156 150204
rect 284254 150152 284306 150204
rect 284392 150152 284444 150204
rect 285542 150152 285594 150204
rect 299480 150152 299532 150204
rect 300354 150152 300406 150204
rect 328460 150152 328512 150204
rect 329242 150152 329294 150204
rect 332692 150152 332744 150204
rect 333750 150152 333802 150204
rect 338396 150152 338448 150204
rect 339454 150152 339506 150204
rect 345112 150152 345164 150204
rect 345894 150152 345946 150204
rect 358912 150152 358964 150204
rect 360062 150152 360114 150204
rect 362960 150152 363012 150204
rect 363926 150152 363978 150204
rect 375564 150152 375616 150204
rect 376714 150152 376766 150204
rect 378140 150152 378192 150204
rect 379290 150152 379342 150204
rect 394976 150152 395028 150204
rect 396034 150152 396086 150204
rect 403164 150152 403216 150204
rect 404314 150152 404366 150204
rect 477684 150152 477736 150204
rect 478834 150152 478886 150204
rect 478972 150152 479024 150204
rect 480122 150152 480174 150204
rect 480260 150152 480312 150204
rect 481410 150152 481462 150204
rect 483204 150152 483256 150204
rect 483986 150152 484038 150204
rect 502340 150152 502392 150204
rect 503214 150152 503266 150204
rect 518026 150152 518078 150204
rect 518808 150152 518860 150204
rect 81348 150084 81400 150136
rect 92480 150084 92532 150136
rect 117228 150084 117280 150136
rect 116492 150016 116544 150068
rect 111156 148316 111208 148368
rect 117044 148316 117096 148368
rect 113088 140700 113140 140752
rect 116124 140700 116176 140752
rect 112996 137912 113048 137964
rect 116124 137912 116176 137964
rect 112904 133832 112956 133884
rect 116032 133832 116084 133884
rect 114192 132608 114244 132660
rect 115204 132608 115256 132660
rect 112812 132404 112864 132456
rect 116124 132404 116176 132456
rect 112720 126896 112772 126948
rect 116124 126896 116176 126948
rect 112628 124108 112680 124160
rect 116124 124108 116176 124160
rect 112536 122748 112588 122800
rect 115940 122748 115992 122800
rect 111708 121388 111760 121440
rect 116124 121388 116176 121440
rect 112444 118600 112496 118652
rect 116124 118600 116176 118652
rect 111616 117240 111668 117292
rect 116124 117240 116176 117292
rect 111524 114452 111576 114504
rect 116124 114452 116176 114504
rect 111432 113092 111484 113144
rect 115940 113092 115992 113144
rect 111340 111732 111392 111784
rect 116124 111732 116176 111784
rect 111156 108944 111208 108996
rect 116124 108944 116176 108996
rect 111248 92420 111300 92472
rect 116124 92420 116176 92472
rect 111064 89632 111116 89684
rect 116124 89632 116176 89684
rect 113824 88272 113876 88324
rect 116032 88272 116084 88324
rect 113916 83920 113968 83972
rect 116584 83920 116636 83972
rect 114008 82764 114060 82816
rect 116216 82764 116268 82816
rect 114100 79976 114152 80028
rect 115940 79976 115992 80028
rect 114192 78616 114244 78668
rect 116124 78616 116176 78668
rect 114192 71748 114244 71800
rect 116584 71748 116636 71800
rect 114100 69028 114152 69080
rect 116308 69028 116360 69080
rect 114008 67600 114060 67652
rect 116124 67600 116176 67652
rect 113916 66240 113968 66292
rect 116584 66240 116636 66292
rect 113364 64676 113416 64728
rect 116584 64676 116636 64728
rect 113824 63520 113876 63572
rect 116216 63520 116268 63572
rect 112444 62092 112496 62144
rect 116124 62092 116176 62144
rect 112536 42780 112588 42832
rect 116124 42780 116176 42832
rect 116676 7896 116728 7948
rect 116860 7896 116912 7948
rect 117044 7760 117096 7812
rect 117320 7760 117372 7812
rect 116860 7692 116912 7744
rect 116768 7624 116820 7676
rect 117228 7624 117280 7676
rect 117044 7420 117096 7472
rect 111708 2864 111760 2916
rect 111800 2796 111852 2848
rect 170312 2456 170364 2508
rect 193588 2456 193640 2508
rect 294788 2456 294840 2508
rect 425796 2456 425848 2508
rect 443644 2456 443696 2508
rect 170312 2320 170364 2372
rect 62396 1844 62448 1896
rect 65340 1844 65392 1896
rect 68008 1844 68060 1896
rect 77116 1844 77168 1896
rect 77760 1844 77812 1896
rect 89260 1844 89312 1896
rect 89352 1844 89404 1896
rect 99656 1844 99708 1896
rect 104348 1844 104400 1896
rect 64144 1776 64196 1828
rect 69388 1776 69440 1828
rect 77024 1776 77076 1828
rect 85948 1776 86000 1828
rect 86040 1776 86092 1828
rect 111064 1912 111116 1964
rect 104532 1844 104584 1896
rect 105728 1844 105780 1896
rect 105820 1844 105872 1896
rect 105912 1844 105964 1896
rect 109224 1844 109276 1896
rect 109316 1844 109368 1896
rect 62672 1708 62724 1760
rect 68836 1708 68888 1760
rect 79968 1708 80020 1760
rect 80796 1708 80848 1760
rect 82636 1708 82688 1760
rect 104072 1708 104124 1760
rect 109592 1776 109644 1828
rect 109960 1708 110012 1760
rect 112444 1708 112496 1760
rect 69296 1640 69348 1692
rect 102600 1640 102652 1692
rect 102692 1640 102744 1692
rect 105820 1640 105872 1692
rect 106188 1640 106240 1692
rect 116584 1640 116636 1692
rect 59360 1572 59412 1624
rect 68468 1572 68520 1624
rect 79324 1572 79376 1624
rect 99472 1572 99524 1624
rect 99564 1572 99616 1624
rect 105912 1572 105964 1624
rect 106004 1572 106056 1624
rect 110144 1572 110196 1624
rect 72700 1504 72752 1556
rect 42616 1436 42668 1488
rect 80428 1436 80480 1488
rect 94136 1436 94188 1488
rect 96620 1436 96672 1488
rect 110512 1504 110564 1556
rect 99656 1436 99708 1488
rect 108212 1436 108264 1488
rect 108304 1436 108356 1488
rect 143632 1436 143684 1488
rect 46020 1368 46072 1420
rect 116492 1368 116544 1420
rect 294788 1368 294840 1420
rect 343640 1368 343692 1420
rect 491300 1368 491352 1420
rect 493600 1368 493652 1420
rect 2688 1300 2740 1352
rect 116308 1300 116360 1352
rect 39304 1232 39356 1284
rect 116400 1232 116452 1284
rect 49332 1164 49384 1216
rect 116768 1164 116820 1216
rect 52644 1096 52696 1148
rect 117228 1096 117280 1148
rect 55956 1028 56008 1080
rect 111800 1028 111852 1080
rect 65984 960 66036 1012
rect 116860 960 116912 1012
rect 76012 892 76064 944
rect 112536 892 112588 944
rect 94688 824 94740 876
rect 100116 824 100168 876
rect 96344 756 96396 808
rect 101864 756 101916 808
<< metal2 >>
rect 386 163200 442 164400
rect 492 163254 1164 163282
rect 400 158030 428 163200
rect 388 158024 440 158030
rect 388 157966 440 157972
rect 492 153882 520 163254
rect 1136 163146 1164 163254
rect 1214 163200 1270 164400
rect 2042 163200 2098 164400
rect 2870 163200 2926 164400
rect 2976 163254 3648 163282
rect 1228 163146 1256 163200
rect 1136 163118 1256 163146
rect 2056 156670 2084 163200
rect 2044 156664 2096 156670
rect 2044 156606 2096 156612
rect 480 153876 532 153882
rect 480 153818 532 153824
rect 2884 152522 2912 163200
rect 2976 153785 3004 163254
rect 3620 163146 3648 163254
rect 3698 163200 3754 164400
rect 4526 163200 4582 164400
rect 5354 163200 5410 164400
rect 6274 163200 6330 164400
rect 7102 163200 7158 164400
rect 7930 163200 7986 164400
rect 8758 163200 8814 164400
rect 8864 163254 9536 163282
rect 3712 163146 3740 163200
rect 3620 163118 3740 163146
rect 4540 155310 4568 163200
rect 4528 155304 4580 155310
rect 4528 155246 4580 155252
rect 5368 155242 5396 163200
rect 6288 159390 6316 163200
rect 6276 159384 6328 159390
rect 6276 159326 6328 159332
rect 5356 155236 5408 155242
rect 5356 155178 5408 155184
rect 7116 153950 7144 163200
rect 7944 155446 7972 163200
rect 7932 155440 7984 155446
rect 7932 155382 7984 155388
rect 8772 155378 8800 163200
rect 8760 155372 8812 155378
rect 8760 155314 8812 155320
rect 7104 153944 7156 153950
rect 7104 153886 7156 153892
rect 2962 153776 3018 153785
rect 2962 153711 3018 153720
rect 2872 152516 2924 152522
rect 2872 152458 2924 152464
rect 8864 152425 8892 163254
rect 9508 163146 9536 163254
rect 9586 163200 9642 164400
rect 9692 163254 10364 163282
rect 9600 163146 9628 163200
rect 9508 163118 9628 163146
rect 9692 154018 9720 163254
rect 10336 163146 10364 163254
rect 10414 163200 10470 164400
rect 11242 163200 11298 164400
rect 12162 163200 12218 164400
rect 12452 163254 12940 163282
rect 10428 163146 10456 163200
rect 10336 163118 10456 163146
rect 11256 156738 11284 163200
rect 11244 156732 11296 156738
rect 11244 156674 11296 156680
rect 12176 155786 12204 163200
rect 12164 155780 12216 155786
rect 12164 155722 12216 155728
rect 9680 154012 9732 154018
rect 9680 153954 9732 153960
rect 12452 152561 12480 163254
rect 12912 163146 12940 163254
rect 12990 163200 13046 164400
rect 13818 163200 13874 164400
rect 14646 163200 14702 164400
rect 15474 163200 15530 164400
rect 16302 163200 16358 164400
rect 16592 163254 17080 163282
rect 13004 163146 13032 163200
rect 12912 163118 13032 163146
rect 13832 154086 13860 163200
rect 14660 156806 14688 163200
rect 14648 156800 14700 156806
rect 14648 156742 14700 156748
rect 15488 154970 15516 163200
rect 16316 159361 16344 163200
rect 16302 159352 16358 159361
rect 16302 159287 16358 159296
rect 15476 154964 15528 154970
rect 15476 154906 15528 154912
rect 13820 154080 13872 154086
rect 13820 154022 13872 154028
rect 16592 153921 16620 163254
rect 17052 163146 17080 163254
rect 17130 163200 17186 164400
rect 18050 163200 18106 164400
rect 18878 163200 18934 164400
rect 19352 163254 19656 163282
rect 17144 163146 17172 163200
rect 17052 163118 17172 163146
rect 18064 156874 18092 163200
rect 18892 159730 18920 163200
rect 18880 159724 18932 159730
rect 18880 159666 18932 159672
rect 18052 156868 18104 156874
rect 18052 156810 18104 156816
rect 16578 153912 16634 153921
rect 16578 153847 16634 153856
rect 19352 152590 19380 163254
rect 19628 163146 19656 163254
rect 19706 163200 19762 164400
rect 19904 163254 20484 163282
rect 19720 163146 19748 163200
rect 19628 163118 19748 163146
rect 19904 154057 19932 163254
rect 20456 163146 20484 163254
rect 20534 163200 20590 164400
rect 21362 163200 21418 164400
rect 22190 163200 22246 164400
rect 23018 163200 23074 164400
rect 23492 163254 23888 163282
rect 20548 163146 20576 163200
rect 20456 163118 20576 163146
rect 21376 156942 21404 163200
rect 21364 156936 21416 156942
rect 21364 156878 21416 156884
rect 19890 154048 19946 154057
rect 19890 153983 19946 153992
rect 22204 152658 22232 163200
rect 23032 159497 23060 163200
rect 23018 159488 23074 159497
rect 23018 159423 23074 159432
rect 23492 154154 23520 163254
rect 23860 163146 23888 163254
rect 23938 163200 23994 164400
rect 24766 163200 24822 164400
rect 25594 163200 25650 164400
rect 26422 163200 26478 164400
rect 27250 163200 27306 164400
rect 28078 163200 28134 164400
rect 28184 163254 28856 163282
rect 23952 163146 23980 163200
rect 23860 163118 23980 163146
rect 24780 157010 24808 163200
rect 25608 160002 25636 163200
rect 25596 159996 25648 160002
rect 25596 159938 25648 159944
rect 24768 157004 24820 157010
rect 24768 156946 24820 156952
rect 23480 154148 23532 154154
rect 23480 154090 23532 154096
rect 23296 153196 23348 153202
rect 23296 153138 23348 153144
rect 22192 152652 22244 152658
rect 22192 152594 22244 152600
rect 19340 152584 19392 152590
rect 12438 152552 12494 152561
rect 19340 152526 19392 152532
rect 12438 152487 12494 152496
rect 8850 152416 8906 152425
rect 8850 152351 8906 152360
rect 9496 152312 9548 152318
rect 9496 152254 9548 152260
rect 6090 150648 6146 150657
rect 6090 150583 6146 150592
rect 2686 150512 2742 150521
rect 2686 150447 2742 150456
rect 2700 149940 2728 150447
rect 6104 149940 6132 150583
rect 9508 149940 9536 152254
rect 19800 152244 19852 152250
rect 19800 152186 19852 152192
rect 16396 151428 16448 151434
rect 16396 151370 16448 151376
rect 12992 151360 13044 151366
rect 12992 151302 13044 151308
rect 13004 149940 13032 151302
rect 16408 149940 16436 151370
rect 19812 149940 19840 152186
rect 23308 149940 23336 153138
rect 26436 152794 26464 163200
rect 27264 154222 27292 163200
rect 28092 156641 28120 163200
rect 28078 156632 28134 156641
rect 28078 156567 28134 156576
rect 27252 154216 27304 154222
rect 27252 154158 27304 154164
rect 26424 152788 26476 152794
rect 26424 152730 26476 152736
rect 28184 152726 28212 163254
rect 28828 163146 28856 163254
rect 28906 163200 28962 164400
rect 29826 163200 29882 164400
rect 30392 163254 30604 163282
rect 28920 163146 28948 163200
rect 28828 163118 28948 163146
rect 29840 159633 29868 163200
rect 29826 159624 29882 159633
rect 29826 159559 29882 159568
rect 30392 154193 30420 163254
rect 30576 163146 30604 163254
rect 30654 163200 30710 164400
rect 31482 163200 31538 164400
rect 32310 163200 32366 164400
rect 33138 163200 33194 164400
rect 33966 163200 34022 164400
rect 34532 163254 34744 163282
rect 30668 163146 30696 163200
rect 30576 163118 30696 163146
rect 31496 156777 31524 163200
rect 32324 159526 32352 163200
rect 32312 159520 32364 159526
rect 32312 159462 32364 159468
rect 31482 156768 31538 156777
rect 31482 156703 31538 156712
rect 30378 154184 30434 154193
rect 30378 154119 30434 154128
rect 33152 152862 33180 163200
rect 33980 158001 34008 163200
rect 33966 157992 34022 158001
rect 33966 157927 34022 157936
rect 34532 154358 34560 163254
rect 34716 163146 34744 163254
rect 34794 163200 34850 164400
rect 35714 163200 35770 164400
rect 36542 163200 36598 164400
rect 37370 163200 37426 164400
rect 37936 163254 38148 163282
rect 34808 163146 34836 163200
rect 34716 163118 34836 163146
rect 35728 157078 35756 163200
rect 36556 159458 36584 163200
rect 36544 159452 36596 159458
rect 36544 159394 36596 159400
rect 37384 158098 37412 163200
rect 37372 158092 37424 158098
rect 37372 158034 37424 158040
rect 35716 157072 35768 157078
rect 35716 157014 35768 157020
rect 34520 154352 34572 154358
rect 34520 154294 34572 154300
rect 37936 154290 37964 163254
rect 38120 163146 38148 163254
rect 38198 163200 38254 164400
rect 39026 163200 39082 164400
rect 39854 163200 39910 164400
rect 40682 163200 40738 164400
rect 41602 163200 41658 164400
rect 42430 163200 42486 164400
rect 43258 163200 43314 164400
rect 44086 163200 44142 164400
rect 44192 163254 44864 163282
rect 38212 163146 38240 163200
rect 38120 163118 38240 163146
rect 39040 157146 39068 163200
rect 39028 157140 39080 157146
rect 39028 157082 39080 157088
rect 39868 155582 39896 163200
rect 40696 158273 40724 163200
rect 40682 158264 40738 158273
rect 40682 158199 40738 158208
rect 39856 155576 39908 155582
rect 39856 155518 39908 155524
rect 37924 154284 37976 154290
rect 37924 154226 37976 154232
rect 41616 153338 41644 163200
rect 42444 157214 42472 163200
rect 43272 159594 43300 163200
rect 43260 159588 43312 159594
rect 43260 159530 43312 159536
rect 44100 158137 44128 163200
rect 44086 158128 44142 158137
rect 44086 158063 44142 158072
rect 42432 157208 42484 157214
rect 42432 157150 42484 157156
rect 44192 154494 44220 163254
rect 44836 163146 44864 163254
rect 44914 163200 44970 164400
rect 45742 163200 45798 164400
rect 46570 163200 46626 164400
rect 47490 163200 47546 164400
rect 48318 163200 48374 164400
rect 49146 163200 49202 164400
rect 49974 163200 50030 164400
rect 50802 163200 50858 164400
rect 51092 163254 51580 163282
rect 44928 163146 44956 163200
rect 44836 163118 44956 163146
rect 45756 157282 45784 163200
rect 45744 157276 45796 157282
rect 45744 157218 45796 157224
rect 46584 155718 46612 163200
rect 47504 158166 47532 163200
rect 47492 158160 47544 158166
rect 47492 158102 47544 158108
rect 46572 155712 46624 155718
rect 46572 155654 46624 155660
rect 44180 154488 44232 154494
rect 44180 154430 44232 154436
rect 48332 153814 48360 163200
rect 49160 157350 49188 163200
rect 49988 159662 50016 163200
rect 49976 159656 50028 159662
rect 49976 159598 50028 159604
rect 50816 158234 50844 163200
rect 50804 158228 50856 158234
rect 50804 158170 50856 158176
rect 49148 157344 49200 157350
rect 49148 157286 49200 157292
rect 51092 154562 51120 163254
rect 51552 163146 51580 163254
rect 51630 163200 51686 164400
rect 52458 163200 52514 164400
rect 53378 163200 53434 164400
rect 54206 163200 54262 164400
rect 54312 163254 54984 163282
rect 51644 163146 51672 163200
rect 51552 163118 51672 163146
rect 52472 156602 52500 163200
rect 52460 156596 52512 156602
rect 52460 156538 52512 156544
rect 53392 155650 53420 163200
rect 54220 158302 54248 163200
rect 54208 158296 54260 158302
rect 54208 158238 54260 158244
rect 53380 155644 53432 155650
rect 53380 155586 53432 155592
rect 51080 154556 51132 154562
rect 51080 154498 51132 154504
rect 54312 154329 54340 163254
rect 54956 163146 54984 163254
rect 55034 163200 55090 164400
rect 55862 163200 55918 164400
rect 56690 163200 56746 164400
rect 57518 163200 57574 164400
rect 57992 163254 58296 163282
rect 55048 163146 55076 163200
rect 54956 163118 55076 163146
rect 55876 156913 55904 163200
rect 56704 159798 56732 163200
rect 56692 159792 56744 159798
rect 56692 159734 56744 159740
rect 57532 158409 57560 163200
rect 57518 158400 57574 158409
rect 57518 158335 57574 158344
rect 55862 156904 55918 156913
rect 55862 156839 55918 156848
rect 54298 154320 54354 154329
rect 54298 154255 54354 154264
rect 48320 153808 48372 153814
rect 48320 153750 48372 153756
rect 57992 153678 58020 163254
rect 58268 163146 58296 163254
rect 58346 163200 58402 164400
rect 59266 163200 59322 164400
rect 60094 163200 60150 164400
rect 60922 163200 60978 164400
rect 61120 163254 61700 163282
rect 58360 163146 58388 163200
rect 58268 163118 58388 163146
rect 59280 156534 59308 163200
rect 59268 156528 59320 156534
rect 59268 156470 59320 156476
rect 60108 155854 60136 163200
rect 60936 158370 60964 163200
rect 60924 158364 60976 158370
rect 60924 158306 60976 158312
rect 60096 155848 60148 155854
rect 60096 155790 60148 155796
rect 61120 153746 61148 163254
rect 61672 163146 61700 163254
rect 61750 163200 61806 164400
rect 62578 163200 62634 164400
rect 63406 163200 63462 164400
rect 64234 163200 64290 164400
rect 65154 163200 65210 164400
rect 65982 163200 66038 164400
rect 66810 163200 66866 164400
rect 67638 163200 67694 164400
rect 68466 163200 68522 164400
rect 69294 163200 69350 164400
rect 70122 163200 70178 164400
rect 71042 163200 71098 164400
rect 71870 163200 71926 164400
rect 72698 163200 72754 164400
rect 73526 163200 73582 164400
rect 74354 163200 74410 164400
rect 75182 163200 75238 164400
rect 76010 163200 76066 164400
rect 76930 163200 76986 164400
rect 77758 163200 77814 164400
rect 78586 163200 78642 164400
rect 78692 163254 79364 163282
rect 61764 163146 61792 163200
rect 61672 163118 61792 163146
rect 62592 155417 62620 163200
rect 63420 160070 63448 163200
rect 63408 160064 63460 160070
rect 63408 160006 63460 160012
rect 64248 158438 64276 163200
rect 64236 158432 64288 158438
rect 64236 158374 64288 158380
rect 65168 155514 65196 163200
rect 65996 155553 66024 163200
rect 66824 155922 66852 163200
rect 67652 158642 67680 163200
rect 67640 158636 67692 158642
rect 67640 158578 67692 158584
rect 66812 155916 66864 155922
rect 66812 155858 66864 155864
rect 66628 155644 66680 155650
rect 66628 155586 66680 155592
rect 65982 155544 66038 155553
rect 65156 155508 65208 155514
rect 65982 155479 66038 155488
rect 65156 155450 65208 155456
rect 62578 155408 62634 155417
rect 62578 155343 62634 155352
rect 61108 153740 61160 153746
rect 61108 153682 61160 153688
rect 57980 153672 58032 153678
rect 57980 153614 58032 153620
rect 41604 153332 41656 153338
rect 41604 153274 41656 153280
rect 33140 152856 33192 152862
rect 33140 152798 33192 152804
rect 28172 152720 28224 152726
rect 28172 152662 28224 152668
rect 66640 152454 66668 155586
rect 68480 155281 68508 163200
rect 69308 156466 69336 163200
rect 70136 159866 70164 163200
rect 70124 159860 70176 159866
rect 70124 159802 70176 159808
rect 71056 158506 71084 163200
rect 71044 158500 71096 158506
rect 71044 158442 71096 158448
rect 69296 156460 69348 156466
rect 69296 156402 69348 156408
rect 71884 155650 71912 163200
rect 72712 157049 72740 163200
rect 73540 159322 73568 163200
rect 73528 159316 73580 159322
rect 73528 159258 73580 159264
rect 74368 158574 74396 163200
rect 74356 158568 74408 158574
rect 74356 158510 74408 158516
rect 72698 157040 72754 157049
rect 72698 156975 72754 156984
rect 75092 155712 75144 155718
rect 75092 155654 75144 155660
rect 71872 155644 71924 155650
rect 71872 155586 71924 155592
rect 68928 155576 68980 155582
rect 68928 155518 68980 155524
rect 68466 155272 68522 155281
rect 68466 155207 68522 155216
rect 66628 152448 66680 152454
rect 66628 152390 66680 152396
rect 33600 152380 33652 152386
rect 33600 152322 33652 152328
rect 30196 151904 30248 151910
rect 30196 151846 30248 151852
rect 26700 151496 26752 151502
rect 26700 151438 26752 151444
rect 26712 149940 26740 151438
rect 30208 149940 30236 151846
rect 33612 149940 33640 152322
rect 68940 152046 68968 155518
rect 71412 152924 71464 152930
rect 71412 152866 71464 152872
rect 68928 152040 68980 152046
rect 68928 151982 68980 151988
rect 40500 151632 40552 151638
rect 40500 151574 40552 151580
rect 37004 150680 37056 150686
rect 37004 150622 37056 150628
rect 37016 149940 37044 150622
rect 40512 149940 40540 151574
rect 68008 151292 68060 151298
rect 68008 151234 68060 151240
rect 64512 151224 64564 151230
rect 64512 151166 64564 151172
rect 61108 151156 61160 151162
rect 61108 151098 61160 151104
rect 57704 151088 57756 151094
rect 57704 151030 57756 151036
rect 54208 151020 54260 151026
rect 54208 150962 54260 150968
rect 50804 150952 50856 150958
rect 50804 150894 50856 150900
rect 47308 150884 47360 150890
rect 47308 150826 47360 150832
rect 43904 150816 43956 150822
rect 43904 150758 43956 150764
rect 43916 149940 43944 150758
rect 47320 149940 47348 150826
rect 50816 149940 50844 150894
rect 54220 149940 54248 150962
rect 57716 149940 57744 151030
rect 61120 149940 61148 151098
rect 64524 149940 64552 151166
rect 68020 149940 68048 151234
rect 71424 149940 71452 152866
rect 75104 151978 75132 155654
rect 75196 155582 75224 163200
rect 76024 155825 76052 163200
rect 76944 159934 76972 163200
rect 76932 159928 76984 159934
rect 76932 159870 76984 159876
rect 77772 157962 77800 163200
rect 77760 157956 77812 157962
rect 77760 157898 77812 157904
rect 76010 155816 76066 155825
rect 76010 155751 76066 155760
rect 78600 155689 78628 163200
rect 78586 155680 78642 155689
rect 78586 155615 78642 155624
rect 75184 155576 75236 155582
rect 75184 155518 75236 155524
rect 78692 153610 78720 163254
rect 79336 163146 79364 163254
rect 79414 163200 79470 164400
rect 80242 163200 80298 164400
rect 81070 163200 81126 164400
rect 81898 163200 81954 164400
rect 82818 163200 82874 164400
rect 83646 163200 83702 164400
rect 84474 163200 84530 164400
rect 85302 163200 85358 164400
rect 85592 163254 86080 163282
rect 79428 163146 79456 163200
rect 79336 163118 79456 163146
rect 80060 159316 80112 159322
rect 80060 159258 80112 159264
rect 78772 155848 78824 155854
rect 78772 155790 78824 155796
rect 78680 153604 78732 153610
rect 78680 153546 78732 153552
rect 78784 152114 78812 155790
rect 80072 153134 80100 159258
rect 80256 159254 80284 163200
rect 80244 159248 80296 159254
rect 80244 159190 80296 159196
rect 81084 158710 81112 163200
rect 81072 158704 81124 158710
rect 81072 158646 81124 158652
rect 81912 155718 81940 163200
rect 82832 156398 82860 163200
rect 83660 159322 83688 163200
rect 83648 159316 83700 159322
rect 83648 159258 83700 159264
rect 84488 157826 84516 163200
rect 84476 157820 84528 157826
rect 84476 157762 84528 157768
rect 82820 156392 82872 156398
rect 82820 156334 82872 156340
rect 85316 155961 85344 163200
rect 85302 155952 85358 155961
rect 82912 155916 82964 155922
rect 85302 155887 85358 155896
rect 82912 155858 82964 155864
rect 81900 155712 81952 155718
rect 81900 155654 81952 155660
rect 80060 153128 80112 153134
rect 80060 153070 80112 153076
rect 82820 152312 82872 152318
rect 82820 152254 82872 152260
rect 78772 152108 78824 152114
rect 78772 152050 78824 152056
rect 75092 151972 75144 151978
rect 75092 151914 75144 151920
rect 74816 151836 74868 151842
rect 81348 151836 81400 151842
rect 74868 151786 74948 151814
rect 74816 151778 74868 151784
rect 74920 149954 74948 151786
rect 81348 151778 81400 151784
rect 78312 150340 78364 150346
rect 78312 150282 78364 150288
rect 74842 149926 74948 149954
rect 78324 149940 78352 150282
rect 81360 150142 81388 151778
rect 81716 150476 81768 150482
rect 81716 150418 81768 150424
rect 81348 150136 81400 150142
rect 81348 150078 81400 150084
rect 81728 149940 81756 150418
rect 82832 149705 82860 152254
rect 82924 152182 82952 155858
rect 85592 154465 85620 163254
rect 86052 163146 86080 163254
rect 86130 163200 86186 164400
rect 86958 163200 87014 164400
rect 87786 163200 87842 164400
rect 88706 163200 88762 164400
rect 89534 163200 89590 164400
rect 90362 163200 90418 164400
rect 91190 163200 91246 164400
rect 92018 163200 92074 164400
rect 92846 163200 92902 164400
rect 93674 163200 93730 164400
rect 94594 163200 94650 164400
rect 95422 163200 95478 164400
rect 96250 163200 96306 164400
rect 96632 163254 97028 163282
rect 86144 163146 86172 163200
rect 86052 163118 86172 163146
rect 86972 159186 87000 163200
rect 86960 159180 87012 159186
rect 86960 159122 87012 159128
rect 87800 157894 87828 163200
rect 87788 157888 87840 157894
rect 87788 157830 87840 157836
rect 88720 155922 88748 163200
rect 88708 155916 88760 155922
rect 88708 155858 88760 155864
rect 89548 155854 89576 163200
rect 90376 158778 90404 163200
rect 91100 159248 91152 159254
rect 91100 159190 91152 159196
rect 90364 158772 90416 158778
rect 90364 158714 90416 158720
rect 89536 155848 89588 155854
rect 89536 155790 89588 155796
rect 85578 154456 85634 154465
rect 85578 154391 85634 154400
rect 91112 152318 91140 159190
rect 91204 157758 91232 163200
rect 91192 157752 91244 157758
rect 91192 157694 91244 157700
rect 92032 155174 92060 163200
rect 92860 158778 92888 163200
rect 93688 159118 93716 163200
rect 93676 159112 93728 159118
rect 93676 159054 93728 159060
rect 92572 158772 92624 158778
rect 92572 158714 92624 158720
rect 92848 158772 92900 158778
rect 92848 158714 92900 158720
rect 92020 155168 92072 155174
rect 92020 155110 92072 155116
rect 92584 152998 92612 158714
rect 94608 157690 94636 163200
rect 94596 157684 94648 157690
rect 94596 157626 94648 157632
rect 95436 155106 95464 163200
rect 96264 158982 96292 163200
rect 96252 158976 96304 158982
rect 96252 158918 96304 158924
rect 95424 155100 95476 155106
rect 95424 155042 95476 155048
rect 92572 152992 92624 152998
rect 92572 152934 92624 152940
rect 96632 152930 96660 163254
rect 97000 163146 97028 163254
rect 97078 163200 97134 164400
rect 97906 163200 97962 164400
rect 98734 163200 98790 164400
rect 99562 163200 99618 164400
rect 100482 163200 100538 164400
rect 101310 163200 101366 164400
rect 102138 163200 102194 164400
rect 102966 163200 103022 164400
rect 103532 163254 103744 163282
rect 97092 163146 97120 163200
rect 97000 163118 97120 163146
rect 97920 157622 97948 163200
rect 97908 157616 97960 157622
rect 97908 157558 97960 157564
rect 98748 155038 98776 163200
rect 99576 156330 99604 163200
rect 100496 159254 100524 163200
rect 100484 159248 100536 159254
rect 100484 159190 100536 159196
rect 99564 156324 99616 156330
rect 99564 156266 99616 156272
rect 101324 156262 101352 163200
rect 101312 156256 101364 156262
rect 101312 156198 101364 156204
rect 98736 155032 98788 155038
rect 98736 154974 98788 154980
rect 102152 153542 102180 163200
rect 102980 158914 103008 163200
rect 102968 158908 103020 158914
rect 102968 158850 103020 158856
rect 102140 153536 102192 153542
rect 102140 153478 102192 153484
rect 103532 153066 103560 163254
rect 103716 163146 103744 163254
rect 103794 163200 103850 164400
rect 104622 163200 104678 164400
rect 104912 163254 105400 163282
rect 103808 163146 103836 163200
rect 103716 163118 103836 163146
rect 104636 158545 104664 163200
rect 104622 158536 104678 158545
rect 104622 158471 104678 158480
rect 104912 153474 104940 163254
rect 105372 163146 105400 163254
rect 105450 163200 105506 164400
rect 106370 163200 106426 164400
rect 107198 163200 107254 164400
rect 108026 163200 108082 164400
rect 108316 163254 108804 163282
rect 105464 163146 105492 163200
rect 105372 163118 105492 163146
rect 106384 154902 106412 163200
rect 107212 159050 107240 163200
rect 107200 159044 107252 159050
rect 107200 158986 107252 158992
rect 108040 156194 108068 163200
rect 108028 156188 108080 156194
rect 108028 156130 108080 156136
rect 106372 154896 106424 154902
rect 106372 154838 106424 154844
rect 104900 153468 104952 153474
rect 104900 153410 104952 153416
rect 108316 153406 108344 163254
rect 108776 163146 108804 163254
rect 108854 163200 108910 164400
rect 109682 163200 109738 164400
rect 110510 163200 110566 164400
rect 111338 163200 111394 164400
rect 112258 163200 112314 164400
rect 113086 163200 113142 164400
rect 113192 163254 113864 163282
rect 108868 163146 108896 163200
rect 108776 163118 108896 163146
rect 109132 159724 109184 159730
rect 109132 159666 109184 159672
rect 109040 154964 109092 154970
rect 109040 154906 109092 154912
rect 108304 153400 108356 153406
rect 108304 153342 108356 153348
rect 103520 153060 103572 153066
rect 103520 153002 103572 153008
rect 92480 152924 92532 152930
rect 92480 152866 92532 152872
rect 96620 152924 96672 152930
rect 96620 152866 96672 152872
rect 91100 152312 91152 152318
rect 91100 152254 91152 152260
rect 82912 152176 82964 152182
rect 82912 152118 82964 152124
rect 92020 151564 92072 151570
rect 92020 151506 92072 151512
rect 88616 150612 88668 150618
rect 88616 150554 88668 150560
rect 85212 150544 85264 150550
rect 85212 150486 85264 150492
rect 85224 149940 85252 150486
rect 88628 149940 88656 150554
rect 92032 149940 92060 151506
rect 92492 150142 92520 152866
rect 109052 152250 109080 154906
rect 109144 154698 109172 159666
rect 109696 158846 109724 163200
rect 109776 159996 109828 160002
rect 109776 159938 109828 159944
rect 109684 158840 109736 158846
rect 109684 158782 109736 158788
rect 109132 154692 109184 154698
rect 109132 154634 109184 154640
rect 109788 152386 109816 159938
rect 110328 155780 110380 155786
rect 110328 155722 110380 155728
rect 109684 152380 109736 152386
rect 109684 152322 109736 152328
rect 109776 152380 109828 152386
rect 109776 152322 109828 152328
rect 97908 152244 97960 152250
rect 97908 152186 97960 152192
rect 109040 152244 109092 152250
rect 109040 152186 109092 152192
rect 95516 150748 95568 150754
rect 95516 150690 95568 150696
rect 92480 150136 92532 150142
rect 92480 150078 92532 150084
rect 95528 149940 95556 150690
rect 97920 150210 97948 152186
rect 105820 151836 105872 151842
rect 105740 151786 105820 151814
rect 102324 151768 102376 151774
rect 102324 151710 102376 151716
rect 98920 151700 98972 151706
rect 98920 151642 98972 151648
rect 97908 150204 97960 150210
rect 97908 150146 97960 150152
rect 98932 149940 98960 151642
rect 102336 149940 102364 151710
rect 105740 149954 105768 151786
rect 105820 151778 105872 151784
rect 105740 149926 105846 149954
rect 82818 149696 82874 149705
rect 82818 149631 82874 149640
rect 109250 149382 109632 149410
rect 109604 148073 109632 149382
rect 109590 148064 109646 148073
rect 109590 147999 109646 148008
rect 109696 132494 109724 152322
rect 110340 151994 110368 155722
rect 110524 154766 110552 163200
rect 111352 157554 111380 163200
rect 111340 157548 111392 157554
rect 111340 157490 111392 157496
rect 112272 155786 112300 163200
rect 113100 159730 113128 163200
rect 113088 159724 113140 159730
rect 113088 159666 113140 159672
rect 112260 155780 112312 155786
rect 112260 155722 112312 155728
rect 110512 154760 110564 154766
rect 110512 154702 110564 154708
rect 113192 153202 113220 163254
rect 113836 163146 113864 163254
rect 113914 163200 113970 164400
rect 114742 163200 114798 164400
rect 115570 163200 115626 164400
rect 115952 163254 116348 163282
rect 113928 163146 113956 163200
rect 113836 163118 113956 163146
rect 114468 158772 114520 158778
rect 114468 158714 114520 158720
rect 114480 154630 114508 158714
rect 114756 157486 114784 163200
rect 114744 157480 114796 157486
rect 114744 157422 114796 157428
rect 115584 157185 115612 163200
rect 115570 157176 115626 157185
rect 115570 157111 115626 157120
rect 114468 154624 114520 154630
rect 114468 154566 114520 154572
rect 115952 154426 115980 163254
rect 116320 163146 116348 163254
rect 116398 163200 116454 164400
rect 117226 163200 117282 164400
rect 118146 163200 118202 164400
rect 118712 163254 118924 163282
rect 116412 163146 116440 163200
rect 116320 163118 116440 163146
rect 117240 160002 117268 163200
rect 117228 159996 117280 160002
rect 117228 159938 117280 159944
rect 118160 156126 118188 163200
rect 118148 156120 118200 156126
rect 118148 156062 118200 156068
rect 115940 154420 115992 154426
rect 115940 154362 115992 154368
rect 118712 153270 118740 163254
rect 118896 163146 118924 163254
rect 118974 163200 119030 164400
rect 119802 163200 119858 164400
rect 120092 163254 120580 163282
rect 118988 163146 119016 163200
rect 118896 163118 119016 163146
rect 119816 158778 119844 163200
rect 119804 158772 119856 158778
rect 119804 158714 119856 158720
rect 118884 158024 118936 158030
rect 118884 157966 118936 157972
rect 118700 153264 118752 153270
rect 118700 153206 118752 153212
rect 110972 153196 111024 153202
rect 110972 153138 111024 153144
rect 113180 153196 113232 153202
rect 113180 153138 113232 153144
rect 110512 152380 110564 152386
rect 110512 152322 110564 152328
rect 110340 151966 110460 151994
rect 110328 151904 110380 151910
rect 110328 151846 110380 151852
rect 110236 151836 110288 151842
rect 110236 151778 110288 151784
rect 110248 146418 110276 151778
rect 110340 150278 110368 151846
rect 110432 151842 110460 151966
rect 110524 151910 110552 152322
rect 110512 151904 110564 151910
rect 110512 151846 110564 151852
rect 110420 151836 110472 151842
rect 110984 151814 111012 153138
rect 110984 151786 111196 151814
rect 110420 151778 110472 151784
rect 110972 151632 111024 151638
rect 110972 151574 111024 151580
rect 110328 150272 110380 150278
rect 110328 150214 110380 150220
rect 110984 147937 111012 151574
rect 111062 150512 111118 150521
rect 111062 150447 111118 150456
rect 110970 147928 111026 147937
rect 110970 147863 111026 147872
rect 110326 146432 110382 146441
rect 110248 146390 110326 146418
rect 110326 146367 110382 146376
rect 109696 132466 110368 132494
rect 110340 106321 110368 132466
rect 110326 106312 110382 106321
rect 110326 106247 110382 106256
rect 111076 89690 111104 150447
rect 111168 148374 111196 151786
rect 116124 151768 116176 151774
rect 116124 151710 116176 151716
rect 116032 151700 116084 151706
rect 116032 151642 116084 151648
rect 113088 151564 113140 151570
rect 113088 151506 113140 151512
rect 112720 151292 112772 151298
rect 112720 151234 112772 151240
rect 112628 151224 112680 151230
rect 112628 151166 112680 151172
rect 112536 151156 112588 151162
rect 112536 151098 112588 151104
rect 111708 151088 111760 151094
rect 111708 151030 111760 151036
rect 111616 150952 111668 150958
rect 111616 150894 111668 150900
rect 111524 150884 111576 150890
rect 111524 150826 111576 150832
rect 111432 150816 111484 150822
rect 111432 150758 111484 150764
rect 111248 150680 111300 150686
rect 111248 150622 111300 150628
rect 111338 150648 111394 150657
rect 111156 148368 111208 148374
rect 111156 148310 111208 148316
rect 111260 148186 111288 150622
rect 111338 150583 111394 150592
rect 111168 148158 111288 148186
rect 111168 109002 111196 148158
rect 111352 148050 111380 150583
rect 111260 148022 111380 148050
rect 111156 108996 111208 109002
rect 111156 108938 111208 108944
rect 111260 92478 111288 148022
rect 111338 147928 111394 147937
rect 111338 147863 111394 147872
rect 111352 111790 111380 147863
rect 111444 113150 111472 150758
rect 111536 114510 111564 150826
rect 111628 117298 111656 150894
rect 111720 121446 111748 151030
rect 112444 151020 112496 151026
rect 112444 150962 112496 150968
rect 111708 121440 111760 121446
rect 111708 121382 111760 121388
rect 112456 118658 112484 150962
rect 112548 122806 112576 151098
rect 112640 124166 112668 151166
rect 112732 126954 112760 151234
rect 112996 150612 113048 150618
rect 112996 150554 113048 150560
rect 112904 150476 112956 150482
rect 112904 150418 112956 150424
rect 112812 150340 112864 150346
rect 112812 150282 112864 150288
rect 112824 132462 112852 150282
rect 112916 133890 112944 150418
rect 113008 137970 113036 150554
rect 113100 140758 113128 151506
rect 115296 150748 115348 150754
rect 115296 150690 115348 150696
rect 115204 150544 115256 150550
rect 115204 150486 115256 150492
rect 113822 144256 113878 144265
rect 113822 144191 113878 144200
rect 113088 140752 113140 140758
rect 113088 140694 113140 140700
rect 112996 137964 113048 137970
rect 112996 137906 113048 137912
rect 112904 133884 112956 133890
rect 112904 133826 112956 133832
rect 112812 132456 112864 132462
rect 112812 132398 112864 132404
rect 112720 126948 112772 126954
rect 112720 126890 112772 126896
rect 112628 124160 112680 124166
rect 112628 124102 112680 124108
rect 112536 122800 112588 122806
rect 112536 122742 112588 122748
rect 112444 118652 112496 118658
rect 112444 118594 112496 118600
rect 111616 117292 111668 117298
rect 111616 117234 111668 117240
rect 111524 114504 111576 114510
rect 111524 114446 111576 114452
rect 111432 113144 111484 113150
rect 111432 113086 111484 113092
rect 111340 111784 111392 111790
rect 111340 111726 111392 111732
rect 111248 92472 111300 92478
rect 111248 92414 111300 92420
rect 111064 89684 111116 89690
rect 111064 89626 111116 89632
rect 113836 88330 113864 144191
rect 115216 135561 115244 150486
rect 115308 141409 115336 150690
rect 116044 143313 116072 151642
rect 116136 145217 116164 151710
rect 116952 151496 117004 151502
rect 116952 151438 117004 151444
rect 116768 151428 116820 151434
rect 116768 151370 116820 151376
rect 116676 151360 116728 151366
rect 116676 151302 116728 151308
rect 116492 150068 116544 150074
rect 116492 150010 116544 150016
rect 116122 145208 116178 145217
rect 116122 145143 116178 145152
rect 116030 143304 116086 143313
rect 116030 143239 116086 143248
rect 115294 141400 115350 141409
rect 115294 141335 115350 141344
rect 116124 140752 116176 140758
rect 116124 140694 116176 140700
rect 116136 139505 116164 140694
rect 116122 139496 116178 139505
rect 116122 139431 116178 139440
rect 116124 137964 116176 137970
rect 116124 137906 116176 137912
rect 116136 137601 116164 137906
rect 116122 137592 116178 137601
rect 116122 137527 116178 137536
rect 115202 135552 115258 135561
rect 115202 135487 115258 135496
rect 116032 133884 116084 133890
rect 116032 133826 116084 133832
rect 116044 133657 116072 133826
rect 116030 133648 116086 133657
rect 116030 133583 116086 133592
rect 114190 132832 114246 132841
rect 114190 132767 114246 132776
rect 114204 132666 114232 132767
rect 114192 132660 114244 132666
rect 114192 132602 114244 132608
rect 115204 132660 115256 132666
rect 115204 132602 115256 132608
rect 113914 121408 113970 121417
rect 113914 121343 113970 121352
rect 113824 88324 113876 88330
rect 113824 88266 113876 88272
rect 113928 83978 113956 121343
rect 114006 110120 114062 110129
rect 114006 110055 114062 110064
rect 113916 83972 113968 83978
rect 113916 83914 113968 83920
rect 114020 82822 114048 110055
rect 114098 98696 114154 98705
rect 114098 98631 114154 98640
rect 114008 82816 114060 82822
rect 114008 82758 114060 82764
rect 114112 80034 114140 98631
rect 114190 87272 114246 87281
rect 114190 87207 114246 87216
rect 114100 80028 114152 80034
rect 114100 79970 114152 79976
rect 114204 78674 114232 87207
rect 115216 85649 115244 132602
rect 116124 132456 116176 132462
rect 116124 132398 116176 132404
rect 116136 131753 116164 132398
rect 116122 131744 116178 131753
rect 116122 131679 116178 131688
rect 116504 129849 116532 150010
rect 116582 149696 116638 149705
rect 116582 149631 116638 149640
rect 116490 129840 116546 129849
rect 116490 129775 116546 129784
rect 116124 126948 116176 126954
rect 116124 126890 116176 126896
rect 116136 126041 116164 126890
rect 116122 126032 116178 126041
rect 116122 125967 116178 125976
rect 116124 124160 116176 124166
rect 116122 124128 116124 124137
rect 116176 124128 116178 124137
rect 116122 124063 116178 124072
rect 115940 122800 115992 122806
rect 115940 122742 115992 122748
rect 115952 122233 115980 122742
rect 115938 122224 115994 122233
rect 115938 122159 115994 122168
rect 116124 121440 116176 121446
rect 116124 121382 116176 121388
rect 116136 120193 116164 121382
rect 116122 120184 116178 120193
rect 116122 120119 116178 120128
rect 116124 118652 116176 118658
rect 116124 118594 116176 118600
rect 116136 118289 116164 118594
rect 116122 118280 116178 118289
rect 116122 118215 116178 118224
rect 116124 117292 116176 117298
rect 116124 117234 116176 117240
rect 116136 116385 116164 117234
rect 116122 116376 116178 116385
rect 116122 116311 116178 116320
rect 116124 114504 116176 114510
rect 116122 114472 116124 114481
rect 116176 114472 116178 114481
rect 116122 114407 116178 114416
rect 115940 113144 115992 113150
rect 115940 113086 115992 113092
rect 115952 112577 115980 113086
rect 115938 112568 115994 112577
rect 115938 112503 115994 112512
rect 116124 111784 116176 111790
rect 116124 111726 116176 111732
rect 116136 110673 116164 111726
rect 116122 110664 116178 110673
rect 116122 110599 116178 110608
rect 116124 108996 116176 109002
rect 116124 108938 116176 108944
rect 116136 108769 116164 108938
rect 116122 108760 116178 108769
rect 116122 108695 116178 108704
rect 116596 93401 116624 149631
rect 116688 95305 116716 151302
rect 116780 97209 116808 151370
rect 116860 150204 116912 150210
rect 116860 150146 116912 150152
rect 116872 99113 116900 150146
rect 116964 102921 116992 151438
rect 117136 150272 117188 150278
rect 117136 150214 117188 150220
rect 117044 148368 117096 148374
rect 117044 148310 117096 148316
rect 116950 102912 117006 102921
rect 116950 102847 117006 102856
rect 117056 101017 117084 148310
rect 117148 104825 117176 150214
rect 117228 150136 117280 150142
rect 117228 150078 117280 150084
rect 117240 132546 117268 150078
rect 118896 149954 118924 157966
rect 119988 154624 120040 154630
rect 119988 154566 120040 154572
rect 120000 154426 120028 154566
rect 119896 154420 119948 154426
rect 119896 154362 119948 154368
rect 119988 154420 120040 154426
rect 119988 154362 120040 154368
rect 119908 153882 119936 154362
rect 119804 153876 119856 153882
rect 119804 153818 119856 153824
rect 119896 153876 119948 153882
rect 119896 153818 119948 153824
rect 119816 150226 119844 153818
rect 120092 152386 120120 163254
rect 120552 163146 120580 163254
rect 120630 163200 120686 164400
rect 121458 163200 121514 164400
rect 122286 163200 122342 164400
rect 123114 163200 123170 164400
rect 124034 163200 124090 164400
rect 124862 163200 124918 164400
rect 125690 163200 125746 164400
rect 126518 163200 126574 164400
rect 126992 163254 127296 163282
rect 120644 163146 120672 163200
rect 120552 163118 120672 163146
rect 120448 156664 120500 156670
rect 120448 156606 120500 156612
rect 120080 152380 120132 152386
rect 120080 152322 120132 152328
rect 120460 150226 120488 156606
rect 121472 156058 121500 163200
rect 121920 158976 121972 158982
rect 121920 158918 121972 158924
rect 121460 156052 121512 156058
rect 121460 155994 121512 156000
rect 121932 153785 121960 158918
rect 122012 155304 122064 155310
rect 122012 155246 122064 155252
rect 121734 153776 121790 153785
rect 121734 153711 121790 153720
rect 121918 153776 121974 153785
rect 121918 153711 121974 153720
rect 121092 152516 121144 152522
rect 121092 152458 121144 152464
rect 121104 150226 121132 152458
rect 121748 150226 121776 153711
rect 122024 151814 122052 155246
rect 122300 154970 122328 163200
rect 123128 159390 123156 163200
rect 122840 159384 122892 159390
rect 122840 159326 122892 159332
rect 123116 159384 123168 159390
rect 123116 159326 123168 159332
rect 122288 154964 122340 154970
rect 122288 154906 122340 154912
rect 122024 151786 122420 151814
rect 122392 150226 122420 151786
rect 119816 150198 119890 150226
rect 120460 150198 120534 150226
rect 121104 150198 121178 150226
rect 121748 150198 121822 150226
rect 122392 150198 122466 150226
rect 122852 150210 122880 159326
rect 124048 158982 124076 163200
rect 124036 158976 124088 158982
rect 124036 158918 124088 158924
rect 124876 156670 124904 163200
rect 125704 161474 125732 163200
rect 125704 161446 125824 161474
rect 125508 158908 125560 158914
rect 125508 158850 125560 158856
rect 124864 156664 124916 156670
rect 124864 156606 124916 156612
rect 124680 155440 124732 155446
rect 124680 155382 124732 155388
rect 123024 155236 123076 155242
rect 123024 155178 123076 155184
rect 123036 150226 123064 155178
rect 124312 153944 124364 153950
rect 124312 153886 124364 153892
rect 124324 150226 124352 153886
rect 124692 151814 124720 155382
rect 125520 153950 125548 158850
rect 125692 155372 125744 155378
rect 125692 155314 125744 155320
rect 125508 153944 125560 153950
rect 125508 153886 125560 153892
rect 124692 151786 124996 151814
rect 124968 150226 124996 151786
rect 125704 150226 125732 155314
rect 125796 154834 125824 161446
rect 126532 160138 126560 163200
rect 126520 160132 126572 160138
rect 126520 160074 126572 160080
rect 126428 159724 126480 159730
rect 126428 159666 126480 159672
rect 126440 159526 126468 159666
rect 126428 159520 126480 159526
rect 126428 159462 126480 159468
rect 126244 159452 126296 159458
rect 126244 159394 126296 159400
rect 126796 159452 126848 159458
rect 126796 159394 126848 159400
rect 126256 158914 126284 159394
rect 126244 158908 126296 158914
rect 126244 158850 126296 158856
rect 125784 154828 125836 154834
rect 125784 154770 125836 154776
rect 126808 152425 126836 159394
rect 126888 154012 126940 154018
rect 126888 153954 126940 153960
rect 126242 152416 126298 152425
rect 126242 152351 126298 152360
rect 126794 152416 126850 152425
rect 126794 152351 126850 152360
rect 118896 149926 119324 149954
rect 119862 149940 119890 150198
rect 120506 149940 120534 150198
rect 121150 149940 121178 150198
rect 121794 149940 121822 150198
rect 122438 149940 122466 150198
rect 122840 150204 122892 150210
rect 123036 150198 123110 150226
rect 122840 150146 122892 150152
rect 123082 149940 123110 150198
rect 123714 150204 123766 150210
rect 124324 150198 124398 150226
rect 124968 150198 125042 150226
rect 123714 150146 123766 150152
rect 123726 149940 123754 150146
rect 124370 149940 124398 150198
rect 125014 149940 125042 150198
rect 125658 150198 125732 150226
rect 126256 150226 126284 152351
rect 126900 150226 126928 153954
rect 126992 152522 127020 163254
rect 127268 163146 127296 163254
rect 127346 163200 127402 164400
rect 128174 163200 128230 164400
rect 129002 163200 129058 164400
rect 129922 163200 129978 164400
rect 130750 163200 130806 164400
rect 131578 163200 131634 164400
rect 132406 163200 132462 164400
rect 133234 163200 133290 164400
rect 134062 163200 134118 164400
rect 134890 163200 134946 164400
rect 135810 163200 135866 164400
rect 136638 163200 136694 164400
rect 137466 163200 137522 164400
rect 138294 163200 138350 164400
rect 139122 163200 139178 164400
rect 139950 163200 140006 164400
rect 140778 163200 140834 164400
rect 141698 163200 141754 164400
rect 142526 163200 142582 164400
rect 143354 163200 143410 164400
rect 144182 163200 144238 164400
rect 145010 163200 145066 164400
rect 145838 163200 145894 164400
rect 146666 163200 146722 164400
rect 147586 163200 147642 164400
rect 148414 163200 148470 164400
rect 149242 163200 149298 164400
rect 150070 163200 150126 164400
rect 150898 163200 150954 164400
rect 151726 163200 151782 164400
rect 151832 163254 152504 163282
rect 127360 163146 127388 163200
rect 127268 163118 127388 163146
rect 127808 159520 127860 159526
rect 127808 159462 127860 159468
rect 127532 156732 127584 156738
rect 127532 156674 127584 156680
rect 126980 152516 127032 152522
rect 126980 152458 127032 152464
rect 127544 150226 127572 156674
rect 127820 153950 127848 159462
rect 128188 156738 128216 163200
rect 128176 156732 128228 156738
rect 128176 156674 128228 156680
rect 129016 155242 129044 163200
rect 129936 159594 129964 163200
rect 129924 159588 129976 159594
rect 129924 159530 129976 159536
rect 129924 159384 129976 159390
rect 129924 159326 129976 159332
rect 129740 158908 129792 158914
rect 129740 158850 129792 158856
rect 129004 155236 129056 155242
rect 129004 155178 129056 155184
rect 129464 154080 129516 154086
rect 129464 154022 129516 154028
rect 127716 153944 127768 153950
rect 127716 153886 127768 153892
rect 127808 153944 127860 153950
rect 127808 153886 127860 153892
rect 127624 153876 127676 153882
rect 127624 153818 127676 153824
rect 127636 153270 127664 153818
rect 127728 153270 127756 153886
rect 127624 153264 127676 153270
rect 127624 153206 127676 153212
rect 127716 153264 127768 153270
rect 127716 153206 127768 153212
rect 128818 152552 128874 152561
rect 128818 152487 128874 152496
rect 128176 151836 128228 151842
rect 128176 151778 128228 151784
rect 128188 150226 128216 151778
rect 128832 150226 128860 152487
rect 129476 150226 129504 154022
rect 129752 151842 129780 158850
rect 129936 158846 129964 159326
rect 130764 158914 130792 163200
rect 131212 159792 131264 159798
rect 131212 159734 131264 159740
rect 131592 159746 131620 163200
rect 131224 159526 131252 159734
rect 131592 159718 131804 159746
rect 131672 159656 131724 159662
rect 131316 159604 131672 159610
rect 131316 159598 131724 159604
rect 131316 159582 131712 159598
rect 131120 159520 131172 159526
rect 131120 159462 131172 159468
rect 131212 159520 131264 159526
rect 131212 159462 131264 159468
rect 131026 159352 131082 159361
rect 131132 159338 131160 159462
rect 131316 159338 131344 159582
rect 131132 159310 131344 159338
rect 131026 159287 131082 159296
rect 130752 158908 130804 158914
rect 130752 158850 130804 158856
rect 129924 158840 129976 158846
rect 129924 158782 129976 158788
rect 130108 156800 130160 156806
rect 130108 156742 130160 156748
rect 129740 151836 129792 151842
rect 129740 151778 129792 151784
rect 130120 150226 130148 156742
rect 130752 152244 130804 152250
rect 130752 152186 130804 152192
rect 130764 150226 130792 152186
rect 131040 151814 131068 159287
rect 131776 158030 131804 159718
rect 131764 158024 131816 158030
rect 131764 157966 131816 157972
rect 132420 153950 132448 163200
rect 133248 158846 133276 163200
rect 133602 159488 133658 159497
rect 133602 159423 133658 159432
rect 133236 158840 133288 158846
rect 133236 158782 133288 158788
rect 132500 156868 132552 156874
rect 132500 156810 132552 156816
rect 132408 153944 132460 153950
rect 132038 153912 132094 153921
rect 132408 153886 132460 153892
rect 132038 153847 132094 153856
rect 131040 151786 131436 151814
rect 131408 150226 131436 151786
rect 132052 150226 132080 153847
rect 132512 151814 132540 156810
rect 133052 154692 133104 154698
rect 133052 154634 133104 154640
rect 133064 151814 133092 154634
rect 133616 153105 133644 159423
rect 133602 153096 133658 153105
rect 133602 153031 133658 153040
rect 133972 152584 134024 152590
rect 133972 152526 134024 152532
rect 132512 151786 132724 151814
rect 133064 151786 133368 151814
rect 132696 150226 132724 151786
rect 133340 150226 133368 151786
rect 133984 150226 134012 152526
rect 134076 152250 134104 163200
rect 134156 160132 134208 160138
rect 134156 160074 134208 160080
rect 134168 159730 134196 160074
rect 134156 159724 134208 159730
rect 134156 159666 134208 159672
rect 134904 156874 134932 163200
rect 135824 156942 135852 163200
rect 136652 159662 136680 163200
rect 136548 159656 136600 159662
rect 136548 159598 136600 159604
rect 136640 159656 136692 159662
rect 136640 159598 136692 159604
rect 136560 159474 136588 159598
rect 136560 159446 136680 159474
rect 135260 156936 135312 156942
rect 135260 156878 135312 156884
rect 135812 156936 135864 156942
rect 135812 156878 135864 156884
rect 134892 156868 134944 156874
rect 134892 156810 134944 156816
rect 134614 154048 134670 154057
rect 134614 153983 134670 153992
rect 134064 152244 134116 152250
rect 134064 152186 134116 152192
rect 134628 150226 134656 153983
rect 135272 150226 135300 156878
rect 136546 153096 136602 153105
rect 136546 153031 136602 153040
rect 135904 152652 135956 152658
rect 135904 152594 135956 152600
rect 135916 150226 135944 152594
rect 136560 150226 136588 153031
rect 136652 152590 136680 159446
rect 137480 159390 137508 163200
rect 138018 159624 138074 159633
rect 138018 159559 138074 159568
rect 137100 159384 137152 159390
rect 137100 159326 137152 159332
rect 137468 159384 137520 159390
rect 137468 159326 137520 159332
rect 137112 154630 137140 159326
rect 138032 157334 138060 159559
rect 138032 157306 138152 157334
rect 137376 157004 137428 157010
rect 137376 156946 137428 156952
rect 137100 154624 137152 154630
rect 137100 154566 137152 154572
rect 136916 154216 136968 154222
rect 136916 154158 136968 154164
rect 136640 152584 136692 152590
rect 136640 152526 136692 152532
rect 126256 150198 126330 150226
rect 126900 150198 126974 150226
rect 127544 150198 127618 150226
rect 128188 150198 128262 150226
rect 128832 150198 128906 150226
rect 129476 150198 129550 150226
rect 130120 150198 130194 150226
rect 130764 150198 130838 150226
rect 131408 150198 131482 150226
rect 132052 150198 132126 150226
rect 132696 150198 132770 150226
rect 133340 150198 133414 150226
rect 133984 150198 134058 150226
rect 134628 150198 134702 150226
rect 135272 150198 135346 150226
rect 135916 150198 135990 150226
rect 136560 150198 136634 150226
rect 136928 150210 136956 154158
rect 137008 154148 137060 154154
rect 137008 154090 137060 154096
rect 137020 151814 137048 154090
rect 137388 151814 137416 156946
rect 138124 152862 138152 157306
rect 138308 157010 138336 163200
rect 138296 157004 138348 157010
rect 138296 156946 138348 156952
rect 139136 156806 139164 163200
rect 139964 159662 139992 163200
rect 139400 159656 139452 159662
rect 139400 159598 139452 159604
rect 139952 159656 140004 159662
rect 139952 159598 140004 159604
rect 139412 157334 139440 159598
rect 139412 157306 139900 157334
rect 139124 156800 139176 156806
rect 139124 156742 139176 156748
rect 139308 154760 139360 154766
rect 139308 154702 139360 154708
rect 138204 154624 138256 154630
rect 138256 154572 138428 154574
rect 138204 154566 138428 154572
rect 138216 154546 138428 154566
rect 138400 154086 138428 154546
rect 138388 154080 138440 154086
rect 138388 154022 138440 154028
rect 138020 152856 138072 152862
rect 138020 152798 138072 152804
rect 138112 152856 138164 152862
rect 138112 152798 138164 152804
rect 138032 152674 138060 152798
rect 139124 152788 139176 152794
rect 139124 152730 139176 152736
rect 138032 152646 138152 152674
rect 138124 152590 138152 152646
rect 138112 152584 138164 152590
rect 138112 152526 138164 152532
rect 138480 151904 138532 151910
rect 138480 151846 138532 151852
rect 137020 151786 137232 151814
rect 137388 151786 137876 151814
rect 137204 150226 137232 151786
rect 137848 150226 137876 151786
rect 125658 149940 125686 150198
rect 126302 149940 126330 150198
rect 126946 149940 126974 150198
rect 127590 149940 127618 150198
rect 128234 149940 128262 150198
rect 128878 149940 128906 150198
rect 129522 149940 129550 150198
rect 130166 149940 130194 150198
rect 130810 149940 130838 150198
rect 131454 149940 131482 150198
rect 132098 149940 132126 150198
rect 132742 149940 132770 150198
rect 133386 149940 133414 150198
rect 134030 149940 134058 150198
rect 134674 149940 134702 150198
rect 135318 149940 135346 150198
rect 135962 149940 135990 150198
rect 136606 149940 136634 150198
rect 136916 150204 136968 150210
rect 137204 150198 137278 150226
rect 137848 150198 137922 150226
rect 136916 150146 136968 150152
rect 137250 149940 137278 150198
rect 137894 149940 137922 150198
rect 138492 150090 138520 151846
rect 139136 150090 139164 152730
rect 139320 151910 139348 154702
rect 139872 153950 139900 157306
rect 140410 156632 140466 156641
rect 140410 156567 140466 156576
rect 139860 153944 139912 153950
rect 139860 153886 139912 153892
rect 139308 151904 139360 151910
rect 139308 151846 139360 151852
rect 139814 150204 139866 150210
rect 139814 150146 139866 150152
rect 138492 150062 138566 150090
rect 139136 150062 139210 150090
rect 138538 149940 138566 150062
rect 139182 149940 139210 150062
rect 139826 149940 139854 150146
rect 140424 150090 140452 156567
rect 140792 152794 140820 163200
rect 141712 157418 141740 163200
rect 141700 157412 141752 157418
rect 141700 157354 141752 157360
rect 142540 155310 142568 163200
rect 143368 159798 143396 163200
rect 143264 159792 143316 159798
rect 143264 159734 143316 159740
rect 143356 159792 143408 159798
rect 143356 159734 143408 159740
rect 143078 156768 143134 156777
rect 143078 156703 143134 156712
rect 142528 155304 142580 155310
rect 142528 155246 142580 155252
rect 142448 154550 142752 154578
rect 142342 154184 142398 154193
rect 142448 154154 142476 154550
rect 142528 154488 142580 154494
rect 142528 154430 142580 154436
rect 142342 154119 142398 154128
rect 142436 154148 142488 154154
rect 141700 152856 141752 152862
rect 141700 152798 141752 152804
rect 140780 152788 140832 152794
rect 140780 152730 140832 152736
rect 141056 152720 141108 152726
rect 141056 152662 141108 152668
rect 141068 150090 141096 152662
rect 141712 150090 141740 152798
rect 142356 150090 142384 154119
rect 142436 154090 142488 154096
rect 142540 153950 142568 154430
rect 142724 154358 142752 154550
rect 142804 154488 142856 154494
rect 142804 154430 142856 154436
rect 142620 154352 142672 154358
rect 142620 154294 142672 154300
rect 142712 154352 142764 154358
rect 142712 154294 142764 154300
rect 142632 154193 142660 154294
rect 142816 154222 142844 154430
rect 142804 154216 142856 154222
rect 142618 154184 142674 154193
rect 142804 154158 142856 154164
rect 142618 154119 142674 154128
rect 142436 153944 142488 153950
rect 142434 153912 142436 153921
rect 142528 153944 142580 153950
rect 142488 153912 142490 153921
rect 142988 153944 143040 153950
rect 142528 153886 142580 153892
rect 142986 153912 142988 153921
rect 143040 153912 143042 153921
rect 142434 153847 142490 153856
rect 142804 153876 142856 153882
rect 142986 153847 143042 153856
rect 142804 153818 142856 153824
rect 142710 153368 142766 153377
rect 142816 153338 142844 153818
rect 142710 153303 142712 153312
rect 142764 153303 142766 153312
rect 142804 153332 142856 153338
rect 142712 153274 142764 153280
rect 142804 153274 142856 153280
rect 142804 152720 142856 152726
rect 142804 152662 142856 152668
rect 142816 152046 142844 152662
rect 142804 152040 142856 152046
rect 142804 151982 142856 151988
rect 143092 150090 143120 156703
rect 143172 154284 143224 154290
rect 143172 154226 143224 154232
rect 143184 154086 143212 154226
rect 143172 154080 143224 154086
rect 143172 154022 143224 154028
rect 143276 152046 143304 159734
rect 144196 159526 144224 163200
rect 144092 159520 144144 159526
rect 144092 159462 144144 159468
rect 144184 159520 144236 159526
rect 144184 159462 144236 159468
rect 144104 159338 144132 159462
rect 144104 159310 144408 159338
rect 143446 154184 143502 154193
rect 143446 154119 143448 154128
rect 143500 154119 143502 154128
rect 143448 154090 143500 154096
rect 143356 154080 143408 154086
rect 143356 154022 143408 154028
rect 143368 153377 143396 154022
rect 143354 153368 143410 153377
rect 143354 153303 143410 153312
rect 144380 152794 144408 159310
rect 144918 157992 144974 158001
rect 144918 157927 144974 157936
rect 144276 152788 144328 152794
rect 144276 152730 144328 152736
rect 144368 152788 144420 152794
rect 144368 152730 144420 152736
rect 144288 152674 144316 152730
rect 144288 152646 144408 152674
rect 144380 152590 144408 152646
rect 144276 152584 144328 152590
rect 144276 152526 144328 152532
rect 144368 152584 144420 152590
rect 144368 152526 144420 152532
rect 143630 152416 143686 152425
rect 143630 152351 143686 152360
rect 143264 152040 143316 152046
rect 143264 151982 143316 151988
rect 140424 150062 140498 150090
rect 141068 150062 141142 150090
rect 141712 150062 141786 150090
rect 142356 150062 142430 150090
rect 140470 149940 140498 150062
rect 141114 149940 141142 150062
rect 141758 149940 141786 150062
rect 142402 149940 142430 150062
rect 143046 150062 143120 150090
rect 143644 150090 143672 152351
rect 144288 150090 144316 152526
rect 144932 150226 144960 157927
rect 145024 155990 145052 163200
rect 145012 155984 145064 155990
rect 145012 155926 145064 155932
rect 145852 155378 145880 163200
rect 146484 160064 146536 160070
rect 146484 160006 146536 160012
rect 146392 158092 146444 158098
rect 146392 158034 146444 158040
rect 146208 157072 146260 157078
rect 146208 157014 146260 157020
rect 145840 155372 145892 155378
rect 145840 155314 145892 155320
rect 145564 154148 145616 154154
rect 145564 154090 145616 154096
rect 144932 150198 145006 150226
rect 143644 150062 143718 150090
rect 144288 150062 144362 150090
rect 143046 149940 143074 150062
rect 143690 149940 143718 150062
rect 144334 149940 144362 150062
rect 144978 149940 145006 150198
rect 145576 150090 145604 154090
rect 146220 150090 146248 157014
rect 146404 150210 146432 158034
rect 146496 152862 146524 160006
rect 146680 158778 146708 163200
rect 146944 160064 146996 160070
rect 146944 160006 146996 160012
rect 146956 159594 146984 160006
rect 146944 159588 146996 159594
rect 146944 159530 146996 159536
rect 147600 159458 147628 163200
rect 147496 159452 147548 159458
rect 147496 159394 147548 159400
rect 147588 159452 147640 159458
rect 147588 159394 147640 159400
rect 147508 159338 147536 159394
rect 147508 159310 147812 159338
rect 146576 158772 146628 158778
rect 146576 158714 146628 158720
rect 146668 158772 146720 158778
rect 146668 158714 146720 158720
rect 146588 158658 146616 158714
rect 146588 158630 147168 158658
rect 147140 154154 147168 158630
rect 147680 157140 147732 157146
rect 147680 157082 147732 157088
rect 147588 154216 147640 154222
rect 147586 154184 147588 154193
rect 147640 154184 147642 154193
rect 147128 154148 147180 154154
rect 147586 154119 147642 154128
rect 147128 154090 147180 154096
rect 146484 152856 146536 152862
rect 146484 152798 146536 152804
rect 146944 152040 146996 152046
rect 146944 151982 146996 151988
rect 146956 151842 146984 151982
rect 146852 151836 146904 151842
rect 146852 151778 146904 151784
rect 146944 151836 146996 151842
rect 146944 151778 146996 151784
rect 146392 150204 146444 150210
rect 146392 150146 146444 150152
rect 146864 150090 146892 151778
rect 147692 150210 147720 157082
rect 147784 154222 147812 159310
rect 148428 158098 148456 163200
rect 148416 158092 148468 158098
rect 148416 158034 148468 158040
rect 149256 155446 149284 163200
rect 149520 159452 149572 159458
rect 149520 159394 149572 159400
rect 149244 155440 149296 155446
rect 149244 155382 149296 155388
rect 147772 154216 147824 154222
rect 147772 154158 147824 154164
rect 148138 154184 148194 154193
rect 148138 154119 148194 154128
rect 148152 150226 148180 154119
rect 149532 152726 149560 159394
rect 149610 158264 149666 158273
rect 149610 158199 149666 158208
rect 149428 152720 149480 152726
rect 149428 152662 149480 152668
rect 149520 152720 149572 152726
rect 149520 152662 149572 152668
rect 149440 150226 149468 152662
rect 149624 151814 149652 158199
rect 150084 157146 150112 163200
rect 150912 159458 150940 163200
rect 150900 159452 150952 159458
rect 150900 159394 150952 159400
rect 151268 157208 151320 157214
rect 151268 157150 151320 157156
rect 150072 157140 150124 157146
rect 150072 157082 150124 157088
rect 150624 154080 150676 154086
rect 150624 154022 150676 154028
rect 149624 151786 150020 151814
rect 149992 150226 150020 151786
rect 150636 150226 150664 154022
rect 151280 150226 151308 157150
rect 151740 157078 151768 163200
rect 151728 157072 151780 157078
rect 151728 157014 151780 157020
rect 151832 154086 151860 163254
rect 152476 163146 152504 163254
rect 152554 163200 152610 164400
rect 153474 163200 153530 164400
rect 153580 163254 154252 163282
rect 152568 163146 152596 163200
rect 152476 163118 152596 163146
rect 153488 159866 153516 163200
rect 153384 159860 153436 159866
rect 153384 159802 153436 159808
rect 153476 159860 153528 159866
rect 153476 159802 153528 159808
rect 153396 159594 153424 159802
rect 153384 159588 153436 159594
rect 153384 159530 153436 159536
rect 152554 158128 152610 158137
rect 152554 158063 152610 158072
rect 151820 154080 151872 154086
rect 151820 154022 151872 154028
rect 151912 152652 151964 152658
rect 151912 152594 151964 152600
rect 151924 150226 151952 152594
rect 152568 150226 152596 158063
rect 153292 153876 153344 153882
rect 153292 153818 153344 153824
rect 153304 150226 153332 153818
rect 153580 152658 153608 163254
rect 154224 163146 154252 163254
rect 154302 163200 154358 164400
rect 155130 163200 155186 164400
rect 155958 163200 156014 164400
rect 156786 163200 156842 164400
rect 157614 163200 157670 164400
rect 158442 163200 158498 164400
rect 159362 163200 159418 164400
rect 160190 163200 160246 164400
rect 161018 163200 161074 164400
rect 161846 163200 161902 164400
rect 162674 163200 162730 164400
rect 163502 163200 163558 164400
rect 164330 163200 164386 164400
rect 165250 163200 165306 164400
rect 165632 163254 166028 163282
rect 154316 163146 154344 163200
rect 154224 163118 154344 163146
rect 154488 160064 154540 160070
rect 154488 160006 154540 160012
rect 153752 157276 153804 157282
rect 153752 157218 153804 157224
rect 153568 152652 153620 152658
rect 153568 152594 153620 152600
rect 153764 151814 153792 157218
rect 154500 154630 154528 160006
rect 155144 158166 155172 163200
rect 155040 158160 155092 158166
rect 155040 158102 155092 158108
rect 155132 158160 155184 158166
rect 155132 158102 155184 158108
rect 155052 157978 155080 158102
rect 155052 157950 155172 157978
rect 154488 154624 154540 154630
rect 154488 154566 154540 154572
rect 155040 154556 155092 154562
rect 155040 154498 155092 154504
rect 155052 153882 155080 154498
rect 155040 153876 155092 153882
rect 155040 153818 155092 153824
rect 154488 151972 154540 151978
rect 154488 151914 154540 151920
rect 153764 151786 153884 151814
rect 147542 150204 147594 150210
rect 147542 150146 147594 150152
rect 147680 150204 147732 150210
rect 148152 150198 148226 150226
rect 147680 150146 147732 150152
rect 145576 150062 145650 150090
rect 146220 150062 146294 150090
rect 146864 150062 146938 150090
rect 145622 149940 145650 150062
rect 146266 149940 146294 150062
rect 146910 149940 146938 150062
rect 147554 149940 147582 150146
rect 148198 149940 148226 150198
rect 148830 150204 148882 150210
rect 149440 150198 149514 150226
rect 149992 150198 150066 150226
rect 150636 150198 150710 150226
rect 151280 150198 151354 150226
rect 151924 150198 151998 150226
rect 152568 150198 152642 150226
rect 148830 150146 148882 150152
rect 148842 149940 148870 150146
rect 149486 149940 149514 150198
rect 150038 149940 150066 150198
rect 150682 149940 150710 150198
rect 151326 149940 151354 150198
rect 151970 149940 151998 150198
rect 152614 149940 152642 150198
rect 153258 150198 153332 150226
rect 153856 150226 153884 151786
rect 154500 150226 154528 151914
rect 155144 150226 155172 157950
rect 155972 154766 156000 163200
rect 156800 160070 156828 163200
rect 156788 160064 156840 160070
rect 156788 160006 156840 160012
rect 156512 159724 156564 159730
rect 156512 159666 156564 159672
rect 156420 157344 156472 157350
rect 156420 157286 156472 157292
rect 155960 154760 156012 154766
rect 155960 154702 156012 154708
rect 155868 154080 155920 154086
rect 155868 154022 155920 154028
rect 155880 153814 155908 154022
rect 155776 153808 155828 153814
rect 155776 153750 155828 153756
rect 155868 153808 155920 153814
rect 155868 153750 155920 153756
rect 155788 150226 155816 153750
rect 156432 150226 156460 157286
rect 156524 157214 156552 159666
rect 157628 159594 157656 163200
rect 156788 159588 156840 159594
rect 156788 159530 156840 159536
rect 157616 159588 157668 159594
rect 157616 159530 157668 159536
rect 156512 157208 156564 157214
rect 156512 157150 156564 157156
rect 156696 154624 156748 154630
rect 156696 154566 156748 154572
rect 156604 154556 156656 154562
rect 156604 154498 156656 154504
rect 156616 154222 156644 154498
rect 156604 154216 156656 154222
rect 156604 154158 156656 154164
rect 156512 154148 156564 154154
rect 156512 154090 156564 154096
rect 156524 153678 156552 154090
rect 156708 154086 156736 154566
rect 156604 154080 156656 154086
rect 156604 154022 156656 154028
rect 156696 154080 156748 154086
rect 156696 154022 156748 154028
rect 156616 153678 156644 154022
rect 156512 153672 156564 153678
rect 156512 153614 156564 153620
rect 156604 153672 156656 153678
rect 156604 153614 156656 153620
rect 156800 152046 156828 159530
rect 158456 158234 158484 163200
rect 158720 158840 158772 158846
rect 158720 158782 158772 158788
rect 157708 158228 157760 158234
rect 157708 158170 157760 158176
rect 158444 158228 158496 158234
rect 158444 158170 158496 158176
rect 156788 152040 156840 152046
rect 156788 151982 156840 151988
rect 157064 151836 157116 151842
rect 157064 151778 157116 151784
rect 157076 150226 157104 151778
rect 157720 150226 157748 158170
rect 158732 157350 158760 158782
rect 158720 157344 158772 157350
rect 158720 157286 158772 157292
rect 159088 157208 159140 157214
rect 159088 157150 159140 157156
rect 159100 156602 159128 157150
rect 158996 156596 159048 156602
rect 158996 156538 159048 156544
rect 159088 156596 159140 156602
rect 159088 156538 159140 156544
rect 158536 154080 158588 154086
rect 158536 154022 158588 154028
rect 158352 153876 158404 153882
rect 158352 153818 158404 153824
rect 158364 150226 158392 153818
rect 158548 153814 158576 154022
rect 158536 153808 158588 153814
rect 158536 153750 158588 153756
rect 159008 150226 159036 156538
rect 159376 154698 159404 163200
rect 160100 159792 160152 159798
rect 160100 159734 160152 159740
rect 160112 157214 160140 159734
rect 160100 157208 160152 157214
rect 160100 157150 160152 157156
rect 159364 154692 159416 154698
rect 159364 154634 159416 154640
rect 160204 154086 160232 163200
rect 161032 159662 161060 163200
rect 161020 159656 161072 159662
rect 161020 159598 161072 159604
rect 161860 158302 161888 163200
rect 162492 159928 162544 159934
rect 162492 159870 162544 159876
rect 160284 158296 160336 158302
rect 160284 158238 160336 158244
rect 161848 158296 161900 158302
rect 161848 158238 161900 158244
rect 160192 154080 160244 154086
rect 160192 154022 160244 154028
rect 159640 152448 159692 152454
rect 159640 152390 159692 152396
rect 159652 150226 159680 152390
rect 160296 150226 160324 158238
rect 161570 156904 161626 156913
rect 161570 156839 161626 156848
rect 160926 154320 160982 154329
rect 160926 154255 160982 154264
rect 160940 150226 160968 154255
rect 161584 150226 161612 156839
rect 162216 152788 162268 152794
rect 162216 152730 162268 152736
rect 162228 150226 162256 152730
rect 162504 151978 162532 159870
rect 162688 154630 162716 163200
rect 162872 159186 163084 159202
rect 162872 159180 163096 159186
rect 162872 159174 163044 159180
rect 162872 159118 162900 159174
rect 163044 159122 163096 159128
rect 162860 159112 162912 159118
rect 162860 159054 162912 159060
rect 163516 158846 163544 163200
rect 164344 161474 164372 163200
rect 164344 161446 164464 161474
rect 163780 159724 163832 159730
rect 163780 159666 163832 159672
rect 163504 158840 163556 158846
rect 163504 158782 163556 158788
rect 162858 158400 162914 158409
rect 162858 158335 162914 158344
rect 162676 154624 162728 154630
rect 162676 154566 162728 154572
rect 162492 151972 162544 151978
rect 162492 151914 162544 151920
rect 162872 150226 162900 158335
rect 163792 157282 163820 159666
rect 164332 158364 164384 158370
rect 164332 158306 164384 158312
rect 163780 157276 163832 157282
rect 163780 157218 163832 157224
rect 164148 156528 164200 156534
rect 164148 156470 164200 156476
rect 163504 154148 163556 154154
rect 163504 154090 163556 154096
rect 163516 150226 163544 154090
rect 164160 150226 164188 156470
rect 153856 150198 153930 150226
rect 154500 150198 154574 150226
rect 155144 150198 155218 150226
rect 155788 150198 155862 150226
rect 156432 150198 156506 150226
rect 157076 150198 157150 150226
rect 157720 150198 157794 150226
rect 158364 150198 158438 150226
rect 159008 150198 159082 150226
rect 159652 150198 159726 150226
rect 160296 150198 160370 150226
rect 160940 150198 161014 150226
rect 161584 150198 161658 150226
rect 162228 150198 162302 150226
rect 162872 150198 162946 150226
rect 163516 150198 163590 150226
rect 164160 150198 164234 150226
rect 164344 150210 164372 158306
rect 164436 152794 164464 161446
rect 165264 158370 165292 163200
rect 165252 158364 165304 158370
rect 165252 158306 165304 158312
rect 165632 154154 165660 163254
rect 166000 163146 166028 163254
rect 166078 163200 166134 164400
rect 166906 163200 166962 164400
rect 167734 163200 167790 164400
rect 168562 163200 168618 164400
rect 169390 163200 169446 164400
rect 170218 163200 170274 164400
rect 171138 163200 171194 164400
rect 171966 163200 172022 164400
rect 172532 163254 172744 163282
rect 166092 163146 166120 163200
rect 166000 163118 166120 163146
rect 166920 159934 166948 163200
rect 166908 159928 166960 159934
rect 166908 159870 166960 159876
rect 167748 159730 167776 163200
rect 167736 159724 167788 159730
rect 167736 159666 167788 159672
rect 167000 159316 167052 159322
rect 167000 159258 167052 159264
rect 166448 157276 166500 157282
rect 166448 157218 166500 157224
rect 166172 157208 166224 157214
rect 166172 157150 166224 157156
rect 166264 157208 166316 157214
rect 166264 157150 166316 157156
rect 166184 156534 166212 157150
rect 166172 156528 166224 156534
rect 166172 156470 166224 156476
rect 166276 156466 166304 157150
rect 166460 156534 166488 157218
rect 166448 156528 166500 156534
rect 166448 156470 166500 156476
rect 166264 156460 166316 156466
rect 166264 156402 166316 156408
rect 166722 155408 166778 155417
rect 166722 155343 166778 155352
rect 165620 154148 165672 154154
rect 165620 154090 165672 154096
rect 166080 153740 166132 153746
rect 166080 153682 166132 153688
rect 164424 152788 164476 152794
rect 164424 152730 164476 152736
rect 164792 152108 164844 152114
rect 164792 152050 164844 152056
rect 164804 150226 164832 152050
rect 166092 150226 166120 153682
rect 166736 150226 166764 155343
rect 167012 152114 167040 159258
rect 168576 158438 168604 163200
rect 167552 158432 167604 158438
rect 167552 158374 167604 158380
rect 168564 158432 168616 158438
rect 168564 158374 168616 158380
rect 167368 152856 167420 152862
rect 167368 152798 167420 152804
rect 167000 152108 167052 152114
rect 167000 152050 167052 152056
rect 167380 150226 167408 152798
rect 167564 151814 167592 158374
rect 168470 155544 168526 155553
rect 169404 155514 169432 163200
rect 170232 159322 170260 163200
rect 171152 159798 171180 163200
rect 171140 159792 171192 159798
rect 171140 159734 171192 159740
rect 170220 159316 170272 159322
rect 170220 159258 170272 159264
rect 169760 159112 169812 159118
rect 169760 159054 169812 159060
rect 169668 158432 169720 158438
rect 169666 158400 169668 158409
rect 169720 158400 169722 158409
rect 169666 158335 169722 158344
rect 168470 155479 168526 155488
rect 168656 155508 168708 155514
rect 167564 151786 168052 151814
rect 168024 150226 168052 151786
rect 153258 149940 153286 150198
rect 153902 149940 153930 150198
rect 154546 149940 154574 150198
rect 155190 149940 155218 150198
rect 155834 149940 155862 150198
rect 156478 149940 156506 150198
rect 157122 149940 157150 150198
rect 157766 149940 157794 150198
rect 158410 149940 158438 150198
rect 159054 149940 159082 150198
rect 159698 149940 159726 150198
rect 160342 149940 160370 150198
rect 160986 149940 161014 150198
rect 161630 149940 161658 150198
rect 162274 149940 162302 150198
rect 162918 149940 162946 150198
rect 163562 149940 163590 150198
rect 164206 149940 164234 150198
rect 164332 150204 164384 150210
rect 164804 150198 164878 150226
rect 164332 150146 164384 150152
rect 164850 149940 164878 150198
rect 165482 150204 165534 150210
rect 166092 150198 166166 150226
rect 166736 150198 166810 150226
rect 167380 150198 167454 150226
rect 168024 150198 168098 150226
rect 168484 150210 168512 155479
rect 168656 155450 168708 155456
rect 169392 155508 169444 155514
rect 169392 155450 169444 155456
rect 168668 150226 168696 155450
rect 169772 151842 169800 159054
rect 171980 158642 172008 163200
rect 172152 159180 172204 159186
rect 172152 159122 172204 159128
rect 170312 158636 170364 158642
rect 170312 158578 170364 158584
rect 171968 158636 172020 158642
rect 171968 158578 172020 158584
rect 169944 152176 169996 152182
rect 169944 152118 169996 152124
rect 169760 151836 169812 151842
rect 169760 151778 169812 151784
rect 169956 150226 169984 152118
rect 170324 151814 170352 158578
rect 171784 158500 171836 158506
rect 171784 158442 171836 158448
rect 171796 157962 171824 158442
rect 171784 157956 171836 157962
rect 171784 157898 171836 157904
rect 171876 157956 171928 157962
rect 171876 157898 171928 157904
rect 171888 157842 171916 157898
rect 171796 157826 171916 157842
rect 171784 157820 171916 157826
rect 171836 157814 171916 157820
rect 171784 157762 171836 157768
rect 171140 157208 171192 157214
rect 171140 157150 171192 157156
rect 170324 151786 170628 151814
rect 170600 150226 170628 151786
rect 165482 150146 165534 150152
rect 165494 149940 165522 150146
rect 166138 149940 166166 150198
rect 166782 149940 166810 150198
rect 167426 149940 167454 150198
rect 168070 149940 168098 150198
rect 168472 150204 168524 150210
rect 168668 150198 168742 150226
rect 168472 150146 168524 150152
rect 168714 149940 168742 150198
rect 169346 150204 169398 150210
rect 169956 150198 170030 150226
rect 170600 150198 170674 150226
rect 171152 150210 171180 157150
rect 171230 155272 171286 155281
rect 171230 155207 171286 155216
rect 171244 150226 171272 155207
rect 172164 152182 172192 159122
rect 172532 154222 172560 163254
rect 172716 163146 172744 163254
rect 172794 163200 172850 164400
rect 173622 163200 173678 164400
rect 173912 163254 174400 163282
rect 172808 163146 172836 163200
rect 172716 163118 172836 163146
rect 173256 159792 173308 159798
rect 173256 159734 173308 159740
rect 173072 158432 173124 158438
rect 173164 158432 173216 158438
rect 173072 158374 173124 158380
rect 173162 158400 173164 158409
rect 173216 158400 173218 158409
rect 172704 155644 172756 155650
rect 172704 155586 172756 155592
rect 172520 154216 172572 154222
rect 172520 154158 172572 154164
rect 172152 152176 172204 152182
rect 172152 152118 172204 152124
rect 172520 152040 172572 152046
rect 172520 151982 172572 151988
rect 172532 150226 172560 151982
rect 169346 150146 169398 150152
rect 169358 149940 169386 150146
rect 170002 149940 170030 150198
rect 170646 149940 170674 150198
rect 171140 150204 171192 150210
rect 171244 150198 171318 150226
rect 171140 150146 171192 150152
rect 171290 149940 171318 150198
rect 171922 150204 171974 150210
rect 172532 150198 172606 150226
rect 172716 150210 172744 155586
rect 173084 151814 173112 158374
rect 173162 158335 173218 158344
rect 173268 152454 173296 159734
rect 173636 159118 173664 163200
rect 173624 159112 173676 159118
rect 173624 159054 173676 159060
rect 173912 152862 173940 163254
rect 174372 163146 174400 163254
rect 174450 163200 174506 164400
rect 175278 163200 175334 164400
rect 176106 163200 176162 164400
rect 177026 163200 177082 164400
rect 177854 163200 177910 164400
rect 178682 163200 178738 164400
rect 179510 163200 179566 164400
rect 180338 163200 180394 164400
rect 180812 163254 181116 163282
rect 174464 163146 174492 163200
rect 174372 163118 174492 163146
rect 175292 158574 175320 163200
rect 175188 158568 175240 158574
rect 175188 158510 175240 158516
rect 175280 158568 175332 158574
rect 175280 158510 175332 158516
rect 175200 158386 175228 158510
rect 175200 158358 175320 158386
rect 175292 157334 175320 158358
rect 175292 157306 175412 157334
rect 174450 157040 174506 157049
rect 174450 156975 174506 156984
rect 173900 152856 173952 152862
rect 173900 152798 173952 152804
rect 173256 152448 173308 152454
rect 173256 152390 173308 152396
rect 173084 151786 173204 151814
rect 173176 150226 173204 151786
rect 174464 150226 174492 156975
rect 175096 153128 175148 153134
rect 175096 153070 175148 153076
rect 175108 150226 175136 153070
rect 175384 151814 175412 157306
rect 176120 155650 176148 163200
rect 176660 158772 176712 158778
rect 176660 158714 176712 158720
rect 176108 155644 176160 155650
rect 176108 155586 176160 155592
rect 176384 155576 176436 155582
rect 176384 155518 176436 155524
rect 175384 151786 175780 151814
rect 175752 150226 175780 151786
rect 176396 150226 176424 155518
rect 176672 153678 176700 158714
rect 177040 157214 177068 163200
rect 177868 159798 177896 163200
rect 177856 159792 177908 159798
rect 177856 159734 177908 159740
rect 178696 158506 178724 163200
rect 179420 159860 179472 159866
rect 179420 159802 179472 159808
rect 178040 158500 178092 158506
rect 178040 158442 178092 158448
rect 178684 158500 178736 158506
rect 178684 158442 178736 158448
rect 177028 157208 177080 157214
rect 177028 157150 177080 157156
rect 177026 155816 177082 155825
rect 177026 155751 177082 155760
rect 176660 153672 176712 153678
rect 176660 153614 176712 153620
rect 177040 150226 177068 155751
rect 177672 151972 177724 151978
rect 177672 151914 177724 151920
rect 177684 150226 177712 151914
rect 178052 151814 178080 158442
rect 179432 157826 179460 159802
rect 179420 157820 179472 157826
rect 179420 157762 179472 157768
rect 178958 155680 179014 155689
rect 178958 155615 179014 155624
rect 178052 151786 178356 151814
rect 178328 150226 178356 151786
rect 178972 150226 179000 155615
rect 179524 155582 179552 163200
rect 180352 158778 180380 163200
rect 180340 158772 180392 158778
rect 180340 158714 180392 158720
rect 179512 155576 179564 155582
rect 179512 155518 179564 155524
rect 179604 153604 179656 153610
rect 179604 153546 179656 153552
rect 179616 150226 179644 153546
rect 180812 153134 180840 163254
rect 181088 163146 181116 163254
rect 181166 163200 181222 164400
rect 181994 163200 182050 164400
rect 182192 163254 182864 163282
rect 181180 163146 181208 163200
rect 181088 163118 181208 163146
rect 182008 158710 182036 163200
rect 180892 158704 180944 158710
rect 180892 158646 180944 158652
rect 181996 158704 182048 158710
rect 181996 158646 182048 158652
rect 180800 153128 180852 153134
rect 180800 153070 180852 153076
rect 180248 152312 180300 152318
rect 180248 152254 180300 152260
rect 180260 150226 180288 152254
rect 180904 150226 180932 158646
rect 182088 156392 182140 156398
rect 182088 156334 182140 156340
rect 180984 155712 181036 155718
rect 180984 155654 181036 155660
rect 180996 151814 181024 155654
rect 180996 151786 181484 151814
rect 171922 150146 171974 150152
rect 171934 149940 171962 150146
rect 172578 149940 172606 150198
rect 172704 150204 172756 150210
rect 173176 150198 173250 150226
rect 172704 150146 172756 150152
rect 173222 149940 173250 150198
rect 173854 150204 173906 150210
rect 174464 150198 174538 150226
rect 175108 150198 175182 150226
rect 175752 150198 175826 150226
rect 176396 150198 176470 150226
rect 177040 150198 177114 150226
rect 177684 150198 177758 150226
rect 178328 150198 178402 150226
rect 178972 150198 179046 150226
rect 179616 150198 179690 150226
rect 180260 150198 180334 150226
rect 173854 150146 173906 150152
rect 173866 149940 173894 150146
rect 174510 149940 174538 150198
rect 175154 149940 175182 150198
rect 175798 149940 175826 150198
rect 176442 149940 176470 150198
rect 177086 149940 177114 150198
rect 177730 149940 177758 150198
rect 178374 149940 178402 150198
rect 179018 149940 179046 150198
rect 179662 149940 179690 150198
rect 180306 149940 180334 150198
rect 180858 150198 180932 150226
rect 181456 150226 181484 151786
rect 182100 150226 182128 156334
rect 182192 153678 182220 163254
rect 182836 163146 182864 163254
rect 182914 163200 182970 164400
rect 183742 163200 183798 164400
rect 184570 163200 184626 164400
rect 185398 163200 185454 164400
rect 186226 163200 186282 164400
rect 187054 163200 187110 164400
rect 187882 163200 187938 164400
rect 188802 163200 188858 164400
rect 189630 163200 189686 164400
rect 190458 163200 190514 164400
rect 191286 163200 191342 164400
rect 192114 163200 192170 164400
rect 192942 163200 192998 164400
rect 193770 163200 193826 164400
rect 194690 163200 194746 164400
rect 195518 163200 195574 164400
rect 196346 163200 196402 164400
rect 197174 163200 197230 164400
rect 198002 163200 198058 164400
rect 198830 163200 198886 164400
rect 199658 163200 199714 164400
rect 200578 163200 200634 164400
rect 201406 163200 201462 164400
rect 202234 163200 202290 164400
rect 203062 163200 203118 164400
rect 203890 163200 203946 164400
rect 204718 163200 204774 164400
rect 205008 163254 205496 163282
rect 182928 163146 182956 163200
rect 182836 163118 182956 163146
rect 183756 159050 183784 163200
rect 184584 159866 184612 163200
rect 184572 159860 184624 159866
rect 184572 159802 184624 159808
rect 184388 159248 184440 159254
rect 184388 159190 184440 159196
rect 183468 159044 183520 159050
rect 183468 158986 183520 158992
rect 183744 159044 183796 159050
rect 183744 158986 183796 158992
rect 182272 157956 182324 157962
rect 182272 157898 182324 157904
rect 182180 153672 182232 153678
rect 182180 153614 182232 153620
rect 181456 150198 181530 150226
rect 182100 150198 182174 150226
rect 182284 150210 182312 157898
rect 183480 152114 183508 158986
rect 184018 155952 184074 155961
rect 184018 155887 184074 155896
rect 182732 152108 182784 152114
rect 182732 152050 182784 152056
rect 183468 152108 183520 152114
rect 183468 152050 183520 152056
rect 182744 150226 182772 152050
rect 184032 150226 184060 155887
rect 184400 151978 184428 159190
rect 185412 157962 185440 163200
rect 185308 157956 185360 157962
rect 185308 157898 185360 157904
rect 185400 157956 185452 157962
rect 185400 157898 185452 157904
rect 185124 157888 185176 157894
rect 185124 157830 185176 157836
rect 185320 157842 185348 157898
rect 185136 155258 185164 157830
rect 185320 157814 185624 157842
rect 185308 157752 185360 157758
rect 185308 157694 185360 157700
rect 185320 157570 185348 157694
rect 185596 157690 185624 157814
rect 185676 157752 185728 157758
rect 185676 157694 185728 157700
rect 185584 157684 185636 157690
rect 185584 157626 185636 157632
rect 185688 157570 185716 157694
rect 185320 157542 185716 157570
rect 186240 155718 186268 163200
rect 186412 159928 186464 159934
rect 186412 159870 186464 159876
rect 186424 157334 186452 159870
rect 187068 159254 187096 163200
rect 187896 161474 187924 163200
rect 187896 161446 188016 161474
rect 187056 159248 187108 159254
rect 187056 159190 187108 159196
rect 186424 157306 186728 157334
rect 186320 155848 186372 155854
rect 186320 155790 186372 155796
rect 186412 155848 186464 155854
rect 186412 155790 186464 155796
rect 186228 155712 186280 155718
rect 186228 155654 186280 155660
rect 185136 155230 185992 155258
rect 184662 154456 184718 154465
rect 184662 154391 184718 154400
rect 185400 154420 185452 154426
rect 184388 151972 184440 151978
rect 184388 151914 184440 151920
rect 184676 150226 184704 154391
rect 185400 154362 185452 154368
rect 185860 154420 185912 154426
rect 185860 154362 185912 154368
rect 185412 154306 185440 154362
rect 185412 154290 185808 154306
rect 185308 154284 185360 154290
rect 185412 154284 185820 154290
rect 185412 154278 185768 154284
rect 185308 154226 185360 154232
rect 185768 154226 185820 154232
rect 185320 154170 185348 154226
rect 185872 154170 185900 154362
rect 185320 154142 185900 154170
rect 185308 151836 185360 151842
rect 185308 151778 185360 151784
rect 185320 150226 185348 151778
rect 185964 150226 185992 155230
rect 186332 155145 186360 155790
rect 186318 155136 186374 155145
rect 186318 155071 186374 155080
rect 186320 155032 186372 155038
rect 186424 155020 186452 155790
rect 186372 154992 186452 155020
rect 186320 154974 186372 154980
rect 186700 154902 186728 157306
rect 186872 155916 186924 155922
rect 186872 155858 186924 155864
rect 186780 155100 186832 155106
rect 186780 155042 186832 155048
rect 186412 154896 186464 154902
rect 186412 154838 186464 154844
rect 186688 154896 186740 154902
rect 186688 154838 186740 154844
rect 186424 154714 186452 154838
rect 186792 154714 186820 155042
rect 186424 154686 186820 154714
rect 186884 154408 186912 155858
rect 187238 155136 187294 155145
rect 187238 155071 187294 155080
rect 186700 154380 186912 154408
rect 186700 150226 186728 154380
rect 186872 154284 186924 154290
rect 186872 154226 186924 154232
rect 186964 154284 187016 154290
rect 186964 154226 187016 154232
rect 186884 154193 186912 154226
rect 186870 154184 186926 154193
rect 186870 154119 186926 154128
rect 186976 153678 187004 154226
rect 186964 153672 187016 153678
rect 186964 153614 187016 153620
rect 180858 149940 180886 150198
rect 181502 149940 181530 150198
rect 182146 149940 182174 150198
rect 182272 150204 182324 150210
rect 182744 150198 182818 150226
rect 182272 150146 182324 150152
rect 182790 149940 182818 150198
rect 183422 150204 183474 150210
rect 184032 150198 184106 150226
rect 184676 150198 184750 150226
rect 185320 150198 185394 150226
rect 185964 150198 186038 150226
rect 183422 150146 183474 150152
rect 183434 149940 183462 150146
rect 184078 149940 184106 150198
rect 184722 149940 184750 150198
rect 185366 149940 185394 150198
rect 186010 149940 186038 150198
rect 186654 150198 186728 150226
rect 186654 149940 186682 150198
rect 187252 150090 187280 155071
rect 187884 152992 187936 152998
rect 187884 152934 187936 152940
rect 187896 150090 187924 152934
rect 187988 152318 188016 161446
rect 188816 157894 188844 163200
rect 188804 157888 188856 157894
rect 188804 157830 188856 157836
rect 188528 157752 188580 157758
rect 188528 157694 188580 157700
rect 188436 154488 188488 154494
rect 188436 154430 188488 154436
rect 188448 153678 188476 154430
rect 188436 153672 188488 153678
rect 188436 153614 188488 153620
rect 187976 152312 188028 152318
rect 187976 152254 188028 152260
rect 188540 150226 188568 157694
rect 189644 155854 189672 163200
rect 190472 157758 190500 163200
rect 191300 159934 191328 163200
rect 191748 160064 191800 160070
rect 191748 160006 191800 160012
rect 191472 159996 191524 160002
rect 191472 159938 191524 159944
rect 191288 159928 191340 159934
rect 191288 159870 191340 159876
rect 190644 157820 190696 157826
rect 190644 157762 190696 157768
rect 190460 157752 190512 157758
rect 190460 157694 190512 157700
rect 190656 157334 190684 157762
rect 190656 157306 191144 157334
rect 189540 155848 189592 155854
rect 189540 155790 189592 155796
rect 189632 155848 189684 155854
rect 189632 155790 189684 155796
rect 189552 155174 189580 155790
rect 189172 155168 189224 155174
rect 189172 155110 189224 155116
rect 189540 155168 189592 155174
rect 189540 155110 189592 155116
rect 188540 150198 188614 150226
rect 187252 150062 187326 150090
rect 187896 150062 187970 150090
rect 187298 149940 187326 150062
rect 187942 149940 187970 150062
rect 188586 149940 188614 150198
rect 189184 150090 189212 155110
rect 191012 154420 191064 154426
rect 191012 154362 191064 154368
rect 189814 154184 189870 154193
rect 189814 154119 189870 154128
rect 189828 150090 189856 154119
rect 191024 153406 191052 154362
rect 191012 153400 191064 153406
rect 191012 153342 191064 153348
rect 190460 152176 190512 152182
rect 190460 152118 190512 152124
rect 190472 150090 190500 152118
rect 191116 150226 191144 157306
rect 191484 152046 191512 159938
rect 191760 157334 191788 160006
rect 191668 157306 191788 157334
rect 191668 153406 191696 157306
rect 192128 157282 192156 163200
rect 192116 157276 192168 157282
rect 192116 157218 192168 157224
rect 192956 155922 192984 163200
rect 193784 159186 193812 163200
rect 193772 159180 193824 159186
rect 193772 159122 193824 159128
rect 194140 158976 194192 158982
rect 194140 158918 194192 158924
rect 193220 157616 193272 157622
rect 193220 157558 193272 157564
rect 193232 157334 193260 157558
rect 193232 157306 193720 157334
rect 192944 155916 192996 155922
rect 192944 155858 192996 155864
rect 191748 155032 191800 155038
rect 191748 154974 191800 154980
rect 191656 153400 191708 153406
rect 191656 153342 191708 153348
rect 191472 152040 191524 152046
rect 191472 151982 191524 151988
rect 191116 150198 191190 150226
rect 189184 150062 189258 150090
rect 189828 150062 189902 150090
rect 190472 150062 190546 150090
rect 189230 149940 189258 150062
rect 189874 149940 189902 150062
rect 190518 149940 190546 150062
rect 191162 149940 191190 150198
rect 191760 150090 191788 154974
rect 192390 153776 192446 153785
rect 192390 153711 192446 153720
rect 192404 150090 192432 153711
rect 193036 152924 193088 152930
rect 193036 152866 193088 152872
rect 193048 150090 193076 152866
rect 193692 150226 193720 157306
rect 194152 152182 194180 158918
rect 194704 158914 194732 163200
rect 194600 158908 194652 158914
rect 194600 158850 194652 158856
rect 194692 158908 194744 158914
rect 194692 158850 194744 158856
rect 194324 155168 194376 155174
rect 194324 155110 194376 155116
rect 194140 152176 194192 152182
rect 194140 152118 194192 152124
rect 193692 150198 193766 150226
rect 191760 150062 191834 150090
rect 192404 150062 192478 150090
rect 193048 150062 193122 150090
rect 191806 149940 191834 150062
rect 192450 149940 192478 150062
rect 193094 149940 193122 150062
rect 193738 149940 193766 150198
rect 194336 150090 194364 155110
rect 194612 152998 194640 158850
rect 195532 157826 195560 163200
rect 195980 158840 196032 158846
rect 195980 158782 196032 158788
rect 195520 157820 195572 157826
rect 195520 157762 195572 157768
rect 195992 156330 196020 158782
rect 194968 156324 195020 156330
rect 194968 156266 195020 156272
rect 195980 156324 196032 156330
rect 195980 156266 196032 156272
rect 194600 152992 194652 152998
rect 194600 152934 194652 152940
rect 194980 150090 195008 156266
rect 196256 156256 196308 156262
rect 196256 156198 196308 156204
rect 195980 153672 196032 153678
rect 195886 153640 195942 153649
rect 196072 153672 196124 153678
rect 195980 153614 196032 153620
rect 196070 153640 196072 153649
rect 196124 153640 196126 153649
rect 195886 153575 195942 153584
rect 195900 153406 195928 153575
rect 195992 153406 196020 153614
rect 196070 153575 196126 153584
rect 195888 153400 195940 153406
rect 195888 153342 195940 153348
rect 195980 153400 196032 153406
rect 195980 153342 196032 153348
rect 195612 151972 195664 151978
rect 195612 151914 195664 151920
rect 195624 150090 195652 151914
rect 196268 150090 196296 156198
rect 196360 155174 196388 163200
rect 197188 160070 197216 163200
rect 197176 160064 197228 160070
rect 197176 160006 197228 160012
rect 198016 160002 198044 163200
rect 198004 159996 198056 160002
rect 198004 159938 198056 159944
rect 197360 159112 197412 159118
rect 197360 159054 197412 159060
rect 197372 157622 197400 159054
rect 198738 158536 198794 158545
rect 198738 158471 198794 158480
rect 197360 157616 197412 157622
rect 197360 157558 197412 157564
rect 196992 156324 197044 156330
rect 196992 156266 197044 156272
rect 196348 155168 196400 155174
rect 196348 155110 196400 155116
rect 196900 153536 196952 153542
rect 196900 153478 196952 153484
rect 196532 153468 196584 153474
rect 196532 153410 196584 153416
rect 196544 150210 196572 153410
rect 196532 150204 196584 150210
rect 196532 150146 196584 150152
rect 196912 150090 196940 153478
rect 197004 153474 197032 156266
rect 198004 156256 198056 156262
rect 198004 156198 198056 156204
rect 198016 156058 198044 156198
rect 198004 156052 198056 156058
rect 198004 155994 198056 156000
rect 196992 153468 197044 153474
rect 196992 153410 197044 153416
rect 197544 153400 197596 153406
rect 197544 153342 197596 153348
rect 197556 150090 197584 153342
rect 198188 153060 198240 153066
rect 198188 153002 198240 153008
rect 198200 150090 198228 153002
rect 198752 150226 198780 158471
rect 198844 156398 198872 163200
rect 198924 159316 198976 159322
rect 198924 159258 198976 159264
rect 198832 156392 198884 156398
rect 198832 156334 198884 156340
rect 198936 153542 198964 159258
rect 199672 155106 199700 163200
rect 200592 158982 200620 163200
rect 201420 159322 201448 163200
rect 201408 159316 201460 159322
rect 201408 159258 201460 159264
rect 201408 159044 201460 159050
rect 201408 158986 201460 158992
rect 200580 158976 200632 158982
rect 200580 158918 200632 158924
rect 200764 156596 200816 156602
rect 200764 156538 200816 156544
rect 200948 156596 201000 156602
rect 200948 156538 201000 156544
rect 200776 156330 200804 156538
rect 200960 156398 200988 156538
rect 200948 156392 201000 156398
rect 200948 156334 201000 156340
rect 200764 156324 200816 156330
rect 200764 156266 200816 156272
rect 200672 156188 200724 156194
rect 200672 156130 200724 156136
rect 199660 155100 199712 155106
rect 199660 155042 199712 155048
rect 200120 155032 200172 155038
rect 200120 154974 200172 154980
rect 198924 153536 198976 153542
rect 198924 153478 198976 153484
rect 198752 150198 198918 150226
rect 194336 150062 194410 150090
rect 194980 150062 195054 150090
rect 195624 150062 195698 150090
rect 196268 150062 196342 150090
rect 196912 150062 196986 150090
rect 197556 150062 197630 150090
rect 198200 150062 198274 150090
rect 194382 149940 194410 150062
rect 195026 149940 195054 150062
rect 195670 149940 195698 150062
rect 196314 149940 196342 150062
rect 196958 149940 196986 150062
rect 197602 149940 197630 150062
rect 198246 149940 198274 150062
rect 198890 149940 198918 150198
rect 199522 150204 199574 150210
rect 199522 150146 199574 150152
rect 199534 149940 199562 150146
rect 200132 150090 200160 154974
rect 200684 152266 200712 156130
rect 201420 153474 201448 158986
rect 202248 156058 202276 163200
rect 203076 156126 203104 163200
rect 203904 159118 203932 163200
rect 204732 159361 204760 163200
rect 204718 159352 204774 159361
rect 204718 159287 204774 159296
rect 203892 159112 203944 159118
rect 203892 159054 203944 159060
rect 203708 158908 203760 158914
rect 203708 158850 203760 158856
rect 203432 157548 203484 157554
rect 203432 157490 203484 157496
rect 203444 157334 203472 157490
rect 203444 157306 203656 157334
rect 203064 156120 203116 156126
rect 203064 156062 203116 156068
rect 202236 156052 202288 156058
rect 202236 155994 202288 156000
rect 202696 154488 202748 154494
rect 202696 154430 202748 154436
rect 202052 154420 202104 154426
rect 202052 154362 202104 154368
rect 201408 153468 201460 153474
rect 201408 153410 201460 153416
rect 200684 152238 201448 152266
rect 200764 152108 200816 152114
rect 200764 152050 200816 152056
rect 200776 150090 200804 152050
rect 201420 150226 201448 152238
rect 201420 150198 201494 150226
rect 200132 150062 200206 150090
rect 200776 150062 200850 150090
rect 200178 149940 200206 150062
rect 200822 149940 200850 150062
rect 201466 149940 201494 150198
rect 202064 150090 202092 154362
rect 202708 150090 202736 154430
rect 203340 151904 203392 151910
rect 203340 151846 203392 151852
rect 203352 150090 203380 151846
rect 203628 150226 203656 157306
rect 203720 153066 203748 158850
rect 204904 158772 204956 158778
rect 204904 158714 204956 158720
rect 204916 157554 204944 158714
rect 204904 157548 204956 157554
rect 204904 157490 204956 157496
rect 204628 155780 204680 155786
rect 204628 155722 204680 155728
rect 203708 153060 203760 153066
rect 203708 153002 203760 153008
rect 203628 150198 204070 150226
rect 202064 150062 202138 150090
rect 202708 150062 202782 150090
rect 203352 150062 203426 150090
rect 202110 149940 202138 150062
rect 202754 149940 202782 150062
rect 203398 149940 203426 150062
rect 204042 149940 204070 150198
rect 204640 150090 204668 155722
rect 205008 154426 205036 163254
rect 205468 163146 205496 163254
rect 205546 163200 205602 164400
rect 206466 163200 206522 164400
rect 207294 163200 207350 164400
rect 208122 163200 208178 164400
rect 208412 163254 208900 163282
rect 205560 163146 205588 163200
rect 205468 163118 205588 163146
rect 206480 155786 206508 163200
rect 207020 160064 207072 160070
rect 207020 160006 207072 160012
rect 206560 157480 206612 157486
rect 206560 157422 206612 157428
rect 206468 155780 206520 155786
rect 206468 155722 206520 155728
rect 204996 154420 205048 154426
rect 204996 154362 205048 154368
rect 205272 154352 205324 154358
rect 205272 154294 205324 154300
rect 205284 150090 205312 154294
rect 205916 153196 205968 153202
rect 205916 153138 205968 153144
rect 205928 150090 205956 153138
rect 206572 150226 206600 157422
rect 207032 155038 207060 160006
rect 207308 158846 207336 163200
rect 208136 158914 208164 163200
rect 208124 158908 208176 158914
rect 208124 158850 208176 158856
rect 207296 158840 207348 158846
rect 207296 158782 207348 158788
rect 207202 157176 207258 157185
rect 207202 157111 207258 157120
rect 207020 155032 207072 155038
rect 207020 154974 207072 154980
rect 206572 150198 206646 150226
rect 204640 150062 204714 150090
rect 205284 150062 205358 150090
rect 205928 150062 206002 150090
rect 204686 149940 204714 150062
rect 205330 149940 205358 150062
rect 205974 149940 206002 150062
rect 206618 149940 206646 150198
rect 207216 150090 207244 157111
rect 208412 154358 208440 163254
rect 208872 163146 208900 163254
rect 208950 163200 209006 164400
rect 209778 163200 209834 164400
rect 210606 163200 210662 164400
rect 211434 163200 211490 164400
rect 211540 163254 212304 163282
rect 208964 163146 208992 163200
rect 208872 163118 208992 163146
rect 209792 157334 209820 163200
rect 210620 158778 210648 163200
rect 211448 160070 211476 163200
rect 211436 160064 211488 160070
rect 211436 160006 211488 160012
rect 210608 158772 210660 158778
rect 210608 158714 210660 158720
rect 210516 157344 210568 157350
rect 209792 157306 209912 157334
rect 209778 156768 209834 156777
rect 209778 156703 209834 156712
rect 209792 156670 209820 156703
rect 209780 156664 209832 156670
rect 209780 156606 209832 156612
rect 209884 156398 209912 157306
rect 210516 157286 210568 157292
rect 210424 156868 210476 156874
rect 210424 156810 210476 156816
rect 209964 156664 210016 156670
rect 209964 156606 210016 156612
rect 209872 156392 209924 156398
rect 209872 156334 209924 156340
rect 209976 156262 210004 156606
rect 210436 156330 210464 156810
rect 210424 156324 210476 156330
rect 210424 156266 210476 156272
rect 210528 156262 210556 157286
rect 210608 156868 210660 156874
rect 210608 156810 210660 156816
rect 210620 156777 210648 156810
rect 210606 156768 210662 156777
rect 210606 156703 210662 156712
rect 209964 156256 210016 156262
rect 209964 156198 210016 156204
rect 210516 156256 210568 156262
rect 210516 156198 210568 156204
rect 209136 156188 209188 156194
rect 209136 156130 209188 156136
rect 208400 154352 208452 154358
rect 208400 154294 208452 154300
rect 207848 153264 207900 153270
rect 207848 153206 207900 153212
rect 207860 150090 207888 153206
rect 208492 152040 208544 152046
rect 208492 151982 208544 151988
rect 208504 150090 208532 151982
rect 209148 150090 209176 156130
rect 211540 153785 211568 163254
rect 212276 163146 212304 163254
rect 212354 163200 212410 164400
rect 213182 163200 213238 164400
rect 214010 163200 214066 164400
rect 214838 163200 214894 164400
rect 215312 163254 215616 163282
rect 212368 163146 212396 163200
rect 212276 163118 212396 163146
rect 213196 160274 213224 163200
rect 213184 160268 213236 160274
rect 213184 160210 213236 160216
rect 214024 159322 214052 163200
rect 212632 159316 212684 159322
rect 212632 159258 212684 159264
rect 214012 159316 214064 159322
rect 214012 159258 214064 159264
rect 212448 158908 212500 158914
rect 212448 158850 212500 158856
rect 211620 156664 211672 156670
rect 211620 156606 211672 156612
rect 211526 153776 211582 153785
rect 210424 153740 210476 153746
rect 211526 153711 211582 153720
rect 210424 153682 210476 153688
rect 209780 153332 209832 153338
rect 209780 153274 209832 153280
rect 209792 150090 209820 153274
rect 210436 150090 210464 153682
rect 211068 152380 211120 152386
rect 211068 152322 211120 152328
rect 211080 150090 211108 152322
rect 211632 150090 211660 156606
rect 212264 154964 212316 154970
rect 212264 154906 212316 154912
rect 212276 150090 212304 154906
rect 212460 152930 212488 158850
rect 212448 152924 212500 152930
rect 212448 152866 212500 152872
rect 212644 152046 212672 159258
rect 214656 159248 214708 159254
rect 214656 159190 214708 159196
rect 212724 159112 212776 159118
rect 212724 159054 212776 159060
rect 212736 152114 212764 159054
rect 214564 157480 214616 157486
rect 214392 157440 214564 157468
rect 214392 157350 214420 157440
rect 214564 157422 214616 157428
rect 214380 157344 214432 157350
rect 214380 157286 214432 157292
rect 214196 156868 214248 156874
rect 214196 156810 214248 156816
rect 212908 154556 212960 154562
rect 212908 154498 212960 154504
rect 212724 152108 212776 152114
rect 212724 152050 212776 152056
rect 212632 152040 212684 152046
rect 212632 151982 212684 151988
rect 212920 150090 212948 154498
rect 213552 152176 213604 152182
rect 213552 152118 213604 152124
rect 213564 150090 213592 152118
rect 214208 150090 214236 156810
rect 214668 154970 214696 159190
rect 214852 159050 214880 163200
rect 214840 159044 214892 159050
rect 214840 158986 214892 158992
rect 214656 154964 214708 154970
rect 214656 154906 214708 154912
rect 214840 154828 214892 154834
rect 214840 154770 214892 154776
rect 214852 150090 214880 154770
rect 215312 154562 215340 163254
rect 215588 163146 215616 163254
rect 215666 163200 215722 164400
rect 216494 163200 216550 164400
rect 217322 163200 217378 164400
rect 218242 163200 218298 164400
rect 218348 163254 219020 163282
rect 215680 163146 215708 163200
rect 215588 163118 215708 163146
rect 215392 158772 215444 158778
rect 215392 158714 215444 158720
rect 215300 154556 215352 154562
rect 215300 154498 215352 154504
rect 215404 153202 215432 158714
rect 216508 156670 216536 163200
rect 217336 158846 217364 163200
rect 218256 159254 218284 163200
rect 218244 159248 218296 159254
rect 218244 159190 218296 159196
rect 218060 159180 218112 159186
rect 218060 159122 218112 159128
rect 217324 158840 217376 158846
rect 217324 158782 217376 158788
rect 216772 156732 216824 156738
rect 216772 156674 216824 156680
rect 216496 156664 216548 156670
rect 216496 156606 216548 156612
rect 215484 156188 215536 156194
rect 215484 156130 215536 156136
rect 215392 153196 215444 153202
rect 215392 153138 215444 153144
rect 215496 150226 215524 156130
rect 216128 152516 216180 152522
rect 216128 152458 216180 152464
rect 216140 150226 216168 152458
rect 216784 150226 216812 156674
rect 218072 156194 218100 159122
rect 218060 156188 218112 156194
rect 218060 156130 218112 156136
rect 217416 155236 217468 155242
rect 217416 155178 217468 155184
rect 217428 150226 217456 155178
rect 218348 154494 218376 163254
rect 218992 163146 219020 163254
rect 219070 163200 219126 164400
rect 219898 163200 219954 164400
rect 220726 163200 220782 164400
rect 221554 163200 221610 164400
rect 222382 163200 222438 164400
rect 223210 163200 223266 164400
rect 224130 163200 224186 164400
rect 224958 163200 225014 164400
rect 225248 163254 225736 163282
rect 219084 163146 219112 163200
rect 218992 163118 219112 163146
rect 219348 158024 219400 158030
rect 219348 157966 219400 157972
rect 218336 154488 218388 154494
rect 218336 154430 218388 154436
rect 218060 153808 218112 153814
rect 218060 153750 218112 153756
rect 218072 150226 218100 153750
rect 218704 152992 218756 152998
rect 218704 152934 218756 152940
rect 218716 150226 218744 152934
rect 219360 150226 219388 157966
rect 219716 156868 219768 156874
rect 219716 156810 219768 156816
rect 219728 156466 219756 156810
rect 219716 156460 219768 156466
rect 219716 156402 219768 156408
rect 219808 156460 219860 156466
rect 219808 156402 219860 156408
rect 219820 156330 219848 156402
rect 219912 156330 219940 163200
rect 220740 159118 220768 163200
rect 221188 160268 221240 160274
rect 221188 160210 221240 160216
rect 220728 159112 220780 159118
rect 220728 159054 220780 159060
rect 220360 158840 220412 158846
rect 220360 158782 220412 158788
rect 219808 156324 219860 156330
rect 219808 156266 219860 156272
rect 219900 156324 219952 156330
rect 219900 156266 219952 156272
rect 219992 156256 220044 156262
rect 219992 156198 220044 156204
rect 219900 154012 219952 154018
rect 219900 153954 219952 153960
rect 215496 150198 215570 150226
rect 216140 150198 216214 150226
rect 216784 150198 216858 150226
rect 217428 150198 217502 150226
rect 218072 150198 218146 150226
rect 218716 150198 218790 150226
rect 219360 150198 219434 150226
rect 207216 150062 207290 150090
rect 207860 150062 207934 150090
rect 208504 150062 208578 150090
rect 209148 150062 209222 150090
rect 209792 150062 209866 150090
rect 210436 150062 210510 150090
rect 211080 150062 211154 150090
rect 211632 150062 211706 150090
rect 212276 150062 212350 150090
rect 212920 150062 212994 150090
rect 213564 150062 213638 150090
rect 214208 150062 214282 150090
rect 214852 150062 214926 150090
rect 207262 149940 207290 150062
rect 207906 149940 207934 150062
rect 208550 149940 208578 150062
rect 209194 149940 209222 150062
rect 209838 149940 209866 150062
rect 210482 149940 210510 150062
rect 211126 149940 211154 150062
rect 211678 149940 211706 150062
rect 212322 149940 212350 150062
rect 212966 149940 212994 150062
rect 213610 149940 213638 150062
rect 214254 149940 214282 150062
rect 214898 149940 214926 150062
rect 215542 149940 215570 150198
rect 216186 149940 216214 150198
rect 216830 149940 216858 150198
rect 217474 149940 217502 150198
rect 218118 149940 218146 150198
rect 218762 149940 218790 150198
rect 219406 149940 219434 150198
rect 219912 150192 219940 153954
rect 220004 151814 220032 156198
rect 220372 152998 220400 158782
rect 221200 157350 221228 160210
rect 221568 158778 221596 163200
rect 222108 159044 222160 159050
rect 222108 158986 222160 158992
rect 221556 158772 221608 158778
rect 221556 158714 221608 158720
rect 221188 157344 221240 157350
rect 221188 157286 221240 157292
rect 221372 156460 221424 156466
rect 221372 156402 221424 156408
rect 220360 152992 220412 152998
rect 220360 152934 220412 152940
rect 221280 152244 221332 152250
rect 221280 152186 221332 152192
rect 220004 151786 220676 151814
rect 220648 150226 220676 151786
rect 221292 150226 221320 152186
rect 221384 151814 221412 156402
rect 222120 152250 222148 158986
rect 222396 154018 222424 163200
rect 222568 156936 222620 156942
rect 222568 156878 222620 156884
rect 222384 154012 222436 154018
rect 222384 153954 222436 153960
rect 222108 152244 222160 152250
rect 222108 152186 222160 152192
rect 221384 151786 221964 151814
rect 221936 150226 221964 151786
rect 222580 150226 222608 156878
rect 223224 156738 223252 163200
rect 223580 159384 223632 159390
rect 223580 159326 223632 159332
rect 223212 156732 223264 156738
rect 223212 156674 223264 156680
rect 223212 153944 223264 153950
rect 223212 153886 223264 153892
rect 223224 150226 223252 153886
rect 223592 151814 223620 159326
rect 224144 159050 224172 163200
rect 224972 159186 225000 163200
rect 224960 159180 225012 159186
rect 224960 159122 225012 159128
rect 224132 159044 224184 159050
rect 224132 158986 224184 158992
rect 224960 158976 225012 158982
rect 224960 158918 225012 158924
rect 224408 158772 224460 158778
rect 224408 158714 224460 158720
rect 224132 157004 224184 157010
rect 224132 156946 224184 156952
rect 224144 151814 224172 156946
rect 224420 152386 224448 158714
rect 224972 156942 225000 158918
rect 224960 156936 225012 156942
rect 224960 156878 225012 156884
rect 225144 156800 225196 156806
rect 225144 156742 225196 156748
rect 225052 156528 225104 156534
rect 225052 156470 225104 156476
rect 224408 152380 224460 152386
rect 224408 152322 224460 152328
rect 223592 151786 223896 151814
rect 224144 151786 224540 151814
rect 223868 150226 223896 151786
rect 224512 150226 224540 151786
rect 220648 150198 220722 150226
rect 221292 150198 221366 150226
rect 221936 150198 222010 150226
rect 222580 150198 222654 150226
rect 223224 150198 223298 150226
rect 223868 150198 223942 150226
rect 224512 150198 224586 150226
rect 225064 150210 225092 156470
rect 225156 150226 225184 156742
rect 225248 153950 225276 163254
rect 225708 163146 225736 163254
rect 225786 163200 225842 164400
rect 226614 163200 226670 164400
rect 227442 163200 227498 164400
rect 227732 163254 228220 163282
rect 225800 163146 225828 163200
rect 225708 163118 225828 163146
rect 225328 159520 225380 159526
rect 225328 159462 225380 159468
rect 225236 153944 225288 153950
rect 225236 153886 225288 153892
rect 225340 152182 225368 159462
rect 226628 156874 226656 163200
rect 227076 157412 227128 157418
rect 227076 157354 227128 157360
rect 226616 156868 226668 156874
rect 226616 156810 226668 156816
rect 226432 152584 226484 152590
rect 226432 152526 226484 152532
rect 225328 152176 225380 152182
rect 225328 152118 225380 152124
rect 226444 150226 226472 152526
rect 227088 150226 227116 157354
rect 227456 152425 227484 163200
rect 227732 152522 227760 163254
rect 228192 163146 228220 163254
rect 228270 163200 228326 164400
rect 229098 163200 229154 164400
rect 230018 163200 230074 164400
rect 230846 163200 230902 164400
rect 231674 163200 231730 164400
rect 231872 163254 232452 163282
rect 228284 163146 228312 163200
rect 228192 163118 228312 163146
rect 228364 156800 228416 156806
rect 228364 156742 228416 156748
rect 227812 155304 227864 155310
rect 227812 155246 227864 155252
rect 227720 152516 227772 152522
rect 227720 152458 227772 152464
rect 227442 152416 227498 152425
rect 227442 152351 227498 152360
rect 227824 150226 227852 155246
rect 219912 150164 220078 150192
rect 220050 149940 220078 150164
rect 220694 149940 220722 150198
rect 221338 149940 221366 150198
rect 221982 149940 222010 150198
rect 222626 149940 222654 150198
rect 223270 149940 223298 150198
rect 223914 149940 223942 150198
rect 224558 149940 224586 150198
rect 225052 150204 225104 150210
rect 225156 150198 225230 150226
rect 225052 150146 225104 150152
rect 225202 149940 225230 150198
rect 225834 150204 225886 150210
rect 226444 150198 226518 150226
rect 227088 150198 227162 150226
rect 225834 150146 225886 150152
rect 225846 149940 225874 150146
rect 226490 149940 226518 150198
rect 227134 149940 227162 150198
rect 227778 150198 227852 150226
rect 228376 150226 228404 156742
rect 229112 153746 229140 163200
rect 230032 156806 230060 163200
rect 230860 159526 230888 163200
rect 230848 159520 230900 159526
rect 230848 159462 230900 159468
rect 231688 159390 231716 163200
rect 231676 159384 231728 159390
rect 231676 159326 231728 159332
rect 230756 158908 230808 158914
rect 230756 158850 230808 158856
rect 230020 156800 230072 156806
rect 230020 156742 230072 156748
rect 230768 156194 230796 158850
rect 230756 156188 230808 156194
rect 230756 156130 230808 156136
rect 229652 155984 229704 155990
rect 229652 155926 229704 155932
rect 229192 155372 229244 155378
rect 229192 155314 229244 155320
rect 229100 153740 229152 153746
rect 229100 153682 229152 153688
rect 229008 152176 229060 152182
rect 229008 152118 229060 152124
rect 229020 150226 229048 152118
rect 228376 150198 228450 150226
rect 229020 150198 229094 150226
rect 229204 150210 229232 155314
rect 229664 150226 229692 155926
rect 231872 153814 231900 163254
rect 232424 163146 232452 163254
rect 232502 163200 232558 164400
rect 233330 163200 233386 164400
rect 234158 163200 234214 164400
rect 234986 163200 235042 164400
rect 235092 163254 235856 163282
rect 232516 163146 232544 163200
rect 232424 163118 232544 163146
rect 233240 159452 233292 159458
rect 233240 159394 233292 159400
rect 231952 158092 232004 158098
rect 231952 158034 232004 158040
rect 231860 153808 231912 153814
rect 231860 153750 231912 153756
rect 230940 153604 230992 153610
rect 230940 153546 230992 153552
rect 230952 150226 230980 153546
rect 231584 152720 231636 152726
rect 231584 152662 231636 152668
rect 231596 150226 231624 152662
rect 231964 151814 231992 158034
rect 232872 155440 232924 155446
rect 232872 155382 232924 155388
rect 231964 151786 232268 151814
rect 232240 150226 232268 151786
rect 232884 150226 232912 155382
rect 227778 149940 227806 150198
rect 228422 149940 228450 150198
rect 229066 149940 229094 150198
rect 229192 150204 229244 150210
rect 229664 150198 229738 150226
rect 229192 150146 229244 150152
rect 229710 149940 229738 150198
rect 230342 150204 230394 150210
rect 230952 150198 231026 150226
rect 231596 150198 231670 150226
rect 232240 150198 232314 150226
rect 232884 150198 232958 150226
rect 233252 150210 233280 159394
rect 233344 155310 233372 163200
rect 233516 157140 233568 157146
rect 233516 157082 233568 157088
rect 233332 155304 233384 155310
rect 233332 155246 233384 155252
rect 233528 150226 233556 157082
rect 234172 152590 234200 163200
rect 235000 159458 235028 163200
rect 234988 159452 235040 159458
rect 234988 159394 235040 159400
rect 234804 157072 234856 157078
rect 234804 157014 234856 157020
rect 234160 152584 234212 152590
rect 234160 152526 234212 152532
rect 234816 150226 234844 157014
rect 235092 153678 235120 163254
rect 235828 163146 235856 163254
rect 235906 163200 235962 164400
rect 236734 163200 236790 164400
rect 237562 163200 237618 164400
rect 238390 163200 238446 164400
rect 238864 163254 239168 163282
rect 235920 163146 235948 163200
rect 235828 163118 235948 163146
rect 236748 158030 236776 163200
rect 237576 158982 237604 163200
rect 237564 158976 237616 158982
rect 237564 158918 237616 158924
rect 238404 158846 238432 163200
rect 238392 158840 238444 158846
rect 238392 158782 238444 158788
rect 237380 158160 237432 158166
rect 237380 158102 237432 158108
rect 236736 158024 236788 158030
rect 236736 157966 236788 157972
rect 236092 157684 236144 157690
rect 236092 157626 236144 157632
rect 235448 153876 235500 153882
rect 235448 153818 235500 153824
rect 235080 153672 235132 153678
rect 235080 153614 235132 153620
rect 235460 150226 235488 153818
rect 236104 150226 236132 157626
rect 236736 152652 236788 152658
rect 236736 152594 236788 152600
rect 236748 150226 236776 152594
rect 237392 150226 237420 158102
rect 238024 154760 238076 154766
rect 238024 154702 238076 154708
rect 238036 150226 238064 154702
rect 238864 153610 238892 163254
rect 239140 163146 239168 163254
rect 239218 163200 239274 164400
rect 240046 163200 240102 164400
rect 240874 163200 240930 164400
rect 241794 163200 241850 164400
rect 241900 163254 242572 163282
rect 239232 163146 239260 163200
rect 239140 163118 239260 163146
rect 239312 159588 239364 159594
rect 239312 159530 239364 159536
rect 238944 158228 238996 158234
rect 238944 158170 238996 158176
rect 238668 153604 238720 153610
rect 238668 153546 238720 153552
rect 238852 153604 238904 153610
rect 238852 153546 238904 153552
rect 238680 150226 238708 153546
rect 230342 150146 230394 150152
rect 230354 149940 230382 150146
rect 230998 149940 231026 150198
rect 231642 149940 231670 150198
rect 232286 149940 232314 150198
rect 232930 149940 232958 150198
rect 233240 150204 233292 150210
rect 233528 150198 233602 150226
rect 233240 150146 233292 150152
rect 233574 149940 233602 150198
rect 234206 150204 234258 150210
rect 234816 150198 234890 150226
rect 235460 150198 235534 150226
rect 236104 150198 236178 150226
rect 236748 150198 236822 150226
rect 237392 150198 237466 150226
rect 238036 150198 238110 150226
rect 238680 150198 238754 150226
rect 238956 150210 238984 158170
rect 239324 150226 239352 159530
rect 240060 155242 240088 163200
rect 240232 159656 240284 159662
rect 240232 159598 240284 159604
rect 240048 155236 240100 155242
rect 240048 155178 240100 155184
rect 240244 152726 240272 159598
rect 240888 158778 240916 163200
rect 241808 158914 241836 163200
rect 241796 158908 241848 158914
rect 241796 158850 241848 158856
rect 241612 158840 241664 158846
rect 241612 158782 241664 158788
rect 240876 158772 240928 158778
rect 240876 158714 240928 158720
rect 240600 154692 240652 154698
rect 240600 154634 240652 154640
rect 240232 152720 240284 152726
rect 240232 152662 240284 152668
rect 240612 150226 240640 154634
rect 241244 154080 241296 154086
rect 241244 154022 241296 154028
rect 241256 150226 241284 154022
rect 241624 151910 241652 158782
rect 241900 153882 241928 163254
rect 242544 163146 242572 163254
rect 242622 163200 242678 164400
rect 243450 163200 243506 164400
rect 244278 163200 244334 164400
rect 244476 163254 245056 163282
rect 242636 163146 242664 163200
rect 242544 163118 242664 163146
rect 243360 158772 243412 158778
rect 243360 158714 243412 158720
rect 242072 158296 242124 158302
rect 242072 158238 242124 158244
rect 241888 153876 241940 153882
rect 241888 153818 241940 153824
rect 241888 152720 241940 152726
rect 241888 152662 241940 152668
rect 241612 151904 241664 151910
rect 241612 151846 241664 151852
rect 241900 150226 241928 152662
rect 242084 151814 242112 158238
rect 243084 154624 243136 154630
rect 243084 154566 243136 154572
rect 242084 151786 242480 151814
rect 242452 150226 242480 151786
rect 243096 150226 243124 154566
rect 243372 151978 243400 158714
rect 243464 158098 243492 163200
rect 244292 159662 244320 163200
rect 244280 159656 244332 159662
rect 244280 159598 244332 159604
rect 243452 158092 243504 158098
rect 243452 158034 243504 158040
rect 243728 153400 243780 153406
rect 243728 153342 243780 153348
rect 243360 151972 243412 151978
rect 243360 151914 243412 151920
rect 243740 150226 243768 153342
rect 244372 152788 244424 152794
rect 244372 152730 244424 152736
rect 244384 150226 244412 152730
rect 244476 152182 244504 163254
rect 245028 163146 245056 163254
rect 245106 163200 245162 164400
rect 245934 163200 245990 164400
rect 246762 163200 246818 164400
rect 247052 163254 247632 163282
rect 245120 163146 245148 163200
rect 245028 163118 245148 163146
rect 245016 158364 245068 158370
rect 245016 158306 245068 158312
rect 244464 152176 244516 152182
rect 244464 152118 244516 152124
rect 245028 150226 245056 158306
rect 245844 154896 245896 154902
rect 245844 154838 245896 154844
rect 245660 154148 245712 154154
rect 245660 154090 245712 154096
rect 245672 150226 245700 154090
rect 245856 151814 245884 154838
rect 245948 154154 245976 163200
rect 246776 158166 246804 163200
rect 246948 159724 247000 159730
rect 246948 159666 247000 159672
rect 246764 158160 246816 158166
rect 246764 158102 246816 158108
rect 245936 154148 245988 154154
rect 245936 154090 245988 154096
rect 245856 151786 246344 151814
rect 246316 150226 246344 151786
rect 246960 150226 246988 159666
rect 247052 152658 247080 163254
rect 247604 163146 247632 163254
rect 247682 163200 247738 164400
rect 248510 163200 248566 164400
rect 248616 163254 249288 163282
rect 247696 163146 247724 163200
rect 247604 163118 247724 163146
rect 248524 159730 248552 163200
rect 248512 159724 248564 159730
rect 248512 159666 248564 159672
rect 247132 158432 247184 158438
rect 247132 158374 247184 158380
rect 247040 152652 247092 152658
rect 247040 152594 247092 152600
rect 247144 151814 247172 158374
rect 248236 155508 248288 155514
rect 248236 155450 248288 155456
rect 247144 151786 247632 151814
rect 247604 150226 247632 151786
rect 248248 150226 248276 155450
rect 248616 154086 248644 163254
rect 249260 163146 249288 163254
rect 249338 163200 249394 164400
rect 250166 163200 250222 164400
rect 250994 163200 251050 164400
rect 251192 163254 251772 163282
rect 249352 163146 249380 163200
rect 249260 163118 249380 163146
rect 250076 158636 250128 158642
rect 250076 158578 250128 158584
rect 248604 154080 248656 154086
rect 248604 154022 248656 154028
rect 248880 153536 248932 153542
rect 248880 153478 248932 153484
rect 248892 150226 248920 153478
rect 249524 152448 249576 152454
rect 249524 152390 249576 152396
rect 249536 150226 249564 152390
rect 250088 151814 250116 158578
rect 250180 155378 250208 163200
rect 251008 159594 251036 163200
rect 250996 159588 251048 159594
rect 250996 159530 251048 159536
rect 250168 155372 250220 155378
rect 250168 155314 250220 155320
rect 250812 154216 250864 154222
rect 250812 154158 250864 154164
rect 250088 151786 250208 151814
rect 250180 150226 250208 151786
rect 250824 150226 250852 154158
rect 251192 152726 251220 163254
rect 251744 163146 251772 163254
rect 251822 163200 251878 164400
rect 252650 163200 252706 164400
rect 253570 163200 253626 164400
rect 254398 163200 254454 164400
rect 255226 163200 255282 164400
rect 255332 163254 256004 163282
rect 251836 163146 251864 163200
rect 251744 163118 251864 163146
rect 251456 157616 251508 157622
rect 251456 157558 251508 157564
rect 251180 152720 251232 152726
rect 251180 152662 251232 152668
rect 251468 150226 251496 157558
rect 252664 153542 252692 163200
rect 252744 158568 252796 158574
rect 252744 158510 252796 158516
rect 252652 153536 252704 153542
rect 252652 153478 252704 153484
rect 252100 152856 252152 152862
rect 252100 152798 252152 152804
rect 252112 150226 252140 152798
rect 252756 150226 252784 158510
rect 253388 155644 253440 155650
rect 253388 155586 253440 155592
rect 253400 150226 253428 155586
rect 253584 155446 253612 163200
rect 253940 159792 253992 159798
rect 253940 159734 253992 159740
rect 253572 155440 253624 155446
rect 253572 155382 253624 155388
rect 234206 150146 234258 150152
rect 234218 149940 234246 150146
rect 234862 149940 234890 150198
rect 235506 149940 235534 150198
rect 236150 149940 236178 150198
rect 236794 149940 236822 150198
rect 237438 149940 237466 150198
rect 238082 149940 238110 150198
rect 238726 149940 238754 150198
rect 238944 150204 238996 150210
rect 239324 150198 239398 150226
rect 238944 150146 238996 150152
rect 239370 149940 239398 150198
rect 240002 150204 240054 150210
rect 240612 150198 240686 150226
rect 241256 150198 241330 150226
rect 241900 150198 241974 150226
rect 242452 150198 242526 150226
rect 243096 150198 243170 150226
rect 243740 150198 243814 150226
rect 244384 150198 244458 150226
rect 245028 150198 245102 150226
rect 245672 150198 245746 150226
rect 246316 150198 246390 150226
rect 246960 150198 247034 150226
rect 247604 150198 247678 150226
rect 248248 150198 248322 150226
rect 248892 150198 248966 150226
rect 249536 150198 249610 150226
rect 250180 150198 250254 150226
rect 250824 150198 250898 150226
rect 251468 150198 251542 150226
rect 252112 150198 252186 150226
rect 252756 150198 252830 150226
rect 253400 150198 253474 150226
rect 253952 150210 253980 159734
rect 254412 158778 254440 163200
rect 255240 159798 255268 163200
rect 255228 159792 255280 159798
rect 255228 159734 255280 159740
rect 254400 158772 254452 158778
rect 254400 158714 254452 158720
rect 254032 157208 254084 157214
rect 254032 157150 254084 157156
rect 254044 150226 254072 157150
rect 255332 154222 255360 163254
rect 255976 163146 256004 163254
rect 256054 163200 256110 164400
rect 256882 163200 256938 164400
rect 257710 163200 257766 164400
rect 258538 163200 258594 164400
rect 259458 163200 259514 164400
rect 260286 163200 260342 164400
rect 261114 163200 261170 164400
rect 261942 163200 261998 164400
rect 262232 163254 262720 163282
rect 256068 163146 256096 163200
rect 255976 163118 256096 163146
rect 255412 158772 255464 158778
rect 255412 158714 255464 158720
rect 255320 154216 255372 154222
rect 255320 154158 255372 154164
rect 255424 152862 255452 158714
rect 256792 158704 256844 158710
rect 256792 158646 256844 158652
rect 255596 158500 255648 158506
rect 255596 158442 255648 158448
rect 255412 152856 255464 152862
rect 255412 152798 255464 152804
rect 255608 152538 255636 158442
rect 255872 157548 255924 157554
rect 255872 157490 255924 157496
rect 255688 155576 255740 155582
rect 255688 155518 255740 155524
rect 255424 152510 255636 152538
rect 255424 150226 255452 152510
rect 255700 151814 255728 155518
rect 255884 151814 255912 157490
rect 255700 151786 255820 151814
rect 255884 151786 256648 151814
rect 240002 150146 240054 150152
rect 240014 149940 240042 150146
rect 240658 149940 240686 150198
rect 241302 149940 241330 150198
rect 241946 149940 241974 150198
rect 242498 149940 242526 150198
rect 243142 149940 243170 150198
rect 243786 149940 243814 150198
rect 244430 149940 244458 150198
rect 245074 149940 245102 150198
rect 245718 149940 245746 150198
rect 246362 149940 246390 150198
rect 247006 149940 247034 150198
rect 247650 149940 247678 150198
rect 248294 149940 248322 150198
rect 248938 149940 248966 150198
rect 249582 149940 249610 150198
rect 250226 149940 250254 150198
rect 250870 149940 250898 150198
rect 251514 149940 251542 150198
rect 252158 149940 252186 150198
rect 252802 149940 252830 150198
rect 253446 149940 253474 150198
rect 253940 150204 253992 150210
rect 254044 150198 254118 150226
rect 253940 150146 253992 150152
rect 254090 149940 254118 150198
rect 254722 150204 254774 150210
rect 254722 150146 254774 150152
rect 255378 150198 255452 150226
rect 255792 150226 255820 151786
rect 256620 150226 256648 151786
rect 255792 150198 256050 150226
rect 256620 150198 256694 150226
rect 256804 150210 256832 158646
rect 256896 158234 256924 163200
rect 256884 158228 256936 158234
rect 256884 158170 256936 158176
rect 257252 153128 257304 153134
rect 257252 153070 257304 153076
rect 257264 150226 257292 153070
rect 257724 152794 257752 163200
rect 258552 158778 258580 163200
rect 258540 158772 258592 158778
rect 258540 158714 258592 158720
rect 258540 154284 258592 154290
rect 258540 154226 258592 154232
rect 257712 152788 257764 152794
rect 257712 152730 257764 152736
rect 258552 150226 258580 154226
rect 259184 153468 259236 153474
rect 259184 153410 259236 153416
rect 259196 150226 259224 153410
rect 259472 153406 259500 163200
rect 259552 159860 259604 159866
rect 259552 159802 259604 159808
rect 259460 153400 259512 153406
rect 259460 153342 259512 153348
rect 259564 151814 259592 159802
rect 260300 155514 260328 163200
rect 261128 158846 261156 163200
rect 261956 159866 261984 163200
rect 261944 159860 261996 159866
rect 261944 159802 261996 159808
rect 261116 158840 261168 158846
rect 261116 158782 261168 158788
rect 260932 158772 260984 158778
rect 260932 158714 260984 158720
rect 260472 157956 260524 157962
rect 260472 157898 260524 157904
rect 260288 155508 260340 155514
rect 260288 155450 260340 155456
rect 259564 151786 259868 151814
rect 259840 150226 259868 151786
rect 260484 150226 260512 157898
rect 260840 155712 260892 155718
rect 260840 155654 260892 155660
rect 260852 151814 260880 155654
rect 260944 152454 260972 158714
rect 261392 154964 261444 154970
rect 261392 154906 261444 154912
rect 260932 152448 260984 152454
rect 260932 152390 260984 152396
rect 261404 151814 261432 154906
rect 262232 154290 262260 163254
rect 262692 163146 262720 163254
rect 262770 163200 262826 164400
rect 263598 163200 263654 164400
rect 264426 163200 264482 164400
rect 264992 163254 265296 163282
rect 262784 163146 262812 163200
rect 262692 163118 262812 163146
rect 263048 157888 263100 157894
rect 263048 157830 263100 157836
rect 262220 154284 262272 154290
rect 262220 154226 262272 154232
rect 262404 152312 262456 152318
rect 262404 152254 262456 152260
rect 260852 151786 261156 151814
rect 261404 151786 261800 151814
rect 261128 150226 261156 151786
rect 261772 150226 261800 151786
rect 262416 150226 262444 152254
rect 263060 150226 263088 157830
rect 263612 155582 263640 163200
rect 264440 158778 264468 163200
rect 264888 159928 264940 159934
rect 264888 159870 264940 159876
rect 264428 158772 264480 158778
rect 264428 158714 264480 158720
rect 263692 157752 263744 157758
rect 263692 157694 263744 157700
rect 263600 155576 263652 155582
rect 263600 155518 263652 155524
rect 263704 150346 263732 157694
rect 263784 155848 263836 155854
rect 263784 155790 263836 155796
rect 263692 150340 263744 150346
rect 263692 150282 263744 150288
rect 263796 150226 263824 155790
rect 264900 151814 264928 159870
rect 264992 153134 265020 163254
rect 265268 163146 265296 163254
rect 265346 163200 265402 164400
rect 265452 163254 266124 163282
rect 265360 163146 265388 163200
rect 265268 163118 265388 163146
rect 265164 157276 265216 157282
rect 265164 157218 265216 157224
rect 264980 153128 265032 153134
rect 264980 153070 265032 153076
rect 265176 151814 265204 157218
rect 265452 153474 265480 163254
rect 266096 163146 266124 163254
rect 266174 163200 266230 164400
rect 267002 163200 267058 164400
rect 267830 163200 267886 164400
rect 268658 163200 268714 164400
rect 269224 163254 269436 163282
rect 266188 163146 266216 163200
rect 266096 163118 266216 163146
rect 266360 158772 266412 158778
rect 266360 158714 266412 158720
rect 266268 155916 266320 155922
rect 266268 155858 266320 155864
rect 265440 153468 265492 153474
rect 265440 153410 265492 153416
rect 264900 151786 265020 151814
rect 265176 151786 265664 151814
rect 254734 149940 254762 150146
rect 255378 149940 255406 150198
rect 256022 149940 256050 150198
rect 256666 149940 256694 150198
rect 256792 150204 256844 150210
rect 257264 150198 257338 150226
rect 256792 150146 256844 150152
rect 257310 149940 257338 150198
rect 257942 150204 257994 150210
rect 258552 150198 258626 150226
rect 259196 150198 259270 150226
rect 259840 150198 259914 150226
rect 260484 150198 260558 150226
rect 261128 150198 261202 150226
rect 261772 150198 261846 150226
rect 262416 150198 262490 150226
rect 263060 150198 263134 150226
rect 257942 150146 257994 150152
rect 257954 149940 257982 150146
rect 258598 149940 258626 150198
rect 259242 149940 259270 150198
rect 259886 149940 259914 150198
rect 260530 149940 260558 150198
rect 261174 149940 261202 150198
rect 261818 149940 261846 150198
rect 262462 149940 262490 150198
rect 263106 149940 263134 150198
rect 263750 150198 263824 150226
rect 264992 150226 265020 151786
rect 265636 150226 265664 151786
rect 266280 150226 266308 155858
rect 266372 152318 266400 158714
rect 266912 156256 266964 156262
rect 266912 156198 266964 156204
rect 266360 152312 266412 152318
rect 266360 152254 266412 152260
rect 266924 150226 266952 156198
rect 267016 155650 267044 163200
rect 267844 158778 267872 163200
rect 268672 159934 268700 163200
rect 269120 159996 269172 160002
rect 269120 159938 269172 159944
rect 268660 159928 268712 159934
rect 268660 159870 268712 159876
rect 267832 158772 267884 158778
rect 267832 158714 267884 158720
rect 267740 157820 267792 157826
rect 267740 157762 267792 157768
rect 267004 155644 267056 155650
rect 267004 155586 267056 155592
rect 267556 153060 267608 153066
rect 267556 153002 267608 153008
rect 267568 150226 267596 153002
rect 267752 151814 267780 157762
rect 268844 155168 268896 155174
rect 268844 155110 268896 155116
rect 267752 151786 268240 151814
rect 268212 150226 268240 151786
rect 268856 150226 268884 155110
rect 264382 150204 264434 150210
rect 263750 149940 263778 150198
rect 264992 150198 265066 150226
rect 265636 150198 265710 150226
rect 266280 150198 266354 150226
rect 266924 150198 266998 150226
rect 267568 150198 267642 150226
rect 268212 150198 268286 150226
rect 268856 150198 268930 150226
rect 269132 150210 269160 159938
rect 269224 153338 269252 163254
rect 269408 163146 269436 163254
rect 269486 163200 269542 164400
rect 270314 163200 270370 164400
rect 271234 163200 271290 164400
rect 272062 163200 272118 164400
rect 272890 163200 272946 164400
rect 273718 163200 273774 164400
rect 274546 163200 274602 164400
rect 275374 163200 275430 164400
rect 276202 163200 276258 164400
rect 277122 163200 277178 164400
rect 277412 163254 277900 163282
rect 269500 163146 269528 163200
rect 269408 163118 269528 163146
rect 270328 155718 270356 163200
rect 271248 160002 271276 163200
rect 272076 161474 272104 163200
rect 272076 161446 272196 161474
rect 271236 159996 271288 160002
rect 271236 159938 271288 159944
rect 272064 156936 272116 156942
rect 272064 156878 272116 156884
rect 270500 156596 270552 156602
rect 270500 156538 270552 156544
rect 270316 155712 270368 155718
rect 270316 155654 270368 155660
rect 269488 155032 269540 155038
rect 269488 154974 269540 154980
rect 269212 153332 269264 153338
rect 269212 153274 269264 153280
rect 269500 150226 269528 154974
rect 270512 151814 270540 156538
rect 271420 155100 271472 155106
rect 271420 155042 271472 155048
rect 270512 151786 270816 151814
rect 270788 150226 270816 151786
rect 271432 150226 271460 155042
rect 272076 150226 272104 156878
rect 272168 153066 272196 161446
rect 272800 159996 272852 160002
rect 272800 159938 272852 159944
rect 272156 153060 272208 153066
rect 272156 153002 272208 153008
rect 272812 152046 272840 159938
rect 272904 153270 272932 163200
rect 273732 157010 273760 163200
rect 274560 159497 274588 163200
rect 275388 160002 275416 163200
rect 275376 159996 275428 160002
rect 275376 159938 275428 159944
rect 274546 159488 274602 159497
rect 274546 159423 274602 159432
rect 275190 159352 275246 159361
rect 275190 159287 275246 159296
rect 273720 157004 273772 157010
rect 273720 156946 273772 156952
rect 273904 156120 273956 156126
rect 273904 156062 273956 156068
rect 273260 156052 273312 156058
rect 273260 155994 273312 156000
rect 272892 153264 272944 153270
rect 272892 153206 272944 153212
rect 272708 152040 272760 152046
rect 272708 151982 272760 151988
rect 272800 152040 272852 152046
rect 272800 151982 272852 151988
rect 272720 150226 272748 151982
rect 264382 150146 264434 150152
rect 264394 149940 264422 150146
rect 265038 149940 265066 150198
rect 265682 149940 265710 150198
rect 266326 149940 266354 150198
rect 266970 149940 266998 150198
rect 267614 149940 267642 150198
rect 268258 149940 268286 150198
rect 268902 149940 268930 150198
rect 269120 150204 269172 150210
rect 269500 150198 269574 150226
rect 269120 150146 269172 150152
rect 269546 149940 269574 150198
rect 270178 150204 270230 150210
rect 270788 150198 270862 150226
rect 271432 150198 271506 150226
rect 272076 150198 272150 150226
rect 272720 150198 272794 150226
rect 270178 150146 270230 150152
rect 270190 149940 270218 150146
rect 270834 149940 270862 150198
rect 271478 149940 271506 150198
rect 272122 149940 272150 150198
rect 272766 149940 272794 150198
rect 273272 150090 273300 155994
rect 273916 150090 273944 156062
rect 274548 152108 274600 152114
rect 274548 152050 274600 152056
rect 274560 150090 274588 152050
rect 275204 150226 275232 159287
rect 275468 154828 275520 154834
rect 275468 154770 275520 154776
rect 275480 154698 275508 154770
rect 275468 154692 275520 154698
rect 275468 154634 275520 154640
rect 276216 154426 276244 163200
rect 277136 156942 277164 163200
rect 277124 156936 277176 156942
rect 277124 156878 277176 156884
rect 277124 156188 277176 156194
rect 277124 156130 277176 156136
rect 276480 155780 276532 155786
rect 276480 155722 276532 155728
rect 275284 154420 275336 154426
rect 275284 154362 275336 154368
rect 276204 154420 276256 154426
rect 276204 154362 276256 154368
rect 275296 150362 275324 154362
rect 275296 150334 275876 150362
rect 275848 150226 275876 150334
rect 275204 150198 275278 150226
rect 275848 150198 275922 150226
rect 273272 150062 273346 150090
rect 273916 150062 273990 150090
rect 274560 150062 274634 150090
rect 273318 149940 273346 150062
rect 273962 149940 273990 150062
rect 274606 149940 274634 150062
rect 275250 149940 275278 150198
rect 275894 149940 275922 150198
rect 276492 150090 276520 155722
rect 277136 150090 277164 156130
rect 277412 152114 277440 163254
rect 277872 163146 277900 163254
rect 277950 163200 278006 164400
rect 278778 163200 278834 164400
rect 278884 163254 279556 163282
rect 277964 163146 277992 163200
rect 277872 163118 277992 163146
rect 278412 154352 278464 154358
rect 278412 154294 278464 154300
rect 277768 152924 277820 152930
rect 277768 152866 277820 152872
rect 277400 152108 277452 152114
rect 277400 152050 277452 152056
rect 277780 150090 277808 152866
rect 278424 150090 278452 154294
rect 278792 152930 278820 163200
rect 278884 154358 278912 163254
rect 279528 163146 279556 163254
rect 279606 163200 279662 164400
rect 280434 163200 280490 164400
rect 281262 163200 281318 164400
rect 282090 163200 282146 164400
rect 283010 163200 283066 164400
rect 283838 163200 283894 164400
rect 284666 163200 284722 164400
rect 285494 163200 285550 164400
rect 285692 163254 286272 163282
rect 279620 163146 279648 163200
rect 279528 163118 279648 163146
rect 280344 160064 280396 160070
rect 280344 160006 280396 160012
rect 279056 156392 279108 156398
rect 279056 156334 279108 156340
rect 278872 154352 278924 154358
rect 278872 154294 278924 154300
rect 278780 152924 278832 152930
rect 278780 152866 278832 152872
rect 279068 150090 279096 156334
rect 279700 153196 279752 153202
rect 279700 153138 279752 153144
rect 279712 150090 279740 153138
rect 280356 150226 280384 160006
rect 280448 157078 280476 163200
rect 281276 160070 281304 163200
rect 281264 160064 281316 160070
rect 281264 160006 281316 160012
rect 282104 159322 282132 163200
rect 281540 159316 281592 159322
rect 281540 159258 281592 159264
rect 282092 159316 282144 159322
rect 282092 159258 282144 159264
rect 281552 157334 281580 159258
rect 281552 157306 282316 157334
rect 281632 157208 281684 157214
rect 281632 157150 281684 157156
rect 280436 157072 280488 157078
rect 280436 157014 280488 157020
rect 280986 153776 281042 153785
rect 280986 153711 281042 153720
rect 280356 150198 280430 150226
rect 276492 150062 276566 150090
rect 277136 150062 277210 150090
rect 277780 150062 277854 150090
rect 278424 150062 278498 150090
rect 279068 150062 279142 150090
rect 279712 150062 279786 150090
rect 276538 149940 276566 150062
rect 277182 149940 277210 150062
rect 277826 149940 277854 150062
rect 278470 149940 278498 150062
rect 279114 149940 279142 150062
rect 279758 149940 279786 150062
rect 280402 149940 280430 150198
rect 281000 150090 281028 153711
rect 281644 150090 281672 157150
rect 282288 150226 282316 157306
rect 283024 154562 283052 163200
rect 283196 159112 283248 159118
rect 283196 159054 283248 159060
rect 283104 156664 283156 156670
rect 283104 156606 283156 156612
rect 283012 154556 283064 154562
rect 283012 154498 283064 154504
rect 282920 152244 282972 152250
rect 282920 152186 282972 152192
rect 282932 150226 282960 152186
rect 282288 150198 282362 150226
rect 282932 150198 283006 150226
rect 283116 150210 283144 156606
rect 283208 151842 283236 159054
rect 283852 157282 283880 163200
rect 284392 159248 284444 159254
rect 284392 159190 284444 159196
rect 283840 157276 283892 157282
rect 283840 157218 283892 157224
rect 283760 154562 283972 154578
rect 283748 154556 283984 154562
rect 283800 154550 283932 154556
rect 283748 154498 283800 154504
rect 283932 154498 283984 154504
rect 283656 154488 283708 154494
rect 283656 154430 283708 154436
rect 283196 151836 283248 151842
rect 283196 151778 283248 151784
rect 283668 150226 283696 154430
rect 281000 150062 281074 150090
rect 281644 150062 281718 150090
rect 281046 149940 281074 150062
rect 281690 149940 281718 150062
rect 282334 149940 282362 150198
rect 282978 149940 283006 150198
rect 283104 150204 283156 150210
rect 283104 150146 283156 150152
rect 283622 150198 283696 150226
rect 284404 150210 284432 159190
rect 284680 159118 284708 163200
rect 284668 159112 284720 159118
rect 284668 159054 284720 159060
rect 285508 153202 285536 163200
rect 285692 154494 285720 163254
rect 286244 163146 286272 163254
rect 286322 163200 286378 164400
rect 287150 163200 287206 164400
rect 287978 163200 288034 164400
rect 288898 163200 288954 164400
rect 289726 163200 289782 164400
rect 290554 163200 290610 164400
rect 291382 163200 291438 164400
rect 292210 163200 292266 164400
rect 293038 163200 293094 164400
rect 293866 163200 293922 164400
rect 294786 163200 294842 164400
rect 295614 163200 295670 164400
rect 296442 163200 296498 164400
rect 297270 163200 297326 164400
rect 298098 163200 298154 164400
rect 298664 163254 298876 163282
rect 286336 163146 286364 163200
rect 286244 163118 286364 163146
rect 285772 159112 285824 159118
rect 285772 159054 285824 159060
rect 285588 154488 285640 154494
rect 285588 154430 285640 154436
rect 285680 154488 285732 154494
rect 285680 154430 285732 154436
rect 285600 154306 285628 154430
rect 285600 154278 285720 154306
rect 285496 153196 285548 153202
rect 285496 153138 285548 153144
rect 284852 152992 284904 152998
rect 284852 152934 284904 152940
rect 284864 150226 284892 152934
rect 285692 151814 285720 154278
rect 285784 152250 285812 159054
rect 287164 157146 287192 163200
rect 287992 159254 288020 163200
rect 287980 159248 288032 159254
rect 287980 159190 288032 159196
rect 288912 159118 288940 163200
rect 288072 159112 288124 159118
rect 288072 159054 288124 159060
rect 288900 159112 288952 159118
rect 288900 159054 288952 159060
rect 287152 157140 287204 157146
rect 287152 157082 287204 157088
rect 286232 156324 286284 156330
rect 286232 156266 286284 156272
rect 285772 152244 285824 152250
rect 285772 152186 285824 152192
rect 286244 151814 286272 156266
rect 288084 152998 288112 159054
rect 289360 156732 289412 156738
rect 289360 156674 289412 156680
rect 288716 154012 288768 154018
rect 288716 153954 288768 153960
rect 288072 152992 288124 152998
rect 288072 152934 288124 152940
rect 288072 152380 288124 152386
rect 288072 152322 288124 152328
rect 287428 151836 287480 151842
rect 285692 151786 286180 151814
rect 286244 151786 286824 151814
rect 286152 150226 286180 151786
rect 286796 150226 286824 151786
rect 287428 151778 287480 151784
rect 287440 150226 287468 151778
rect 288084 150226 288112 152322
rect 288728 150226 288756 153954
rect 289372 150226 289400 156674
rect 289740 155786 289768 163200
rect 290568 156738 290596 163200
rect 290648 159180 290700 159186
rect 290648 159122 290700 159128
rect 290556 156732 290608 156738
rect 290556 156674 290608 156680
rect 289728 155780 289780 155786
rect 289728 155722 289780 155728
rect 290004 152992 290056 152998
rect 290004 152934 290056 152940
rect 290016 150226 290044 152934
rect 290660 150226 290688 159122
rect 291292 153944 291344 153950
rect 291292 153886 291344 153892
rect 291304 150226 291332 153886
rect 291396 152998 291424 163200
rect 291936 156868 291988 156874
rect 291936 156810 291988 156816
rect 291384 152992 291436 152998
rect 291384 152934 291436 152940
rect 291948 150226 291976 156810
rect 292224 152386 292252 163200
rect 293052 155854 293080 163200
rect 293880 156874 293908 163200
rect 294800 159526 294828 163200
rect 293960 159520 294012 159526
rect 293960 159462 294012 159468
rect 294788 159520 294840 159526
rect 294788 159462 294840 159468
rect 293972 159186 294000 159462
rect 295628 159390 295656 163200
rect 295524 159384 295576 159390
rect 295524 159326 295576 159332
rect 295616 159384 295668 159390
rect 295616 159326 295668 159332
rect 293960 159180 294012 159186
rect 293960 159122 294012 159128
rect 295156 159180 295208 159186
rect 295156 159122 295208 159128
rect 293868 156868 293920 156874
rect 293868 156810 293920 156816
rect 294052 156800 294104 156806
rect 294052 156742 294104 156748
rect 293040 155848 293092 155854
rect 293040 155790 293092 155796
rect 293868 153740 293920 153746
rect 293868 153682 293920 153688
rect 293224 152516 293276 152522
rect 293224 152458 293276 152464
rect 292578 152416 292634 152425
rect 292212 152380 292264 152386
rect 292578 152351 292634 152360
rect 292212 152322 292264 152328
rect 292592 150226 292620 152351
rect 293236 150226 293264 152458
rect 293880 150226 293908 153682
rect 294064 151814 294092 156742
rect 294064 151786 294552 151814
rect 294524 150226 294552 151786
rect 295168 150226 295196 159122
rect 295536 151814 295564 159326
rect 296456 155922 296484 163200
rect 297284 156806 297312 163200
rect 298008 159452 298060 159458
rect 298008 159394 298060 159400
rect 297272 156800 297324 156806
rect 297272 156742 297324 156748
rect 296444 155916 296496 155922
rect 296444 155858 296496 155864
rect 297088 155304 297140 155310
rect 297088 155246 297140 155252
rect 296444 153808 296496 153814
rect 296444 153750 296496 153756
rect 295536 151786 295840 151814
rect 295812 150226 295840 151786
rect 296456 150226 296484 153750
rect 297100 150226 297128 155246
rect 297732 152584 297784 152590
rect 297732 152526 297784 152532
rect 297744 150226 297772 152526
rect 298020 151814 298048 159394
rect 298112 159050 298140 163200
rect 298100 159044 298152 159050
rect 298100 158986 298152 158992
rect 298664 152522 298692 163254
rect 298848 163146 298876 163254
rect 298926 163200 298982 164400
rect 299754 163200 299810 164400
rect 300674 163200 300730 164400
rect 301502 163200 301558 164400
rect 302330 163200 302386 164400
rect 303158 163200 303214 164400
rect 303632 163254 303936 163282
rect 298940 163146 298968 163200
rect 298848 163118 298968 163146
rect 299480 158976 299532 158982
rect 299480 158918 299532 158924
rect 299020 153672 299072 153678
rect 299020 153614 299072 153620
rect 298652 152516 298704 152522
rect 298652 152458 298704 152464
rect 298020 151786 298416 151814
rect 298388 150226 298416 151786
rect 299032 150226 299060 153614
rect 284254 150204 284306 150210
rect 283622 149940 283650 150198
rect 284254 150146 284306 150152
rect 284392 150204 284444 150210
rect 284864 150198 284938 150226
rect 284392 150146 284444 150152
rect 284266 149940 284294 150146
rect 284910 149940 284938 150198
rect 285542 150204 285594 150210
rect 286152 150198 286226 150226
rect 286796 150198 286870 150226
rect 287440 150198 287514 150226
rect 288084 150198 288158 150226
rect 288728 150198 288802 150226
rect 289372 150198 289446 150226
rect 290016 150198 290090 150226
rect 290660 150198 290734 150226
rect 291304 150198 291378 150226
rect 291948 150198 292022 150226
rect 292592 150198 292666 150226
rect 293236 150198 293310 150226
rect 293880 150198 293954 150226
rect 294524 150198 294598 150226
rect 295168 150198 295242 150226
rect 295812 150198 295886 150226
rect 296456 150198 296530 150226
rect 297100 150198 297174 150226
rect 297744 150198 297818 150226
rect 298388 150198 298462 150226
rect 299032 150198 299106 150226
rect 299492 150210 299520 158918
rect 299664 158024 299716 158030
rect 299664 157966 299716 157972
rect 299676 150226 299704 157966
rect 299768 155310 299796 163200
rect 300400 159044 300452 159050
rect 300400 158986 300452 158992
rect 299756 155304 299808 155310
rect 299756 155246 299808 155252
rect 300412 151842 300440 158986
rect 300688 157214 300716 163200
rect 301516 159458 301544 163200
rect 301504 159452 301556 159458
rect 301504 159394 301556 159400
rect 302344 159186 302372 163200
rect 302332 159180 302384 159186
rect 302332 159122 302384 159128
rect 300676 157208 300728 157214
rect 300676 157150 300728 157156
rect 302516 155236 302568 155242
rect 302516 155178 302568 155184
rect 301596 153604 301648 153610
rect 301596 153546 301648 153552
rect 300952 151904 301004 151910
rect 300952 151846 301004 151852
rect 300400 151836 300452 151842
rect 300400 151778 300452 151784
rect 300964 150226 300992 151846
rect 301608 150226 301636 153546
rect 302528 151814 302556 155178
rect 303172 155106 303200 163200
rect 303528 158908 303580 158914
rect 303528 158850 303580 158856
rect 303160 155100 303212 155106
rect 303160 155042 303212 155048
rect 302884 151972 302936 151978
rect 302884 151914 302936 151920
rect 302344 151786 302556 151814
rect 302344 150226 302372 151786
rect 285542 150146 285594 150152
rect 285554 149940 285582 150146
rect 286198 149940 286226 150198
rect 286842 149940 286870 150198
rect 287486 149940 287514 150198
rect 288130 149940 288158 150198
rect 288774 149940 288802 150198
rect 289418 149940 289446 150198
rect 290062 149940 290090 150198
rect 290706 149940 290734 150198
rect 291350 149940 291378 150198
rect 291994 149940 292022 150198
rect 292638 149940 292666 150198
rect 293282 149940 293310 150198
rect 293926 149940 293954 150198
rect 294570 149940 294598 150198
rect 295214 149940 295242 150198
rect 295858 149940 295886 150198
rect 296502 149940 296530 150198
rect 297146 149940 297174 150198
rect 297790 149940 297818 150198
rect 298434 149940 298462 150198
rect 299078 149940 299106 150198
rect 299480 150204 299532 150210
rect 299676 150198 299750 150226
rect 299480 150146 299532 150152
rect 299722 149940 299750 150198
rect 300354 150204 300406 150210
rect 300964 150198 301038 150226
rect 301608 150198 301682 150226
rect 300354 150146 300406 150152
rect 300366 149940 300394 150146
rect 301010 149940 301038 150198
rect 301654 149940 301682 150198
rect 302298 150198 302372 150226
rect 302896 150226 302924 151914
rect 303540 150226 303568 158850
rect 303632 152590 303660 163254
rect 303908 163146 303936 163254
rect 303986 163200 304042 164400
rect 304184 163254 304764 163282
rect 304000 163146 304028 163200
rect 303908 163118 304028 163146
rect 304080 153876 304132 153882
rect 304080 153818 304132 153824
rect 303620 152584 303672 152590
rect 303620 152526 303672 152532
rect 304092 150226 304120 153818
rect 304184 151978 304212 163254
rect 304736 163146 304764 163254
rect 304814 163200 304870 164400
rect 305642 163200 305698 164400
rect 306562 163200 306618 164400
rect 307390 163200 307446 164400
rect 308218 163200 308274 164400
rect 309046 163200 309102 164400
rect 309152 163254 309824 163282
rect 304828 163146 304856 163200
rect 304736 163118 304856 163146
rect 305368 159656 305420 159662
rect 305368 159598 305420 159604
rect 304724 158092 304776 158098
rect 304724 158034 304776 158040
rect 304172 151972 304224 151978
rect 304172 151914 304224 151920
rect 304736 150226 304764 158034
rect 305380 150226 305408 159598
rect 305656 158914 305684 163200
rect 305644 158908 305696 158914
rect 305644 158850 305696 158856
rect 306576 155242 306604 163200
rect 307404 159050 307432 163200
rect 308232 159730 308260 163200
rect 308220 159724 308272 159730
rect 308220 159666 308272 159672
rect 309060 159662 309088 163200
rect 308588 159656 308640 159662
rect 308588 159598 308640 159604
rect 309048 159656 309100 159662
rect 309048 159598 309100 159604
rect 307392 159044 307444 159050
rect 307392 158986 307444 158992
rect 307392 158908 307444 158914
rect 307392 158850 307444 158856
rect 306932 158160 306984 158166
rect 306932 158102 306984 158108
rect 306564 155236 306616 155242
rect 306564 155178 306616 155184
rect 306656 154148 306708 154154
rect 306656 154090 306708 154096
rect 306012 152176 306064 152182
rect 306012 152118 306064 152124
rect 306024 150226 306052 152118
rect 306668 150226 306696 154090
rect 306944 151814 306972 158102
rect 307404 151910 307432 158850
rect 307944 152652 307996 152658
rect 307944 152594 307996 152600
rect 307392 151904 307444 151910
rect 307392 151846 307444 151852
rect 306944 151786 307340 151814
rect 307312 150226 307340 151786
rect 307956 150226 307984 152594
rect 308600 150226 308628 159598
rect 309152 153882 309180 163254
rect 309796 163146 309824 163254
rect 309874 163200 309930 164400
rect 310702 163200 310758 164400
rect 311530 163200 311586 164400
rect 312450 163200 312506 164400
rect 313278 163200 313334 164400
rect 314106 163200 314162 164400
rect 314934 163200 314990 164400
rect 315762 163200 315818 164400
rect 316052 163254 316540 163282
rect 309888 163146 309916 163200
rect 309796 163118 309916 163146
rect 310612 159588 310664 159594
rect 310612 159530 310664 159536
rect 309876 155372 309928 155378
rect 309876 155314 309928 155320
rect 309232 154080 309284 154086
rect 309232 154022 309284 154028
rect 309140 153876 309192 153882
rect 309140 153818 309192 153824
rect 309244 150226 309272 154022
rect 309888 150226 309916 155314
rect 310624 150226 310652 159530
rect 310716 158914 310744 163200
rect 310704 158908 310756 158914
rect 310704 158850 310756 158856
rect 311164 152720 311216 152726
rect 311164 152662 311216 152668
rect 302896 150198 302970 150226
rect 303540 150198 303614 150226
rect 304092 150198 304166 150226
rect 304736 150198 304810 150226
rect 305380 150198 305454 150226
rect 306024 150198 306098 150226
rect 306668 150198 306742 150226
rect 307312 150198 307386 150226
rect 307956 150198 308030 150226
rect 308600 150198 308674 150226
rect 309244 150198 309318 150226
rect 309888 150198 309962 150226
rect 302298 149940 302326 150198
rect 302942 149940 302970 150198
rect 303586 149940 303614 150198
rect 304138 149940 304166 150198
rect 304782 149940 304810 150198
rect 305426 149940 305454 150198
rect 306070 149940 306098 150198
rect 306714 149940 306742 150198
rect 307358 149940 307386 150198
rect 308002 149940 308030 150198
rect 308646 149940 308674 150198
rect 309290 149940 309318 150198
rect 309934 149940 309962 150198
rect 310578 150198 310652 150226
rect 311176 150226 311204 152662
rect 311544 152658 311572 163200
rect 312464 159866 312492 163200
rect 312360 159860 312412 159866
rect 312360 159802 312412 159808
rect 312452 159860 312504 159866
rect 312452 159802 312504 159808
rect 312372 158914 312400 159802
rect 312176 158908 312228 158914
rect 312176 158850 312228 158856
rect 312360 158908 312412 158914
rect 312360 158850 312412 158856
rect 311808 153536 311860 153542
rect 311808 153478 311860 153484
rect 311532 152652 311584 152658
rect 311532 152594 311584 152600
rect 311820 150226 311848 153478
rect 312188 152726 312216 158850
rect 312452 155440 312504 155446
rect 312452 155382 312504 155388
rect 312176 152720 312228 152726
rect 312176 152662 312228 152668
rect 312464 150226 312492 155382
rect 313292 154018 313320 163200
rect 313372 159860 313424 159866
rect 313372 159802 313424 159808
rect 313280 154012 313332 154018
rect 313280 153954 313332 153960
rect 313096 152856 313148 152862
rect 313096 152798 313148 152804
rect 313108 150226 313136 152798
rect 313384 152425 313412 159802
rect 314120 159798 314148 163200
rect 313464 159792 313516 159798
rect 313464 159734 313516 159740
rect 314108 159792 314160 159798
rect 314108 159734 314160 159740
rect 313370 152416 313426 152425
rect 313370 152351 313426 152360
rect 313476 151814 313504 159734
rect 314948 158982 314976 163200
rect 315776 159594 315804 163200
rect 315764 159588 315816 159594
rect 315764 159530 315816 159536
rect 314936 158976 314988 158982
rect 314936 158918 314988 158924
rect 315028 158228 315080 158234
rect 315028 158170 315080 158176
rect 314384 154216 314436 154222
rect 314384 154158 314436 154164
rect 313476 151786 313780 151814
rect 313752 150226 313780 151786
rect 314396 150226 314424 154158
rect 315040 150226 315068 158170
rect 316052 153950 316080 163254
rect 316512 163146 316540 163254
rect 316590 163200 316646 164400
rect 317418 163200 317474 164400
rect 317524 163254 318288 163282
rect 316604 163146 316632 163200
rect 316512 163118 316632 163146
rect 317052 158840 317104 158846
rect 317052 158782 317104 158788
rect 316040 153944 316092 153950
rect 316040 153886 316092 153892
rect 316960 153400 317012 153406
rect 316960 153342 317012 153348
rect 315672 152788 315724 152794
rect 315672 152730 315724 152736
rect 315684 150226 315712 152730
rect 316316 152448 316368 152454
rect 316316 152390 316368 152396
rect 316328 150226 316356 152390
rect 316972 150226 317000 153342
rect 317064 152862 317092 158782
rect 317052 152856 317104 152862
rect 317052 152798 317104 152804
rect 317432 152794 317460 163200
rect 317420 152788 317472 152794
rect 317420 152730 317472 152736
rect 317524 152454 317552 163254
rect 318260 163146 318288 163254
rect 318338 163200 318394 164400
rect 319166 163200 319222 164400
rect 319994 163200 320050 164400
rect 320822 163200 320878 164400
rect 321650 163200 321706 164400
rect 322478 163200 322534 164400
rect 323306 163200 323362 164400
rect 324226 163200 324282 164400
rect 324332 163254 325004 163282
rect 318352 163146 318380 163200
rect 318260 163118 318380 163146
rect 318892 158908 318944 158914
rect 318892 158850 318944 158856
rect 317604 155508 317656 155514
rect 317604 155450 317656 155456
rect 317512 152448 317564 152454
rect 317512 152390 317564 152396
rect 317616 150226 317644 155450
rect 318248 152856 318300 152862
rect 318248 152798 318300 152804
rect 318260 150226 318288 152798
rect 318904 150226 318932 158850
rect 319180 158846 319208 163200
rect 319168 158840 319220 158846
rect 319168 158782 319220 158788
rect 320008 155378 320036 163200
rect 320836 158914 320864 163200
rect 320824 158908 320876 158914
rect 320824 158850 320876 158856
rect 321664 158846 321692 163200
rect 322492 159866 322520 163200
rect 322480 159860 322532 159866
rect 322480 159802 322532 159808
rect 321652 158840 321704 158846
rect 321652 158782 321704 158788
rect 320272 158772 320324 158778
rect 320272 158714 320324 158720
rect 320180 155576 320232 155582
rect 320180 155518 320232 155524
rect 319996 155372 320048 155378
rect 319996 155314 320048 155320
rect 319536 154284 319588 154290
rect 319536 154226 319588 154232
rect 319548 150226 319576 154226
rect 320192 150226 320220 155518
rect 320284 152794 320312 158714
rect 321560 158704 321612 158710
rect 321560 158646 321612 158652
rect 321468 153128 321520 153134
rect 321468 153070 321520 153076
rect 320272 152788 320324 152794
rect 320272 152730 320324 152736
rect 320640 152652 320692 152658
rect 320640 152594 320692 152600
rect 320824 152652 320876 152658
rect 320824 152594 320876 152600
rect 320652 152182 320680 152594
rect 320836 152538 320864 152594
rect 320744 152510 320864 152538
rect 320744 152454 320772 152510
rect 320732 152448 320784 152454
rect 320732 152390 320784 152396
rect 320824 152448 320876 152454
rect 320824 152390 320876 152396
rect 320640 152176 320692 152182
rect 320640 152118 320692 152124
rect 320836 152046 320864 152390
rect 320916 152312 320968 152318
rect 320916 152254 320968 152260
rect 320824 152040 320876 152046
rect 320824 151982 320876 151988
rect 320928 150226 320956 152254
rect 311176 150198 311250 150226
rect 311820 150198 311894 150226
rect 312464 150198 312538 150226
rect 313108 150198 313182 150226
rect 313752 150198 313826 150226
rect 314396 150198 314470 150226
rect 315040 150198 315114 150226
rect 315684 150198 315758 150226
rect 316328 150198 316402 150226
rect 316972 150198 317046 150226
rect 317616 150198 317690 150226
rect 318260 150198 318334 150226
rect 318904 150198 318978 150226
rect 319548 150198 319622 150226
rect 320192 150198 320266 150226
rect 310578 149940 310606 150198
rect 311222 149940 311250 150198
rect 311866 149940 311894 150198
rect 312510 149940 312538 150198
rect 313154 149940 313182 150198
rect 313798 149940 313826 150198
rect 314442 149940 314470 150198
rect 315086 149940 315114 150198
rect 315730 149940 315758 150198
rect 316374 149940 316402 150198
rect 317018 149940 317046 150198
rect 317662 149940 317690 150198
rect 318306 149940 318334 150198
rect 318950 149940 318978 150198
rect 319594 149940 319622 150198
rect 320238 149940 320266 150198
rect 320882 150198 320956 150226
rect 321480 150226 321508 153070
rect 321572 152046 321600 158646
rect 322112 155644 322164 155650
rect 322112 155586 322164 155592
rect 322020 153468 322072 153474
rect 322020 153410 322072 153416
rect 321560 152040 321612 152046
rect 321560 151982 321612 151988
rect 322032 150498 322060 153410
rect 322124 151814 322152 155586
rect 323320 154086 323348 163200
rect 324044 159928 324096 159934
rect 324044 159870 324096 159876
rect 323308 154080 323360 154086
rect 323308 154022 323360 154028
rect 323124 152788 323176 152794
rect 323124 152730 323176 152736
rect 323136 151814 323164 152730
rect 322124 151786 322796 151814
rect 323136 151786 323440 151814
rect 322032 150470 322152 150498
rect 322124 150226 322152 150470
rect 322768 150226 322796 151786
rect 323412 150226 323440 151786
rect 324056 150226 324084 159870
rect 324240 152794 324268 163200
rect 324332 153134 324360 163254
rect 324976 163146 325004 163254
rect 325054 163200 325110 164400
rect 325882 163200 325938 164400
rect 326710 163200 326766 164400
rect 327538 163200 327594 164400
rect 328366 163200 328422 164400
rect 329194 163200 329250 164400
rect 330114 163200 330170 164400
rect 330942 163200 330998 164400
rect 331232 163254 331720 163282
rect 325068 163146 325096 163200
rect 324976 163118 325096 163146
rect 325896 157334 325924 163200
rect 325896 157306 326108 157334
rect 325332 155712 325384 155718
rect 325332 155654 325384 155660
rect 324688 153332 324740 153338
rect 324688 153274 324740 153280
rect 324320 153128 324372 153134
rect 324320 153070 324372 153076
rect 324228 152788 324280 152794
rect 324228 152730 324280 152736
rect 324700 150226 324728 153274
rect 325344 150226 325372 155654
rect 326080 152454 326108 157306
rect 326724 154154 326752 163200
rect 327552 158778 327580 163200
rect 328380 159934 328408 163200
rect 329208 160002 329236 163200
rect 328460 159996 328512 160002
rect 328460 159938 328512 159944
rect 329196 159996 329248 160002
rect 329196 159938 329248 159944
rect 328368 159928 328420 159934
rect 328368 159870 328420 159876
rect 327540 158772 327592 158778
rect 327540 158714 327592 158720
rect 327908 157004 327960 157010
rect 327908 156946 327960 156952
rect 326712 154148 326764 154154
rect 326712 154090 326764 154096
rect 327264 153264 327316 153270
rect 327264 153206 327316 153212
rect 326620 153060 326672 153066
rect 326620 153002 326672 153008
rect 325976 152448 326028 152454
rect 325976 152390 326028 152396
rect 326068 152448 326120 152454
rect 326068 152390 326120 152396
rect 325988 150226 326016 152390
rect 326632 150226 326660 153002
rect 327276 150226 327304 153206
rect 327920 150226 327948 156946
rect 321480 150198 321554 150226
rect 322124 150198 322198 150226
rect 322768 150198 322842 150226
rect 323412 150198 323486 150226
rect 324056 150198 324130 150226
rect 324700 150198 324774 150226
rect 325344 150198 325418 150226
rect 325988 150198 326062 150226
rect 326632 150198 326706 150226
rect 327276 150198 327350 150226
rect 327920 150198 327994 150226
rect 328472 150210 328500 159938
rect 328550 159488 328606 159497
rect 328550 159423 328606 159432
rect 328564 150226 328592 159423
rect 330128 155446 330156 163200
rect 330484 156936 330536 156942
rect 330484 156878 330536 156884
rect 330116 155440 330168 155446
rect 330116 155382 330168 155388
rect 329932 154420 329984 154426
rect 329932 154362 329984 154368
rect 329944 150226 329972 154362
rect 320882 149940 320910 150198
rect 321526 149940 321554 150198
rect 322170 149940 322198 150198
rect 322814 149940 322842 150198
rect 323458 149940 323486 150198
rect 324102 149940 324130 150198
rect 324746 149940 324774 150198
rect 325390 149940 325418 150198
rect 326034 149940 326062 150198
rect 326678 149940 326706 150198
rect 327322 149940 327350 150198
rect 327966 149940 327994 150198
rect 328460 150204 328512 150210
rect 328564 150198 328638 150226
rect 328460 150146 328512 150152
rect 328610 149940 328638 150198
rect 329242 150204 329294 150210
rect 329242 150146 329294 150152
rect 329898 150198 329972 150226
rect 330496 150226 330524 156878
rect 330956 153066 330984 163200
rect 330944 153060 330996 153066
rect 330944 153002 330996 153008
rect 331232 152318 331260 163254
rect 331692 163146 331720 163254
rect 331770 163200 331826 164400
rect 332598 163200 332654 164400
rect 333426 163200 333482 164400
rect 334254 163200 334310 164400
rect 335082 163200 335138 164400
rect 335372 163254 335952 163282
rect 331784 163146 331812 163200
rect 331692 163118 331812 163146
rect 332416 154352 332468 154358
rect 332416 154294 332468 154300
rect 331772 152924 331824 152930
rect 331772 152866 331824 152872
rect 331220 152312 331272 152318
rect 331220 152254 331272 152260
rect 331128 152108 331180 152114
rect 331128 152050 331180 152056
rect 331140 150226 331168 152050
rect 331784 150226 331812 152866
rect 332428 150226 332456 154294
rect 332612 152930 332640 163200
rect 332692 160064 332744 160070
rect 332692 160006 332744 160012
rect 332600 152924 332652 152930
rect 332600 152866 332652 152872
rect 330496 150198 330570 150226
rect 331140 150198 331214 150226
rect 331784 150198 331858 150226
rect 332428 150198 332502 150226
rect 332704 150210 332732 160006
rect 333060 157072 333112 157078
rect 333060 157014 333112 157020
rect 333072 150226 333100 157014
rect 333440 155514 333468 163200
rect 334268 160070 334296 163200
rect 334256 160064 334308 160070
rect 334256 160006 334308 160012
rect 335096 159322 335124 163200
rect 334348 159316 334400 159322
rect 334348 159258 334400 159264
rect 335084 159316 335136 159322
rect 335084 159258 335136 159264
rect 333428 155508 333480 155514
rect 333428 155450 333480 155456
rect 334360 150226 334388 159258
rect 334900 154556 334952 154562
rect 334900 154498 334952 154504
rect 334912 150226 334940 154498
rect 335372 152114 335400 163254
rect 335924 163146 335952 163254
rect 336002 163200 336058 164400
rect 336830 163200 336886 164400
rect 337658 163200 337714 164400
rect 338486 163200 338542 164400
rect 339314 163200 339370 164400
rect 339512 163254 340092 163282
rect 336016 163146 336044 163200
rect 335924 163118 336044 163146
rect 335544 157276 335596 157282
rect 335544 157218 335596 157224
rect 335360 152108 335412 152114
rect 335360 152050 335412 152056
rect 335556 150226 335584 157218
rect 336844 154358 336872 163200
rect 337672 155582 337700 163200
rect 338500 159118 338528 163200
rect 339328 159254 339356 163200
rect 338764 159248 338816 159254
rect 338764 159190 338816 159196
rect 339316 159248 339368 159254
rect 339316 159190 339368 159196
rect 338396 159112 338448 159118
rect 338396 159054 338448 159060
rect 338488 159112 338540 159118
rect 338488 159054 338540 159060
rect 338120 157140 338172 157146
rect 338120 157082 338172 157088
rect 337660 155576 337712 155582
rect 337660 155518 337712 155524
rect 337476 154488 337528 154494
rect 337476 154430 337528 154436
rect 336832 154352 336884 154358
rect 336832 154294 336884 154300
rect 336832 153196 336884 153202
rect 336832 153138 336884 153144
rect 336188 152244 336240 152250
rect 336188 152186 336240 152192
rect 336200 150226 336228 152186
rect 336844 150226 336872 153138
rect 337488 150226 337516 154430
rect 338132 150226 338160 157082
rect 329254 149940 329282 150146
rect 329898 149940 329926 150198
rect 330542 149940 330570 150198
rect 331186 149940 331214 150198
rect 331830 149940 331858 150198
rect 332474 149940 332502 150198
rect 332692 150204 332744 150210
rect 333072 150198 333146 150226
rect 332692 150146 332744 150152
rect 333118 149940 333146 150198
rect 333750 150204 333802 150210
rect 334360 150198 334434 150226
rect 334912 150198 334986 150226
rect 335556 150198 335630 150226
rect 336200 150198 336274 150226
rect 336844 150198 336918 150226
rect 337488 150198 337562 150226
rect 338132 150198 338206 150226
rect 338408 150210 338436 159054
rect 338776 150226 338804 159190
rect 339512 154290 339540 163254
rect 340064 163146 340092 163254
rect 340142 163200 340198 164400
rect 340970 163200 341026 164400
rect 341890 163200 341946 164400
rect 341996 163254 342208 163282
rect 340156 163146 340184 163200
rect 340064 163118 340184 163146
rect 339684 159112 339736 159118
rect 339684 159054 339736 159060
rect 339592 155780 339644 155786
rect 339592 155722 339644 155728
rect 339500 154284 339552 154290
rect 339500 154226 339552 154232
rect 339604 151814 339632 155722
rect 339696 153202 339724 159054
rect 340052 156732 340104 156738
rect 340052 156674 340104 156680
rect 339684 153196 339736 153202
rect 339684 153138 339736 153144
rect 340064 151814 340092 156674
rect 340984 155650 341012 163200
rect 341904 163146 341932 163200
rect 341996 163146 342024 163254
rect 341904 163118 342024 163146
rect 341616 159656 341668 159662
rect 341616 159598 341668 159604
rect 342180 159610 342208 163254
rect 342718 163200 342774 164400
rect 343546 163200 343602 164400
rect 344374 163200 344430 164400
rect 345202 163200 345258 164400
rect 346030 163200 346086 164400
rect 346412 163254 346808 163282
rect 342732 159730 342760 163200
rect 342628 159724 342680 159730
rect 342628 159666 342680 159672
rect 342720 159724 342772 159730
rect 342720 159666 342772 159672
rect 342640 159610 342668 159666
rect 342812 159656 342864 159662
rect 341628 159526 341656 159598
rect 342180 159582 342392 159610
rect 342640 159604 342812 159610
rect 342640 159598 342864 159604
rect 342640 159582 342852 159598
rect 341616 159520 341668 159526
rect 341616 159462 341668 159468
rect 342364 159458 342392 159582
rect 341432 159452 341484 159458
rect 341432 159394 341484 159400
rect 342260 159452 342312 159458
rect 342260 159394 342312 159400
rect 342352 159452 342404 159458
rect 342352 159394 342404 159400
rect 341444 159186 341472 159394
rect 341432 159180 341484 159186
rect 341432 159122 341484 159128
rect 340972 155644 341024 155650
rect 340972 155586 341024 155592
rect 342272 152998 342300 159394
rect 342444 159384 342496 159390
rect 342444 159326 342496 159332
rect 342352 155848 342404 155854
rect 342352 155790 342404 155796
rect 341340 152992 341392 152998
rect 341340 152934 341392 152940
rect 342260 152992 342312 152998
rect 342260 152934 342312 152940
rect 339604 151786 340000 151814
rect 340064 151786 340736 151814
rect 339972 150226 340000 151786
rect 340708 150226 340736 151786
rect 341352 150226 341380 152934
rect 341984 152380 342036 152386
rect 341984 152322 342036 152328
rect 341996 150226 342024 152322
rect 342364 151814 342392 155790
rect 342456 152250 342484 159326
rect 342536 156868 342588 156874
rect 342536 156810 342588 156816
rect 342444 152244 342496 152250
rect 342444 152186 342496 152192
rect 342548 151814 342576 156810
rect 343560 154222 343588 163200
rect 343824 159724 343876 159730
rect 343824 159666 343876 159672
rect 343548 154216 343600 154222
rect 343548 154158 343600 154164
rect 343836 152386 343864 159666
rect 344388 155718 344416 163200
rect 345216 157334 345244 163200
rect 346044 159390 346072 163200
rect 346032 159384 346084 159390
rect 345584 159310 345796 159338
rect 346032 159326 346084 159332
rect 345584 159050 345612 159310
rect 345768 159186 345796 159310
rect 345664 159180 345716 159186
rect 345664 159122 345716 159128
rect 345756 159180 345808 159186
rect 345756 159122 345808 159128
rect 345676 159066 345704 159122
rect 345676 159050 345888 159066
rect 345572 159044 345624 159050
rect 345676 159044 345900 159050
rect 345676 159038 345848 159044
rect 345572 158986 345624 158992
rect 345848 158986 345900 158992
rect 345216 157306 345336 157334
rect 345112 156800 345164 156806
rect 345112 156742 345164 156748
rect 344376 155712 344428 155718
rect 344376 155654 344428 155660
rect 343916 152992 343968 152998
rect 343916 152934 343968 152940
rect 343824 152380 343876 152386
rect 343824 152322 343876 152328
rect 342364 151786 342484 151814
rect 342548 151786 343312 151814
rect 342456 150226 342484 151786
rect 343284 150226 343312 151786
rect 343928 150226 343956 152934
rect 344560 152244 344612 152250
rect 344560 152186 344612 152192
rect 344572 150226 344600 152186
rect 333750 150146 333802 150152
rect 333762 149940 333790 150146
rect 334406 149940 334434 150198
rect 334958 149940 334986 150198
rect 335602 149940 335630 150198
rect 336246 149940 336274 150198
rect 336890 149940 336918 150198
rect 337534 149940 337562 150198
rect 338178 149940 338206 150198
rect 338396 150204 338448 150210
rect 338776 150198 338850 150226
rect 338396 150146 338448 150152
rect 338822 149940 338850 150198
rect 339454 150204 339506 150210
rect 339972 150198 340138 150226
rect 340708 150198 340782 150226
rect 341352 150198 341426 150226
rect 341996 150198 342070 150226
rect 342456 150198 342714 150226
rect 343284 150198 343358 150226
rect 343928 150198 344002 150226
rect 344572 150198 344646 150226
rect 345124 150210 345152 156742
rect 345204 155916 345256 155922
rect 345204 155858 345256 155864
rect 345216 150226 345244 155858
rect 345308 152998 345336 157306
rect 346412 154426 346440 163254
rect 346780 163146 346808 163254
rect 346858 163200 346914 164400
rect 347778 163200 347834 164400
rect 348160 163254 348556 163282
rect 346872 163146 346900 163200
rect 346780 163118 346900 163146
rect 347792 159730 347820 163200
rect 347780 159724 347832 159730
rect 347780 159666 347832 159672
rect 348056 157208 348108 157214
rect 348056 157150 348108 157156
rect 347872 155304 347924 155310
rect 347872 155246 347924 155252
rect 346400 154420 346452 154426
rect 346400 154362 346452 154368
rect 345296 152992 345348 152998
rect 345296 152934 345348 152940
rect 347136 152516 347188 152522
rect 347136 152458 347188 152464
rect 346492 151836 346544 151842
rect 346492 151778 346544 151784
rect 346504 150226 346532 151778
rect 347148 150226 347176 152458
rect 347884 150226 347912 155246
rect 348068 151814 348096 157150
rect 348160 152522 348188 163254
rect 348528 163146 348556 163254
rect 348606 163200 348662 164400
rect 349172 163254 349384 163282
rect 348620 163146 348648 163200
rect 348528 163118 348648 163146
rect 349068 159044 349120 159050
rect 349068 158986 349120 158992
rect 348148 152516 348200 152522
rect 348148 152458 348200 152464
rect 348068 151786 348464 151814
rect 339454 150146 339506 150152
rect 339466 149940 339494 150146
rect 340110 149940 340138 150198
rect 340754 149940 340782 150198
rect 341398 149940 341426 150198
rect 342042 149940 342070 150198
rect 342686 149940 342714 150198
rect 343330 149940 343358 150198
rect 343974 149940 344002 150198
rect 344618 149940 344646 150198
rect 345112 150204 345164 150210
rect 345216 150198 345290 150226
rect 345112 150146 345164 150152
rect 345262 149940 345290 150198
rect 345894 150204 345946 150210
rect 346504 150198 346578 150226
rect 347148 150198 347222 150226
rect 345894 150146 345946 150152
rect 345906 149940 345934 150146
rect 346550 149940 346578 150198
rect 347194 149940 347222 150198
rect 347838 150198 347912 150226
rect 348436 150226 348464 151786
rect 349080 150226 349108 158986
rect 349172 152250 349200 163254
rect 349356 163146 349384 163254
rect 349434 163200 349490 164400
rect 349540 163254 350212 163282
rect 349448 163146 349476 163200
rect 349356 163118 349476 163146
rect 349344 159452 349396 159458
rect 349344 159394 349396 159400
rect 349356 159118 349384 159394
rect 349252 159112 349304 159118
rect 349252 159054 349304 159060
rect 349344 159112 349396 159118
rect 349344 159054 349396 159060
rect 349160 152244 349212 152250
rect 349160 152186 349212 152192
rect 349264 151814 349292 159054
rect 349540 154494 349568 163254
rect 350184 163146 350212 163254
rect 350262 163200 350318 164400
rect 351090 163200 351146 164400
rect 351918 163200 351974 164400
rect 352024 163254 352696 163282
rect 350276 163146 350304 163200
rect 350184 163118 350304 163146
rect 351104 159050 351132 163200
rect 351932 159186 351960 163200
rect 351828 159180 351880 159186
rect 351828 159122 351880 159128
rect 351920 159180 351972 159186
rect 351920 159122 351972 159128
rect 351840 159066 351868 159122
rect 351092 159044 351144 159050
rect 351840 159038 351960 159066
rect 351092 158986 351144 158992
rect 350356 155100 350408 155106
rect 350356 155042 350408 155048
rect 349528 154488 349580 154494
rect 349528 154430 349580 154436
rect 349804 152380 349856 152386
rect 349804 152322 349856 152328
rect 349896 152380 349948 152386
rect 349896 152322 349948 152328
rect 349816 151842 349844 152322
rect 349908 152250 349936 152322
rect 349896 152244 349948 152250
rect 349896 152186 349948 152192
rect 349804 151836 349856 151842
rect 349264 151786 349752 151814
rect 349724 150226 349752 151786
rect 349804 151778 349856 151784
rect 350368 150226 350396 155042
rect 351000 152584 351052 152590
rect 351000 152526 351052 152532
rect 351012 150226 351040 152526
rect 351932 152250 351960 159038
rect 352024 152590 352052 163254
rect 352668 163146 352696 163254
rect 352746 163200 352802 164400
rect 353666 163200 353722 164400
rect 354494 163200 354550 164400
rect 354692 163254 355272 163282
rect 352760 163146 352788 163200
rect 352668 163118 352788 163146
rect 352472 155236 352524 155242
rect 352472 155178 352524 155184
rect 352012 152584 352064 152590
rect 352012 152526 352064 152532
rect 351920 152244 351972 152250
rect 351920 152186 351972 152192
rect 351644 151972 351696 151978
rect 351644 151914 351696 151920
rect 351656 150226 351684 151914
rect 352288 151904 352340 151910
rect 352288 151846 352340 151852
rect 352300 150226 352328 151846
rect 352484 151814 352512 155178
rect 353680 154562 353708 163200
rect 354220 159656 354272 159662
rect 354220 159598 354272 159604
rect 353668 154556 353720 154562
rect 353668 154498 353720 154504
rect 353484 152244 353536 152250
rect 353484 152186 353536 152192
rect 353496 151814 353524 152186
rect 352484 151786 352972 151814
rect 353496 151786 353616 151814
rect 352944 150226 352972 151786
rect 353588 150226 353616 151786
rect 354232 150226 354260 159598
rect 354508 152250 354536 163200
rect 354496 152244 354548 152250
rect 354496 152186 354548 152192
rect 354692 151978 354720 163254
rect 355244 163146 355272 163254
rect 355322 163200 355378 164400
rect 356150 163200 356206 164400
rect 356256 163254 356928 163282
rect 355336 163146 355364 163200
rect 355244 163118 355364 163146
rect 356164 159526 356192 163200
rect 354864 159520 354916 159526
rect 354864 159462 354916 159468
rect 356152 159520 356204 159526
rect 356152 159462 356204 159468
rect 354680 151972 354732 151978
rect 354680 151914 354732 151920
rect 354876 150226 354904 159462
rect 356256 153882 356284 163254
rect 356900 163146 356928 163254
rect 356978 163200 357034 164400
rect 357806 163200 357862 164400
rect 358634 163200 358690 164400
rect 358832 163254 359504 163282
rect 356992 163146 357020 163200
rect 356900 163118 357020 163146
rect 357440 159656 357492 159662
rect 357440 159598 357492 159604
rect 357452 158846 357480 159598
rect 357820 158982 357848 163200
rect 357992 159792 358044 159798
rect 357992 159734 358044 159740
rect 357532 158976 357584 158982
rect 357532 158918 357584 158924
rect 357808 158976 357860 158982
rect 357808 158918 357860 158924
rect 357440 158840 357492 158846
rect 357440 158782 357492 158788
rect 355508 153876 355560 153882
rect 355508 153818 355560 153824
rect 356244 153876 356296 153882
rect 356244 153818 356296 153824
rect 355520 150226 355548 153818
rect 356152 152720 356204 152726
rect 356152 152662 356204 152668
rect 356164 150226 356192 152662
rect 357438 152416 357494 152425
rect 357438 152351 357494 152360
rect 356796 152176 356848 152182
rect 356796 152118 356848 152124
rect 356808 150226 356836 152118
rect 357452 150226 357480 152351
rect 357544 152182 357572 158918
rect 357900 154012 357952 154018
rect 357900 153954 357952 153960
rect 357532 152176 357584 152182
rect 357532 152118 357584 152124
rect 357912 150498 357940 153954
rect 358004 151814 358032 159734
rect 358648 159458 358676 163200
rect 358636 159452 358688 159458
rect 358636 159394 358688 159400
rect 358832 152726 358860 163254
rect 359476 163146 359504 163254
rect 359554 163200 359610 164400
rect 360382 163200 360438 164400
rect 361210 163200 361266 164400
rect 361592 163254 361988 163282
rect 359568 163146 359596 163200
rect 359476 163118 359596 163146
rect 358912 159588 358964 159594
rect 358912 159530 358964 159536
rect 358820 152720 358872 152726
rect 358820 152662 358872 152668
rect 358004 151786 358768 151814
rect 357912 150470 358124 150498
rect 358096 150226 358124 150470
rect 358740 150226 358768 151786
rect 348436 150198 348510 150226
rect 349080 150198 349154 150226
rect 349724 150198 349798 150226
rect 350368 150198 350442 150226
rect 351012 150198 351086 150226
rect 351656 150198 351730 150226
rect 352300 150198 352374 150226
rect 352944 150198 353018 150226
rect 353588 150198 353662 150226
rect 354232 150198 354306 150226
rect 354876 150198 354950 150226
rect 355520 150198 355594 150226
rect 356164 150198 356238 150226
rect 356808 150198 356882 150226
rect 357452 150198 357526 150226
rect 358096 150198 358170 150226
rect 358740 150198 358814 150226
rect 358924 150210 358952 159530
rect 360396 153814 360424 163200
rect 361224 158914 361252 163200
rect 361212 158908 361264 158914
rect 361212 158850 361264 158856
rect 360660 153944 360712 153950
rect 360660 153886 360712 153892
rect 360384 153808 360436 153814
rect 360384 153750 360436 153756
rect 359372 152176 359424 152182
rect 359372 152118 359424 152124
rect 359384 150226 359412 152118
rect 360672 150226 360700 153886
rect 361592 152862 361620 163254
rect 361960 163146 361988 163254
rect 362038 163200 362094 164400
rect 362866 163200 362922 164400
rect 363064 163254 363644 163282
rect 362052 163146 362080 163200
rect 361960 163118 362080 163146
rect 362880 159594 362908 163200
rect 362868 159588 362920 159594
rect 362868 159530 362920 159536
rect 362960 158840 363012 158846
rect 362960 158782 363012 158788
rect 361304 152856 361356 152862
rect 361304 152798 361356 152804
rect 361580 152856 361632 152862
rect 361580 152798 361632 152804
rect 361316 150226 361344 152798
rect 361948 152652 362000 152658
rect 361948 152594 362000 152600
rect 361960 150226 361988 152594
rect 362592 152040 362644 152046
rect 362592 151982 362644 151988
rect 362604 150226 362632 151982
rect 347838 149940 347866 150198
rect 348482 149940 348510 150198
rect 349126 149940 349154 150198
rect 349770 149940 349798 150198
rect 350414 149940 350442 150198
rect 351058 149940 351086 150198
rect 351702 149940 351730 150198
rect 352346 149940 352374 150198
rect 352990 149940 353018 150198
rect 353634 149940 353662 150198
rect 354278 149940 354306 150198
rect 354922 149940 354950 150198
rect 355566 149940 355594 150198
rect 356210 149940 356238 150198
rect 356854 149940 356882 150198
rect 357498 149940 357526 150198
rect 358142 149940 358170 150198
rect 358786 149940 358814 150198
rect 358912 150204 358964 150210
rect 359384 150198 359458 150226
rect 358912 150146 358964 150152
rect 359430 149940 359458 150198
rect 360062 150204 360114 150210
rect 360672 150198 360746 150226
rect 361316 150198 361390 150226
rect 361960 150198 362034 150226
rect 362604 150198 362678 150226
rect 362972 150210 363000 158782
rect 363064 153950 363092 163254
rect 363616 163146 363644 163254
rect 363694 163200 363750 164400
rect 364522 163200 364578 164400
rect 365442 163200 365498 164400
rect 365732 163254 366220 163282
rect 363708 163146 363736 163200
rect 363616 163118 363736 163146
rect 363144 159656 363196 159662
rect 363144 159598 363196 159604
rect 363052 153944 363104 153950
rect 363052 153886 363104 153892
rect 363156 151910 363184 159598
rect 363236 155372 363288 155378
rect 363236 155314 363288 155320
rect 363144 151904 363196 151910
rect 363144 151846 363196 151852
rect 363248 150226 363276 155314
rect 364536 152182 364564 163200
rect 365168 159860 365220 159866
rect 365168 159802 365220 159808
rect 364524 152176 364576 152182
rect 364524 152118 364576 152124
rect 364524 151904 364576 151910
rect 364524 151846 364576 151852
rect 364536 150226 364564 151846
rect 365180 150226 365208 159802
rect 365456 159798 365484 163200
rect 365444 159792 365496 159798
rect 365444 159734 365496 159740
rect 365732 152658 365760 163254
rect 366192 163146 366220 163254
rect 366270 163200 366326 164400
rect 367098 163200 367154 164400
rect 367926 163200 367982 164400
rect 368492 163254 368704 163282
rect 366284 163146 366312 163200
rect 366192 163118 366312 163146
rect 365812 154080 365864 154086
rect 365812 154022 365864 154028
rect 365720 152652 365772 152658
rect 365720 152594 365772 152600
rect 365824 150226 365852 154022
rect 367112 154018 367140 163200
rect 367940 158846 367968 163200
rect 367928 158840 367980 158846
rect 367928 158782 367980 158788
rect 367192 158772 367244 158778
rect 367192 158714 367244 158720
rect 367100 154012 367152 154018
rect 367100 153954 367152 153960
rect 367204 153134 367232 158714
rect 368296 154148 368348 154154
rect 368296 154090 368348 154096
rect 367008 153128 367060 153134
rect 367008 153070 367060 153076
rect 367192 153128 367244 153134
rect 367192 153070 367244 153076
rect 366364 152788 366416 152794
rect 366364 152730 366416 152736
rect 360062 150146 360114 150152
rect 360074 149940 360102 150146
rect 360718 149940 360746 150198
rect 361362 149940 361390 150198
rect 362006 149940 362034 150198
rect 362650 149940 362678 150198
rect 362960 150204 363012 150210
rect 363248 150198 363322 150226
rect 362960 150146 363012 150152
rect 363294 149940 363322 150198
rect 363926 150204 363978 150210
rect 364536 150198 364610 150226
rect 365180 150198 365254 150226
rect 363926 150146 363978 150152
rect 363938 149940 363966 150146
rect 364582 149940 364610 150198
rect 365226 149940 365254 150198
rect 365778 150198 365852 150226
rect 366376 150226 366404 152730
rect 367020 150226 367048 153070
rect 367652 152448 367704 152454
rect 367652 152390 367704 152396
rect 367664 150226 367692 152390
rect 368308 150226 368336 154090
rect 368492 152794 368520 163254
rect 368676 163146 368704 163254
rect 368754 163200 368810 164400
rect 369582 163200 369638 164400
rect 370410 163200 370466 164400
rect 371330 163200 371386 164400
rect 372158 163200 372214 164400
rect 372632 163254 372936 163282
rect 368768 163146 368796 163200
rect 368676 163118 368796 163146
rect 369492 159928 369544 159934
rect 369492 159870 369544 159876
rect 368940 153128 368992 153134
rect 368940 153070 368992 153076
rect 368480 152788 368532 152794
rect 368480 152730 368532 152736
rect 368952 150226 368980 153070
rect 369504 151814 369532 159870
rect 369596 159662 369624 163200
rect 369952 159996 370004 160002
rect 369952 159938 370004 159944
rect 369584 159656 369636 159662
rect 369584 159598 369636 159604
rect 369964 151814 369992 159938
rect 370424 155242 370452 163200
rect 370872 155440 370924 155446
rect 370872 155382 370924 155388
rect 370412 155236 370464 155242
rect 370412 155178 370464 155184
rect 369504 151786 369624 151814
rect 369964 151786 370268 151814
rect 369596 150226 369624 151786
rect 370240 150226 370268 151786
rect 370884 150226 370912 155382
rect 371344 152454 371372 163200
rect 372172 159934 372200 163200
rect 372160 159928 372212 159934
rect 372160 159870 372212 159876
rect 372632 153066 372660 163254
rect 372908 163146 372936 163254
rect 372986 163200 373042 164400
rect 373814 163200 373870 164400
rect 374642 163200 374698 164400
rect 375470 163200 375526 164400
rect 376298 163200 376354 164400
rect 376864 163254 377168 163282
rect 373000 163146 373028 163200
rect 372908 163118 373028 163146
rect 373448 155508 373500 155514
rect 373448 155450 373500 155456
rect 371516 153060 371568 153066
rect 371516 153002 371568 153008
rect 372620 153060 372672 153066
rect 372620 153002 372672 153008
rect 371332 152448 371384 152454
rect 371332 152390 371384 152396
rect 371528 150226 371556 153002
rect 372804 152924 372856 152930
rect 372804 152866 372856 152872
rect 372160 152312 372212 152318
rect 372160 152254 372212 152260
rect 372172 150226 372200 152254
rect 372816 150226 372844 152866
rect 373460 150226 373488 155450
rect 373828 155310 373856 163200
rect 374092 160064 374144 160070
rect 374092 160006 374144 160012
rect 373816 155304 373868 155310
rect 373816 155246 373868 155252
rect 374104 150226 374132 160006
rect 374656 160002 374684 163200
rect 374644 159996 374696 160002
rect 374644 159938 374696 159944
rect 374736 159316 374788 159322
rect 374736 159258 374788 159264
rect 374748 150226 374776 159258
rect 375484 153134 375512 163200
rect 376312 159866 376340 163200
rect 376300 159860 376352 159866
rect 376300 159802 376352 159808
rect 376760 158908 376812 158914
rect 376760 158850 376812 158856
rect 376772 158642 376800 158850
rect 376760 158636 376812 158642
rect 376760 158578 376812 158584
rect 375564 155576 375616 155582
rect 375564 155518 375616 155524
rect 375472 153128 375524 153134
rect 375472 153070 375524 153076
rect 375380 152108 375432 152114
rect 375380 152050 375432 152056
rect 375392 150226 375420 152050
rect 366376 150198 366450 150226
rect 367020 150198 367094 150226
rect 367664 150198 367738 150226
rect 368308 150198 368382 150226
rect 368952 150198 369026 150226
rect 369596 150198 369670 150226
rect 370240 150198 370314 150226
rect 370884 150198 370958 150226
rect 371528 150198 371602 150226
rect 372172 150198 372246 150226
rect 372816 150198 372890 150226
rect 373460 150198 373534 150226
rect 374104 150198 374178 150226
rect 374748 150198 374822 150226
rect 375392 150198 375466 150226
rect 375576 150210 375604 155518
rect 376024 154352 376076 154358
rect 376024 154294 376076 154300
rect 376036 150226 376064 154294
rect 376864 154154 376892 163254
rect 377140 163146 377168 163254
rect 377218 163200 377274 164400
rect 378046 163200 378102 164400
rect 378874 163200 378930 164400
rect 379702 163200 379758 164400
rect 380176 163254 380480 163282
rect 377232 163146 377260 163200
rect 377140 163118 377260 163146
rect 377956 159248 378008 159254
rect 377956 159190 378008 159196
rect 376944 159112 376996 159118
rect 376944 159054 376996 159060
rect 376956 158914 376984 159054
rect 376944 158908 376996 158914
rect 376944 158850 376996 158856
rect 376852 154148 376904 154154
rect 376852 154090 376904 154096
rect 377312 153196 377364 153202
rect 377312 153138 377364 153144
rect 377324 150226 377352 153138
rect 377968 150226 377996 159190
rect 378060 159118 378088 163200
rect 378888 160070 378916 163200
rect 378876 160064 378928 160070
rect 378876 160006 378928 160012
rect 379716 159730 379744 163200
rect 378784 159724 378836 159730
rect 378784 159666 378836 159672
rect 379704 159724 379756 159730
rect 379704 159666 379756 159672
rect 378048 159112 378100 159118
rect 378048 159054 378100 159060
rect 378232 158908 378284 158914
rect 378232 158850 378284 158856
rect 378140 155644 378192 155650
rect 378140 155586 378192 155592
rect 365778 149940 365806 150198
rect 366422 149940 366450 150198
rect 367066 149940 367094 150198
rect 367710 149940 367738 150198
rect 368354 149940 368382 150198
rect 368998 149940 369026 150198
rect 369642 149940 369670 150198
rect 370286 149940 370314 150198
rect 370930 149940 370958 150198
rect 371574 149940 371602 150198
rect 372218 149940 372246 150198
rect 372862 149940 372890 150198
rect 373506 149940 373534 150198
rect 374150 149940 374178 150198
rect 374794 149940 374822 150198
rect 375438 149940 375466 150198
rect 375564 150204 375616 150210
rect 376036 150198 376110 150226
rect 375564 150146 375616 150152
rect 376082 149940 376110 150198
rect 376714 150204 376766 150210
rect 377324 150198 377398 150226
rect 377968 150198 378042 150226
rect 378152 150210 378180 155586
rect 378244 153202 378272 158850
rect 378600 154284 378652 154290
rect 378600 154226 378652 154232
rect 378232 153196 378284 153202
rect 378232 153138 378284 153144
rect 378612 150226 378640 154226
rect 378796 152046 378824 159666
rect 380176 154086 380204 163254
rect 380452 163146 380480 163254
rect 380530 163200 380586 164400
rect 381004 163254 381308 163282
rect 380544 163146 380572 163200
rect 380452 163118 380572 163146
rect 380164 154080 380216 154086
rect 380164 154022 380216 154028
rect 381004 153202 381032 163254
rect 381280 163146 381308 163254
rect 381358 163200 381414 164400
rect 382186 163200 382242 164400
rect 383106 163200 383162 164400
rect 383672 163254 383884 163282
rect 381372 163146 381400 163200
rect 381280 163118 381400 163146
rect 381820 155712 381872 155718
rect 381820 155654 381872 155660
rect 381176 154216 381228 154222
rect 381176 154158 381228 154164
rect 379888 153196 379940 153202
rect 379888 153138 379940 153144
rect 380992 153196 381044 153202
rect 380992 153138 381044 153144
rect 378784 152040 378836 152046
rect 378784 151982 378836 151988
rect 379900 150226 379928 153138
rect 380532 151836 380584 151842
rect 380532 151778 380584 151784
rect 380544 150226 380572 151778
rect 381188 150226 381216 154158
rect 381832 150226 381860 155654
rect 382200 152930 382228 163200
rect 383120 159390 383148 163200
rect 382832 159384 382884 159390
rect 382832 159326 382884 159332
rect 383108 159384 383160 159390
rect 383108 159326 383160 159332
rect 382556 159044 382608 159050
rect 382556 158986 382608 158992
rect 382568 152998 382596 158986
rect 382464 152992 382516 152998
rect 382464 152934 382516 152940
rect 382556 152992 382608 152998
rect 382556 152934 382608 152940
rect 382188 152924 382240 152930
rect 382188 152866 382240 152872
rect 382476 150226 382504 152934
rect 382844 151814 382872 159326
rect 383672 154222 383700 163254
rect 383856 163146 383884 163254
rect 383934 163200 383990 164400
rect 384762 163200 384818 164400
rect 385590 163200 385646 164400
rect 386418 163200 386474 164400
rect 386524 163254 387196 163282
rect 383948 163146 383976 163200
rect 383856 163118 383976 163146
rect 384776 158778 384804 163200
rect 385604 159254 385632 163200
rect 385500 159248 385552 159254
rect 385500 159190 385552 159196
rect 385592 159248 385644 159254
rect 385592 159190 385644 159196
rect 384948 158976 385000 158982
rect 384948 158918 385000 158924
rect 384764 158772 384816 158778
rect 384764 158714 384816 158720
rect 383752 154420 383804 154426
rect 383752 154362 383804 154368
rect 383660 154216 383712 154222
rect 383660 154158 383712 154164
rect 382844 151786 383148 151814
rect 383120 150226 383148 151786
rect 383764 150226 383792 154362
rect 384960 152318 384988 158918
rect 385512 152522 385540 159190
rect 386144 158908 386196 158914
rect 386144 158850 386196 158856
rect 385040 152516 385092 152522
rect 385040 152458 385092 152464
rect 385500 152516 385552 152522
rect 385500 152458 385552 152464
rect 384948 152312 385000 152318
rect 384948 152254 385000 152260
rect 384396 152040 384448 152046
rect 384396 151982 384448 151988
rect 384408 150226 384436 151982
rect 385052 150226 385080 152458
rect 385684 152380 385736 152386
rect 385684 152322 385736 152328
rect 385696 150226 385724 152322
rect 386156 151910 386184 158850
rect 386236 158840 386288 158846
rect 386236 158782 386288 158788
rect 386144 151904 386196 151910
rect 386144 151846 386196 151852
rect 386248 151842 386276 158782
rect 386328 154488 386380 154494
rect 386328 154430 386380 154436
rect 386236 151836 386288 151842
rect 386236 151778 386288 151784
rect 386340 150226 386368 154430
rect 386432 152386 386460 163200
rect 386524 154290 386552 163254
rect 387168 163146 387196 163254
rect 387246 163200 387302 164400
rect 388074 163200 388130 164400
rect 388994 163200 389050 164400
rect 389822 163200 389878 164400
rect 390650 163200 390706 164400
rect 391478 163200 391534 164400
rect 392306 163200 392362 164400
rect 393134 163200 393190 164400
rect 393332 163254 393912 163282
rect 387260 163146 387288 163200
rect 387168 163118 387288 163146
rect 388088 158846 388116 163200
rect 388352 159996 388404 160002
rect 388352 159938 388404 159944
rect 388076 158840 388128 158846
rect 388076 158782 388128 158788
rect 386512 154284 386564 154290
rect 386512 154226 386564 154232
rect 386972 152992 387024 152998
rect 386972 152934 387024 152940
rect 386420 152380 386472 152386
rect 386420 152322 386472 152328
rect 386984 150226 387012 152934
rect 388260 152584 388312 152590
rect 388260 152526 388312 152532
rect 387616 152516 387668 152522
rect 387616 152458 387668 152464
rect 387708 152516 387760 152522
rect 387708 152458 387760 152464
rect 387628 150226 387656 152458
rect 387720 152386 387748 152458
rect 387708 152380 387760 152386
rect 387708 152322 387760 152328
rect 388272 150226 388300 152526
rect 388364 152046 388392 159938
rect 389008 159322 389036 163200
rect 389836 160002 389864 163200
rect 389824 159996 389876 160002
rect 389824 159938 389876 159944
rect 390560 159520 390612 159526
rect 390560 159462 390612 159468
rect 388996 159316 389048 159322
rect 388996 159258 389048 159264
rect 388444 159180 388496 159186
rect 388444 159122 388496 159128
rect 388456 152114 388484 159122
rect 390376 158840 390428 158846
rect 390376 158782 390428 158788
rect 389180 158772 389232 158778
rect 389180 158714 389232 158720
rect 388904 154556 388956 154562
rect 388904 154498 388956 154504
rect 388444 152108 388496 152114
rect 388444 152050 388496 152056
rect 388352 152040 388404 152046
rect 388352 151982 388404 151988
rect 388916 150226 388944 154498
rect 389192 152386 389220 158714
rect 390388 152998 390416 158782
rect 390376 152992 390428 152998
rect 390376 152934 390428 152940
rect 389180 152380 389232 152386
rect 389180 152322 389232 152328
rect 389548 152244 389600 152250
rect 389548 152186 389600 152192
rect 389560 150226 389588 152186
rect 390192 151972 390244 151978
rect 390192 151914 390244 151920
rect 390204 150226 390232 151914
rect 390572 151814 390600 159462
rect 390664 154494 390692 163200
rect 391492 158914 391520 163200
rect 392320 159186 392348 163200
rect 392768 159452 392820 159458
rect 392768 159394 392820 159400
rect 392308 159180 392360 159186
rect 392308 159122 392360 159128
rect 391480 158908 391532 158914
rect 391480 158850 391532 158856
rect 390652 154488 390704 154494
rect 390652 154430 390704 154436
rect 391480 153876 391532 153882
rect 391480 153818 391532 153824
rect 390572 151786 390876 151814
rect 390848 150226 390876 151786
rect 391492 150226 391520 153818
rect 392124 152312 392176 152318
rect 392124 152254 392176 152260
rect 392136 150226 392164 152254
rect 392780 150226 392808 159394
rect 393148 152590 393176 163200
rect 393332 154426 393360 163254
rect 393884 163146 393912 163254
rect 393962 163200 394018 164400
rect 394882 163200 394938 164400
rect 395710 163200 395766 164400
rect 396538 163200 396594 164400
rect 397366 163200 397422 164400
rect 397472 163254 398144 163282
rect 393976 163146 394004 163200
rect 393884 163118 394004 163146
rect 393688 158908 393740 158914
rect 393688 158850 393740 158856
rect 393320 154420 393372 154426
rect 393320 154362 393372 154368
rect 393412 152720 393464 152726
rect 393412 152662 393464 152668
rect 393136 152584 393188 152590
rect 393136 152526 393188 152532
rect 393424 150226 393452 152662
rect 393700 152318 393728 158850
rect 394056 153808 394108 153814
rect 394056 153750 394108 153756
rect 393688 152312 393740 152318
rect 393688 152254 393740 152260
rect 394068 150226 394096 153750
rect 394896 152726 394924 163200
rect 395528 159792 395580 159798
rect 395528 159734 395580 159740
rect 394976 159588 395028 159594
rect 394976 159530 395028 159536
rect 394884 152720 394936 152726
rect 394884 152662 394936 152668
rect 394700 151836 394752 151842
rect 394700 151778 394752 151784
rect 394712 150226 394740 151778
rect 376714 150146 376766 150152
rect 376726 149940 376754 150146
rect 377370 149940 377398 150198
rect 378014 149940 378042 150198
rect 378140 150204 378192 150210
rect 378612 150198 378686 150226
rect 378140 150146 378192 150152
rect 378658 149940 378686 150198
rect 379290 150204 379342 150210
rect 379900 150198 379974 150226
rect 380544 150198 380618 150226
rect 381188 150198 381262 150226
rect 381832 150198 381906 150226
rect 382476 150198 382550 150226
rect 383120 150198 383194 150226
rect 383764 150198 383838 150226
rect 384408 150198 384482 150226
rect 385052 150198 385126 150226
rect 385696 150198 385770 150226
rect 386340 150198 386414 150226
rect 386984 150198 387058 150226
rect 387628 150198 387702 150226
rect 388272 150198 388346 150226
rect 388916 150198 388990 150226
rect 389560 150198 389634 150226
rect 390204 150198 390278 150226
rect 390848 150198 390922 150226
rect 391492 150198 391566 150226
rect 392136 150198 392210 150226
rect 392780 150198 392854 150226
rect 393424 150198 393498 150226
rect 394068 150198 394142 150226
rect 394712 150198 394786 150226
rect 394988 150210 395016 159530
rect 395540 152862 395568 159734
rect 395724 159118 395752 163200
rect 396172 159928 396224 159934
rect 396172 159870 396224 159876
rect 395712 159112 395764 159118
rect 395712 159054 395764 159060
rect 395252 152856 395304 152862
rect 395252 152798 395304 152804
rect 395528 152856 395580 152862
rect 395528 152798 395580 152804
rect 395264 151814 395292 152798
rect 396184 151978 396212 159870
rect 396552 159798 396580 163200
rect 396540 159792 396592 159798
rect 396540 159734 396592 159740
rect 397380 154358 397408 163200
rect 397368 154352 397420 154358
rect 397368 154294 397420 154300
rect 396540 153944 396592 153950
rect 396540 153886 396592 153892
rect 396172 151972 396224 151978
rect 396172 151914 396224 151920
rect 395264 151786 395384 151814
rect 395356 150226 395384 151786
rect 396552 150226 396580 153886
rect 397472 153882 397500 163254
rect 398116 163146 398144 163254
rect 398194 163200 398250 164400
rect 399022 163200 399078 164400
rect 399220 163254 399800 163282
rect 398208 163146 398236 163200
rect 398116 163118 398236 163146
rect 398104 160064 398156 160070
rect 398104 160006 398156 160012
rect 397460 153876 397512 153882
rect 397460 153818 397512 153824
rect 397828 152856 397880 152862
rect 397828 152798 397880 152804
rect 397184 152176 397236 152182
rect 397184 152118 397236 152124
rect 397196 150226 397224 152118
rect 397840 150226 397868 152798
rect 398116 152250 398144 160006
rect 399036 159594 399064 163200
rect 399024 159588 399076 159594
rect 399024 159530 399076 159536
rect 398840 159248 398892 159254
rect 398840 159190 398892 159196
rect 398472 152652 398524 152658
rect 398472 152594 398524 152600
rect 398104 152244 398156 152250
rect 398104 152186 398156 152192
rect 398484 150226 398512 152594
rect 398852 151842 398880 159190
rect 399116 154012 399168 154018
rect 399116 153954 399168 153960
rect 398840 151836 398892 151842
rect 398840 151778 398892 151784
rect 399128 150226 399156 153954
rect 399220 152658 399248 163254
rect 399772 163146 399800 163254
rect 399850 163200 399906 164400
rect 400770 163200 400826 164400
rect 401598 163200 401654 164400
rect 402426 163200 402482 164400
rect 403254 163200 403310 164400
rect 404082 163200 404138 164400
rect 404372 163254 404860 163282
rect 399864 163146 399892 163200
rect 399772 163118 399892 163146
rect 400784 159526 400812 163200
rect 401048 159656 401100 159662
rect 401048 159598 401100 159604
rect 400772 159520 400824 159526
rect 400772 159462 400824 159468
rect 400404 152788 400456 152794
rect 400404 152730 400456 152736
rect 399208 152652 399260 152658
rect 399208 152594 399260 152600
rect 399760 151904 399812 151910
rect 399760 151846 399812 151852
rect 399772 150226 399800 151846
rect 400416 150226 400444 152730
rect 401060 150226 401088 159598
rect 401612 153950 401640 163200
rect 401784 155236 401836 155242
rect 401784 155178 401836 155184
rect 401600 153944 401652 153950
rect 401600 153886 401652 153892
rect 401796 150226 401824 155178
rect 402440 152862 402468 163200
rect 403268 159934 403296 163200
rect 403256 159928 403308 159934
rect 403256 159870 403308 159876
rect 404096 159458 404124 163200
rect 404084 159452 404136 159458
rect 404084 159394 404136 159400
rect 403900 159316 403952 159322
rect 403900 159258 403952 159264
rect 403164 155304 403216 155310
rect 403164 155246 403216 155252
rect 402428 152856 402480 152862
rect 402428 152798 402480 152804
rect 402336 152448 402388 152454
rect 402336 152390 402388 152396
rect 379290 150146 379342 150152
rect 379302 149940 379330 150146
rect 379946 149940 379974 150198
rect 380590 149940 380618 150198
rect 381234 149940 381262 150198
rect 381878 149940 381906 150198
rect 382522 149940 382550 150198
rect 383166 149940 383194 150198
rect 383810 149940 383838 150198
rect 384454 149940 384482 150198
rect 385098 149940 385126 150198
rect 385742 149940 385770 150198
rect 386386 149940 386414 150198
rect 387030 149940 387058 150198
rect 387674 149940 387702 150198
rect 388318 149940 388346 150198
rect 388962 149940 388990 150198
rect 389606 149940 389634 150198
rect 390250 149940 390278 150198
rect 390894 149940 390922 150198
rect 391538 149940 391566 150198
rect 392182 149940 392210 150198
rect 392826 149940 392854 150198
rect 393470 149940 393498 150198
rect 394114 149940 394142 150198
rect 394758 149940 394786 150198
rect 394976 150204 395028 150210
rect 395356 150198 395430 150226
rect 394976 150146 395028 150152
rect 395402 149940 395430 150198
rect 396034 150204 396086 150210
rect 396552 150198 396626 150226
rect 397196 150198 397270 150226
rect 397840 150198 397914 150226
rect 398484 150198 398558 150226
rect 399128 150198 399202 150226
rect 399772 150198 399846 150226
rect 400416 150198 400490 150226
rect 401060 150198 401134 150226
rect 396034 150146 396086 150152
rect 396046 149940 396074 150146
rect 396598 149940 396626 150198
rect 397242 149940 397270 150198
rect 397886 149940 397914 150198
rect 398530 149940 398558 150198
rect 399174 149940 399202 150198
rect 399818 149940 399846 150198
rect 400462 149940 400490 150198
rect 401106 149940 401134 150198
rect 401750 150198 401824 150226
rect 402348 150226 402376 152390
rect 402980 151972 403032 151978
rect 402980 151914 403032 151920
rect 402992 150226 403020 151914
rect 402348 150198 402422 150226
rect 402992 150198 403066 150226
rect 403176 150210 403204 155246
rect 403532 153060 403584 153066
rect 403532 153002 403584 153008
rect 403544 151814 403572 153002
rect 403912 152454 403940 159258
rect 404268 159180 404320 159186
rect 404268 159122 404320 159128
rect 403900 152448 403952 152454
rect 403900 152390 403952 152396
rect 404280 151978 404308 159122
rect 404372 152794 404400 163254
rect 404832 163146 404860 163254
rect 404910 163200 404966 164400
rect 405738 163200 405794 164400
rect 406658 163200 406714 164400
rect 407486 163200 407542 164400
rect 407684 163254 408264 163282
rect 404924 163146 404952 163200
rect 404832 163118 404952 163146
rect 404636 159112 404688 159118
rect 404636 159054 404688 159060
rect 404360 152788 404412 152794
rect 404360 152730 404412 152736
rect 404648 152182 404676 159054
rect 405752 158778 405780 163200
rect 406200 159860 406252 159866
rect 406200 159802 406252 159808
rect 405832 159724 405884 159730
rect 405832 159666 405884 159672
rect 405740 158772 405792 158778
rect 405740 158714 405792 158720
rect 405844 153134 405872 159666
rect 405556 153128 405608 153134
rect 405556 153070 405608 153076
rect 405832 153128 405884 153134
rect 405832 153070 405884 153076
rect 404636 152176 404688 152182
rect 404636 152118 404688 152124
rect 404912 152040 404964 152046
rect 404912 151982 404964 151988
rect 404268 151972 404320 151978
rect 404268 151914 404320 151920
rect 403544 151786 403664 151814
rect 403636 150226 403664 151786
rect 404924 150226 404952 151982
rect 405568 150226 405596 153070
rect 406212 150226 406240 159802
rect 406672 153066 406700 163200
rect 407500 159662 407528 163200
rect 407488 159656 407540 159662
rect 407488 159598 407540 159604
rect 406844 154148 406896 154154
rect 406844 154090 406896 154096
rect 406660 153060 406712 153066
rect 406660 153002 406712 153008
rect 406856 150226 406884 154090
rect 407684 152425 407712 163254
rect 408236 163146 408264 163254
rect 408314 163200 408370 164400
rect 409142 163200 409198 164400
rect 409970 163200 410026 164400
rect 410798 163200 410854 164400
rect 411272 163254 411576 163282
rect 408328 163146 408356 163200
rect 408236 163118 408356 163146
rect 408500 159588 408552 159594
rect 408500 159530 408552 159536
rect 407670 152416 407726 152425
rect 407670 152351 407726 152360
rect 408132 152244 408184 152250
rect 408132 152186 408184 152192
rect 407488 152108 407540 152114
rect 407488 152050 407540 152056
rect 407500 150226 407528 152050
rect 408144 150226 408172 152186
rect 408512 152114 408540 159530
rect 409156 158846 409184 163200
rect 409984 160070 410012 163200
rect 409972 160064 410024 160070
rect 409972 160006 410024 160012
rect 410812 159594 410840 163200
rect 410800 159588 410852 159594
rect 410800 159530 410852 159536
rect 409144 158840 409196 158846
rect 409144 158782 409196 158788
rect 410800 158840 410852 158846
rect 410800 158782 410852 158788
rect 409236 158772 409288 158778
rect 409236 158714 409288 158720
rect 408776 153128 408828 153134
rect 408776 153070 408828 153076
rect 408500 152108 408552 152114
rect 408500 152050 408552 152056
rect 408788 150226 408816 153070
rect 409248 152250 409276 158714
rect 409420 154080 409472 154086
rect 409420 154022 409472 154028
rect 409236 152244 409288 152250
rect 409236 152186 409288 152192
rect 409432 150226 409460 154022
rect 410064 153196 410116 153202
rect 410064 153138 410116 153144
rect 410076 150226 410104 153138
rect 410812 153134 410840 158782
rect 410800 153128 410852 153134
rect 410800 153070 410852 153076
rect 411272 152930 411300 163254
rect 411548 163146 411576 163254
rect 411626 163200 411682 164400
rect 412546 163200 412602 164400
rect 413374 163200 413430 164400
rect 414202 163200 414258 164400
rect 414308 163254 414980 163282
rect 411640 163146 411668 163200
rect 411548 163118 411668 163146
rect 411352 159384 411404 159390
rect 411352 159326 411404 159332
rect 410708 152924 410760 152930
rect 410708 152866 410760 152872
rect 411260 152924 411312 152930
rect 411260 152866 411312 152872
rect 410720 150226 410748 152866
rect 411364 150226 411392 159326
rect 412560 158914 412588 163200
rect 412548 158908 412600 158914
rect 412548 158850 412600 158856
rect 412916 158908 412968 158914
rect 412916 158850 412968 158856
rect 411996 154216 412048 154222
rect 411996 154158 412048 154164
rect 412008 150226 412036 154158
rect 412928 153202 412956 158850
rect 413388 158778 413416 163200
rect 413836 159996 413888 160002
rect 413836 159938 413888 159944
rect 413744 159792 413796 159798
rect 413744 159734 413796 159740
rect 413376 158772 413428 158778
rect 413376 158714 413428 158720
rect 412916 153196 412968 153202
rect 412916 153138 412968 153144
rect 412640 152380 412692 152386
rect 412640 152322 412692 152328
rect 412652 150226 412680 152322
rect 413756 152046 413784 159734
rect 413848 152386 413876 159938
rect 414216 159390 414244 163200
rect 414204 159384 414256 159390
rect 414204 159326 414256 159332
rect 414308 152522 414336 163254
rect 414952 163146 414980 163254
rect 415030 163200 415086 164400
rect 415412 163254 415808 163282
rect 415044 163146 415072 163200
rect 414952 163118 415072 163146
rect 414572 154284 414624 154290
rect 414572 154226 414624 154232
rect 413928 152516 413980 152522
rect 413928 152458 413980 152464
rect 414296 152516 414348 152522
rect 414296 152458 414348 152464
rect 413836 152380 413888 152386
rect 413836 152322 413888 152328
rect 413744 152040 413796 152046
rect 413744 151982 413796 151988
rect 413284 151836 413336 151842
rect 413284 151778 413336 151784
rect 413296 150226 413324 151778
rect 413940 150226 413968 152458
rect 414584 150226 414612 154226
rect 415412 152998 415440 163254
rect 415780 163146 415808 163254
rect 415858 163200 415914 164400
rect 416686 163200 416742 164400
rect 417514 163200 417570 164400
rect 418172 163254 418384 163282
rect 415872 163146 415900 163200
rect 415780 163118 415900 163146
rect 416596 159928 416648 159934
rect 416596 159870 416648 159876
rect 415216 152992 415268 152998
rect 415216 152934 415268 152940
rect 415400 152992 415452 152998
rect 415400 152934 415452 152940
rect 415228 150226 415256 152934
rect 415860 152448 415912 152454
rect 415860 152390 415912 152396
rect 415872 150226 415900 152390
rect 416608 152386 416636 159870
rect 416700 158846 416728 163200
rect 417528 159730 417556 163200
rect 417884 160064 417936 160070
rect 417884 160006 417936 160012
rect 417516 159724 417568 159730
rect 417516 159666 417568 159672
rect 416688 158840 416740 158846
rect 416688 158782 416740 158788
rect 417148 154488 417200 154494
rect 417148 154430 417200 154436
rect 416504 152380 416556 152386
rect 416504 152322 416556 152328
rect 416596 152380 416648 152386
rect 416596 152322 416648 152328
rect 416516 150226 416544 152322
rect 417160 150226 417188 154430
rect 417424 152652 417476 152658
rect 417424 152594 417476 152600
rect 417436 151910 417464 152594
rect 417896 152318 417924 160006
rect 418172 152454 418200 163254
rect 418356 163146 418384 163254
rect 418434 163200 418490 164400
rect 418632 163254 419212 163282
rect 418448 163146 418476 163200
rect 418356 163118 418476 163146
rect 418632 152658 418660 163254
rect 419184 163146 419212 163254
rect 419262 163200 419318 164400
rect 420090 163200 420146 164400
rect 420918 163200 420974 164400
rect 421024 163254 421696 163282
rect 419276 163146 419304 163200
rect 419184 163118 419304 163146
rect 420104 158982 420132 163200
rect 420932 159798 420960 163200
rect 420920 159792 420972 159798
rect 420920 159734 420972 159740
rect 420092 158976 420144 158982
rect 420092 158918 420144 158924
rect 419540 158840 419592 158846
rect 419540 158782 419592 158788
rect 418620 152652 418672 152658
rect 418620 152594 418672 152600
rect 419080 152584 419132 152590
rect 419080 152526 419132 152532
rect 418160 152448 418212 152454
rect 418160 152390 418212 152396
rect 417792 152312 417844 152318
rect 417792 152254 417844 152260
rect 417884 152312 417936 152318
rect 417884 152254 417936 152260
rect 417424 151904 417476 151910
rect 417424 151846 417476 151852
rect 417804 150226 417832 152254
rect 418436 151972 418488 151978
rect 418436 151914 418488 151920
rect 418448 150226 418476 151914
rect 419092 150226 419120 152526
rect 419552 152046 419580 158782
rect 419632 158772 419684 158778
rect 419632 158714 419684 158720
rect 419540 152040 419592 152046
rect 419540 151982 419592 151988
rect 419644 151842 419672 158714
rect 419724 154420 419776 154426
rect 419724 154362 419776 154368
rect 419632 151836 419684 151842
rect 419632 151778 419684 151784
rect 419736 150226 419764 154362
rect 421024 152726 421052 163254
rect 421668 163146 421696 163254
rect 421746 163200 421802 164400
rect 422574 163200 422630 164400
rect 423402 163200 423458 164400
rect 424322 163200 424378 164400
rect 425150 163200 425206 164400
rect 425978 163200 426034 164400
rect 426452 163254 426756 163282
rect 421760 163146 421788 163200
rect 421668 163118 421788 163146
rect 422484 154352 422536 154358
rect 422484 154294 422536 154300
rect 420368 152720 420420 152726
rect 420368 152662 420420 152668
rect 421012 152720 421064 152726
rect 421012 152662 421064 152668
rect 420380 150226 420408 152662
rect 421748 152312 421800 152318
rect 421748 152254 421800 152260
rect 421012 152176 421064 152182
rect 421012 152118 421064 152124
rect 421024 150226 421052 152118
rect 421760 151978 421788 152254
rect 421656 151972 421708 151978
rect 421656 151914 421708 151920
rect 421748 151972 421800 151978
rect 421748 151914 421800 151920
rect 421668 150226 421696 151914
rect 422496 151814 422524 154294
rect 422588 152182 422616 163200
rect 423036 153876 423088 153882
rect 423036 153818 423088 153824
rect 422576 152176 422628 152182
rect 422576 152118 422628 152124
rect 422852 151972 422904 151978
rect 422852 151914 422904 151920
rect 422404 151786 422524 151814
rect 422404 150226 422432 151786
rect 422864 151774 422892 151914
rect 422852 151768 422904 151774
rect 422852 151710 422904 151716
rect 423048 150226 423076 153818
rect 423416 152658 423444 163200
rect 424336 159866 424364 163200
rect 424324 159860 424376 159866
rect 424324 159802 424376 159808
rect 424876 159520 424928 159526
rect 424876 159462 424928 159468
rect 423496 158976 423548 158982
rect 423496 158918 423548 158924
rect 423404 152652 423456 152658
rect 423404 152594 423456 152600
rect 423508 151978 423536 158918
rect 423588 152108 423640 152114
rect 423588 152050 423640 152056
rect 423496 151972 423548 151978
rect 423496 151914 423548 151920
rect 401750 149940 401778 150198
rect 402394 149940 402422 150198
rect 403038 149940 403066 150198
rect 403164 150204 403216 150210
rect 403636 150198 403710 150226
rect 403164 150146 403216 150152
rect 403682 149940 403710 150198
rect 404314 150204 404366 150210
rect 404924 150198 404998 150226
rect 405568 150198 405642 150226
rect 406212 150198 406286 150226
rect 406856 150198 406930 150226
rect 407500 150198 407574 150226
rect 408144 150198 408218 150226
rect 408788 150198 408862 150226
rect 409432 150198 409506 150226
rect 410076 150198 410150 150226
rect 410720 150198 410794 150226
rect 411364 150198 411438 150226
rect 412008 150198 412082 150226
rect 412652 150198 412726 150226
rect 413296 150198 413370 150226
rect 413940 150198 414014 150226
rect 414584 150198 414658 150226
rect 415228 150198 415302 150226
rect 415872 150198 415946 150226
rect 416516 150198 416590 150226
rect 417160 150198 417234 150226
rect 417804 150198 417878 150226
rect 418448 150198 418522 150226
rect 419092 150198 419166 150226
rect 419736 150198 419810 150226
rect 420380 150198 420454 150226
rect 421024 150198 421098 150226
rect 421668 150198 421742 150226
rect 404314 150146 404366 150152
rect 404326 149940 404354 150146
rect 404970 149940 404998 150198
rect 405614 149940 405642 150198
rect 406258 149940 406286 150198
rect 406902 149940 406930 150198
rect 407546 149940 407574 150198
rect 408190 149940 408218 150198
rect 408834 149940 408862 150198
rect 409478 149940 409506 150198
rect 410122 149940 410150 150198
rect 410766 149940 410794 150198
rect 411410 149940 411438 150198
rect 412054 149940 412082 150198
rect 412698 149940 412726 150198
rect 413342 149940 413370 150198
rect 413986 149940 414014 150198
rect 414630 149940 414658 150198
rect 415274 149940 415302 150198
rect 415918 149940 415946 150198
rect 416562 149940 416590 150198
rect 417206 149940 417234 150198
rect 417850 149940 417878 150198
rect 418494 149940 418522 150198
rect 419138 149940 419166 150198
rect 419782 149940 419810 150198
rect 420426 149940 420454 150198
rect 421070 149940 421098 150198
rect 421714 149940 421742 150198
rect 422358 150198 422432 150226
rect 423002 150198 423076 150226
rect 423600 150226 423628 152050
rect 424140 151904 424192 151910
rect 424140 151846 424192 151852
rect 424152 151814 424180 151846
rect 424152 151786 424272 151814
rect 424244 150226 424272 151786
rect 424888 150226 424916 159462
rect 425164 152114 425192 163200
rect 425520 153944 425572 153950
rect 425520 153886 425572 153892
rect 425152 152108 425204 152114
rect 425152 152050 425204 152056
rect 425532 150226 425560 153886
rect 425992 152386 426020 163200
rect 426452 152862 426480 163254
rect 426728 163146 426756 163254
rect 426806 163200 426862 164400
rect 427634 163200 427690 164400
rect 427832 163254 428412 163282
rect 426820 163146 426848 163200
rect 426728 163118 426848 163146
rect 427648 159458 427676 163200
rect 427360 159452 427412 159458
rect 427360 159394 427412 159400
rect 427636 159452 427688 159458
rect 427636 159394 427688 159400
rect 426164 152856 426216 152862
rect 426164 152798 426216 152804
rect 426440 152856 426492 152862
rect 426440 152798 426492 152804
rect 425980 152380 426032 152386
rect 425980 152322 426032 152328
rect 426176 150226 426204 152798
rect 427084 152652 427136 152658
rect 427084 152594 427136 152600
rect 427096 152386 427124 152594
rect 427084 152380 427136 152386
rect 427084 152322 427136 152328
rect 426808 152312 426860 152318
rect 426808 152254 426860 152260
rect 426820 150226 426848 152254
rect 427372 150226 427400 159394
rect 427832 152658 427860 163254
rect 428384 163146 428412 163254
rect 428462 163200 428518 164400
rect 429290 163200 429346 164400
rect 429396 163254 430160 163282
rect 428476 163146 428504 163200
rect 428384 163118 428504 163146
rect 429200 153060 429252 153066
rect 429200 153002 429252 153008
rect 428004 152788 428056 152794
rect 428004 152730 428056 152736
rect 427820 152652 427872 152658
rect 427820 152594 427872 152600
rect 428016 150226 428044 152730
rect 428648 152244 428700 152250
rect 428648 152186 428700 152192
rect 428660 150226 428688 152186
rect 429212 151814 429240 153002
rect 429304 152250 429332 163200
rect 429396 152794 429424 163254
rect 430132 163146 430160 163254
rect 430210 163200 430266 164400
rect 430684 163254 430988 163282
rect 430224 163146 430252 163200
rect 430132 163118 430252 163146
rect 429936 159656 429988 159662
rect 429936 159598 429988 159604
rect 429384 152788 429436 152794
rect 429384 152730 429436 152736
rect 429292 152244 429344 152250
rect 429292 152186 429344 152192
rect 429212 151786 429332 151814
rect 429304 150226 429332 151786
rect 429948 150226 429976 159598
rect 430684 153134 430712 163254
rect 430960 163146 430988 163254
rect 431038 163200 431094 164400
rect 431866 163200 431922 164400
rect 431972 163254 432644 163282
rect 431052 163146 431080 163200
rect 430960 163118 431080 163146
rect 430672 153128 430724 153134
rect 430672 153070 430724 153076
rect 431224 153060 431276 153066
rect 431224 153002 431276 153008
rect 430578 152416 430634 152425
rect 430578 152351 430634 152360
rect 430592 150226 430620 152351
rect 431236 150226 431264 153002
rect 431880 152561 431908 163200
rect 431972 153066 432000 163254
rect 432616 163146 432644 163254
rect 432694 163200 432750 164400
rect 433522 163200 433578 164400
rect 434350 163200 434406 164400
rect 434732 163254 435128 163282
rect 432708 163146 432736 163200
rect 432616 163118 432736 163146
rect 432512 159588 432564 159594
rect 432512 159530 432564 159536
rect 431960 153060 432012 153066
rect 431960 153002 432012 153008
rect 431866 152552 431922 152561
rect 431866 152487 431922 152496
rect 431776 151836 431828 151842
rect 431828 151786 431908 151814
rect 431776 151778 431828 151784
rect 431880 150226 431908 151786
rect 432524 150226 432552 159530
rect 433536 152930 433564 163200
rect 434364 153202 434392 163200
rect 433800 153196 433852 153202
rect 433800 153138 433852 153144
rect 434352 153196 434404 153202
rect 434352 153138 434404 153144
rect 433156 152924 433208 152930
rect 433156 152866 433208 152872
rect 433524 152924 433576 152930
rect 433524 152866 433576 152872
rect 433168 150226 433196 152866
rect 433812 150226 433840 153138
rect 434444 151904 434496 151910
rect 434444 151846 434496 151852
rect 434456 150226 434484 151846
rect 434732 151842 434760 163254
rect 435100 163146 435128 163254
rect 435178 163200 435234 164400
rect 436098 163200 436154 164400
rect 436204 163254 436876 163282
rect 435192 163146 435220 163200
rect 435100 163118 435220 163146
rect 435088 159384 435140 159390
rect 435088 159326 435140 159332
rect 434720 151836 434772 151842
rect 434720 151778 434772 151784
rect 435100 150226 435128 159326
rect 435364 152720 435416 152726
rect 435364 152662 435416 152668
rect 435376 151910 435404 152662
rect 435468 152658 435680 152674
rect 435456 152652 435692 152658
rect 435508 152646 435640 152652
rect 435456 152594 435508 152600
rect 435640 152594 435692 152600
rect 435732 152516 435784 152522
rect 435732 152458 435784 152464
rect 435364 151904 435416 151910
rect 435364 151846 435416 151852
rect 435744 150226 435772 152458
rect 436112 152454 436140 163200
rect 436204 152590 436232 163254
rect 436848 163146 436876 163254
rect 436926 163200 436982 164400
rect 437754 163200 437810 164400
rect 438582 163200 438638 164400
rect 438872 163254 439360 163282
rect 436940 163146 436968 163200
rect 436848 163118 436968 163146
rect 437664 159724 437716 159730
rect 437664 159666 437716 159672
rect 436376 152992 436428 152998
rect 436376 152934 436428 152940
rect 436192 152584 436244 152590
rect 436192 152526 436244 152532
rect 436100 152448 436152 152454
rect 436100 152390 436152 152396
rect 436388 150226 436416 152934
rect 437112 152448 437164 152454
rect 437112 152390 437164 152396
rect 437124 152046 437152 152390
rect 437020 152040 437072 152046
rect 437020 151982 437072 151988
rect 437112 152040 437164 152046
rect 437112 151982 437164 151988
rect 437032 150226 437060 151982
rect 437676 150226 437704 159666
rect 437768 152454 437796 163200
rect 438308 152516 438360 152522
rect 438308 152458 438360 152464
rect 438400 152516 438452 152522
rect 438400 152458 438452 152464
rect 437756 152448 437808 152454
rect 437756 152390 437808 152396
rect 438320 150226 438348 152458
rect 438412 151910 438440 152458
rect 438596 151910 438624 163200
rect 438872 152998 438900 163254
rect 439332 163146 439360 163254
rect 439410 163200 439466 164400
rect 440238 163200 440294 164400
rect 440344 163254 441016 163282
rect 439424 163146 439452 163200
rect 439332 163118 439452 163146
rect 438860 152992 438912 152998
rect 438860 152934 438912 152940
rect 440252 152726 440280 163200
rect 438952 152720 439004 152726
rect 438952 152662 439004 152668
rect 440240 152720 440292 152726
rect 440240 152662 440292 152668
rect 438400 151904 438452 151910
rect 438400 151846 438452 151852
rect 438584 151904 438636 151910
rect 438584 151846 438636 151852
rect 438964 150226 438992 152662
rect 440344 152046 440372 163254
rect 440988 163146 441016 163254
rect 441066 163200 441122 164400
rect 441986 163200 442042 164400
rect 442814 163200 442870 164400
rect 443012 163254 443592 163282
rect 441080 163146 441108 163200
rect 440988 163118 441108 163146
rect 442000 161474 442028 163200
rect 441908 161446 442028 161474
rect 440424 159792 440476 159798
rect 440424 159734 440476 159740
rect 440240 152040 440292 152046
rect 440240 151982 440292 151988
rect 440332 152040 440384 152046
rect 440332 151982 440384 151988
rect 439596 151972 439648 151978
rect 439596 151914 439648 151920
rect 439608 150226 439636 151914
rect 440252 151842 440280 151982
rect 440056 151836 440108 151842
rect 440240 151836 440292 151842
rect 440108 151796 440188 151824
rect 440056 151778 440108 151784
rect 440160 151706 440188 151796
rect 440436 151814 440464 159734
rect 441620 153196 441672 153202
rect 441620 153138 441672 153144
rect 441712 153196 441764 153202
rect 441712 153138 441764 153144
rect 441632 152726 441660 153138
rect 441724 153066 441752 153138
rect 441712 153060 441764 153066
rect 441712 153002 441764 153008
rect 441804 153060 441856 153066
rect 441804 153002 441856 153008
rect 441816 152946 441844 153002
rect 441724 152930 441844 152946
rect 441908 152930 441936 161446
rect 442724 159860 442776 159866
rect 442724 159802 442776 159808
rect 441712 152924 441844 152930
rect 441764 152918 441844 152924
rect 441896 152924 441948 152930
rect 441712 152866 441764 152872
rect 441896 152866 441948 152872
rect 440516 152720 440568 152726
rect 440516 152662 440568 152668
rect 441620 152720 441672 152726
rect 441620 152662 441672 152668
rect 440528 151978 440556 152662
rect 440884 152516 440936 152522
rect 440884 152458 440936 152464
rect 442080 152516 442132 152522
rect 442080 152458 442132 152464
rect 440516 151972 440568 151978
rect 440516 151914 440568 151920
rect 440240 151778 440292 151784
rect 440344 151786 440464 151814
rect 440148 151700 440200 151706
rect 440148 151642 440200 151648
rect 440344 150226 440372 151786
rect 423600 150198 423674 150226
rect 424244 150198 424318 150226
rect 424888 150198 424962 150226
rect 425532 150198 425606 150226
rect 426176 150198 426250 150226
rect 426820 150198 426894 150226
rect 427372 150198 427446 150226
rect 428016 150198 428090 150226
rect 428660 150198 428734 150226
rect 429304 150198 429378 150226
rect 429948 150198 430022 150226
rect 430592 150198 430666 150226
rect 431236 150198 431310 150226
rect 431880 150198 431954 150226
rect 432524 150198 432598 150226
rect 433168 150198 433242 150226
rect 433812 150198 433886 150226
rect 434456 150198 434530 150226
rect 435100 150198 435174 150226
rect 435744 150198 435818 150226
rect 436388 150198 436462 150226
rect 437032 150198 437106 150226
rect 437676 150198 437750 150226
rect 438320 150198 438394 150226
rect 438964 150198 439038 150226
rect 439608 150198 439682 150226
rect 422358 149940 422386 150198
rect 423002 149940 423030 150198
rect 423646 149940 423674 150198
rect 424290 149940 424318 150198
rect 424934 149940 424962 150198
rect 425578 149940 425606 150198
rect 426222 149940 426250 150198
rect 426866 149940 426894 150198
rect 427418 149940 427446 150198
rect 428062 149940 428090 150198
rect 428706 149940 428734 150198
rect 429350 149940 429378 150198
rect 429994 149940 430022 150198
rect 430638 149940 430666 150198
rect 431282 149940 431310 150198
rect 431926 149940 431954 150198
rect 432570 149940 432598 150198
rect 433214 149940 433242 150198
rect 433858 149940 433886 150198
rect 434502 149940 434530 150198
rect 435146 149940 435174 150198
rect 435790 149940 435818 150198
rect 436434 149940 436462 150198
rect 437078 149940 437106 150198
rect 437722 149940 437750 150198
rect 438366 149940 438394 150198
rect 439010 149940 439038 150198
rect 439654 149940 439682 150198
rect 440298 150198 440372 150226
rect 440896 150226 440924 152458
rect 442092 152250 442120 152458
rect 442172 152380 442224 152386
rect 442172 152322 442224 152328
rect 442080 152244 442132 152250
rect 442080 152186 442132 152192
rect 441528 152176 441580 152182
rect 441528 152118 441580 152124
rect 441540 150226 441568 152118
rect 442184 150226 442212 152322
rect 442736 151814 442764 159802
rect 442828 152386 442856 163200
rect 443012 153202 443040 163254
rect 443564 163146 443592 163254
rect 443642 163200 443698 164400
rect 444470 163200 444526 164400
rect 445298 163200 445354 164400
rect 446126 163200 446182 164400
rect 446324 163254 446904 163282
rect 443656 163146 443684 163200
rect 443564 163118 443684 163146
rect 443000 153196 443052 153202
rect 443000 153138 443052 153144
rect 444196 153196 444248 153202
rect 444196 153138 444248 153144
rect 442816 152380 442868 152386
rect 442816 152322 442868 152328
rect 444208 152318 444236 153138
rect 444104 152312 444156 152318
rect 444104 152254 444156 152260
rect 444196 152312 444248 152318
rect 444196 152254 444248 152260
rect 443460 152244 443512 152250
rect 443460 152186 443512 152192
rect 442736 151786 442856 151814
rect 442828 150226 442856 151786
rect 443472 150226 443500 152186
rect 443736 152040 443788 152046
rect 443564 151988 443736 151994
rect 443564 151982 443788 151988
rect 443564 151966 443776 151982
rect 443564 151910 443592 151966
rect 443552 151904 443604 151910
rect 443552 151846 443604 151852
rect 444116 150226 444144 152254
rect 444484 152114 444512 163200
rect 444748 152856 444800 152862
rect 444748 152798 444800 152804
rect 444472 152108 444524 152114
rect 444472 152050 444524 152056
rect 444760 150226 444788 152798
rect 445312 152726 445340 163200
rect 445392 159452 445444 159458
rect 445392 159394 445444 159400
rect 445208 152720 445260 152726
rect 445208 152662 445260 152668
rect 445300 152720 445352 152726
rect 445300 152662 445352 152668
rect 445220 152250 445248 152662
rect 445208 152244 445260 152250
rect 445208 152186 445260 152192
rect 445404 150226 445432 159394
rect 446140 158982 446168 163200
rect 446128 158976 446180 158982
rect 446128 158918 446180 158924
rect 446324 152862 446352 163254
rect 446876 163146 446904 163254
rect 446954 163200 447010 164400
rect 447874 163200 447930 164400
rect 448702 163200 448758 164400
rect 449530 163200 449586 164400
rect 450358 163200 450414 164400
rect 451186 163200 451242 164400
rect 452014 163200 452070 164400
rect 452842 163200 452898 164400
rect 453762 163200 453818 164400
rect 454590 163200 454646 164400
rect 455418 163200 455474 164400
rect 456246 163200 456302 164400
rect 457074 163200 457130 164400
rect 457902 163200 457958 164400
rect 458730 163200 458786 164400
rect 459650 163200 459706 164400
rect 460478 163200 460534 164400
rect 461306 163200 461362 164400
rect 462134 163200 462190 164400
rect 462962 163200 463018 164400
rect 463790 163200 463846 164400
rect 464618 163200 464674 164400
rect 465538 163200 465594 164400
rect 466366 163200 466422 164400
rect 467194 163200 467250 164400
rect 468022 163200 468078 164400
rect 468850 163200 468906 164400
rect 469678 163200 469734 164400
rect 470506 163200 470562 164400
rect 471426 163200 471482 164400
rect 472254 163200 472310 164400
rect 473082 163200 473138 164400
rect 473910 163200 473966 164400
rect 474738 163200 474794 164400
rect 475566 163200 475622 164400
rect 476394 163200 476450 164400
rect 477314 163200 477370 164400
rect 478142 163200 478198 164400
rect 478970 163200 479026 164400
rect 479798 163200 479854 164400
rect 480626 163200 480682 164400
rect 481454 163200 481510 164400
rect 482282 163200 482338 164400
rect 483202 163200 483258 164400
rect 484030 163200 484086 164400
rect 484412 163254 484808 163282
rect 446968 163146 446996 163200
rect 446876 163118 446996 163146
rect 447888 159390 447916 163200
rect 448716 159526 448744 163200
rect 449544 160002 449572 163200
rect 449532 159996 449584 160002
rect 449532 159938 449584 159944
rect 450372 159866 450400 163200
rect 450360 159860 450412 159866
rect 450360 159802 450412 159808
rect 448704 159520 448756 159526
rect 448704 159462 448756 159468
rect 451200 159458 451228 163200
rect 451188 159452 451240 159458
rect 451188 159394 451240 159400
rect 447876 159384 447928 159390
rect 447876 159326 447928 159332
rect 452028 159118 452056 163200
rect 452016 159112 452068 159118
rect 452016 159054 452068 159060
rect 452856 158846 452884 163200
rect 452844 158840 452896 158846
rect 452844 158782 452896 158788
rect 453776 158778 453804 163200
rect 453948 158976 454000 158982
rect 453948 158918 454000 158924
rect 453764 158772 453816 158778
rect 453764 158714 453816 158720
rect 453960 153202 453988 158918
rect 454604 158914 454632 163200
rect 455432 159050 455460 163200
rect 456156 159996 456208 160002
rect 456156 159938 456208 159944
rect 456064 159520 456116 159526
rect 456064 159462 456116 159468
rect 455420 159044 455472 159050
rect 455420 158986 455472 158992
rect 454592 158908 454644 158914
rect 454592 158850 454644 158856
rect 449256 153196 449308 153202
rect 449256 153138 449308 153144
rect 453948 153196 454000 153202
rect 453948 153138 454000 153144
rect 447968 153128 448020 153134
rect 447968 153070 448020 153076
rect 446956 152924 447008 152930
rect 446956 152866 447008 152872
rect 446312 152856 446364 152862
rect 446312 152798 446364 152804
rect 446036 152652 446088 152658
rect 446036 152594 446088 152600
rect 446048 150226 446076 152594
rect 446680 152516 446732 152522
rect 446680 152458 446732 152464
rect 446772 152516 446824 152522
rect 446772 152458 446824 152464
rect 446692 150226 446720 152458
rect 446784 152386 446812 152458
rect 446772 152380 446824 152386
rect 446772 152322 446824 152328
rect 446968 152318 446996 152866
rect 447324 152788 447376 152794
rect 447324 152730 447376 152736
rect 446956 152312 447008 152318
rect 446956 152254 447008 152260
rect 447336 150226 447364 152730
rect 447980 150226 448008 153070
rect 448610 152552 448666 152561
rect 448610 152487 448666 152496
rect 448624 150226 448652 152487
rect 449268 150226 449296 153138
rect 449900 153060 449952 153066
rect 449900 153002 449952 153008
rect 449912 150226 449940 153002
rect 454408 152992 454460 152998
rect 454408 152934 454460 152940
rect 452476 152584 452528 152590
rect 452476 152526 452528 152532
rect 450544 152244 450596 152250
rect 450544 152186 450596 152192
rect 450556 150226 450584 152186
rect 451832 151904 451884 151910
rect 451832 151846 451884 151852
rect 451096 151836 451148 151842
rect 451148 151786 451228 151814
rect 451096 151778 451148 151784
rect 451200 150226 451228 151786
rect 451844 150226 451872 151846
rect 452488 150226 452516 152526
rect 453120 152448 453172 152454
rect 453120 152390 453172 152396
rect 453132 150226 453160 152390
rect 453764 152040 453816 152046
rect 453764 151982 453816 151988
rect 453776 150226 453804 151982
rect 454420 150226 454448 152934
rect 455696 152176 455748 152182
rect 455696 152118 455748 152124
rect 455052 151972 455104 151978
rect 455052 151914 455104 151920
rect 455064 150226 455092 151914
rect 455708 150226 455736 152118
rect 456076 151978 456104 159462
rect 456064 151972 456116 151978
rect 456064 151914 456116 151920
rect 456168 151842 456196 159938
rect 456260 158982 456288 163200
rect 457088 160002 457116 163200
rect 457076 159996 457128 160002
rect 457076 159938 457128 159944
rect 456892 159860 456944 159866
rect 456892 159802 456944 159808
rect 456800 159452 456852 159458
rect 456800 159394 456852 159400
rect 456248 158976 456300 158982
rect 456248 158918 456300 158924
rect 456812 152930 456840 159394
rect 456800 152924 456852 152930
rect 456800 152866 456852 152872
rect 456340 152312 456392 152318
rect 456340 152254 456392 152260
rect 456156 151836 456208 151842
rect 456156 151778 456208 151784
rect 456352 150226 456380 152254
rect 456904 152046 456932 159802
rect 457916 159526 457944 163200
rect 458744 159866 458772 163200
rect 458732 159860 458784 159866
rect 458732 159802 458784 159808
rect 457904 159520 457956 159526
rect 457904 159462 457956 159468
rect 459664 159458 459692 163200
rect 459652 159452 459704 159458
rect 459652 159394 459704 159400
rect 456984 159384 457036 159390
rect 456984 159326 457036 159332
rect 456996 153134 457024 159326
rect 460492 159322 460520 163200
rect 460480 159316 460532 159322
rect 460480 159258 460532 159264
rect 461320 159186 461348 163200
rect 461308 159180 461360 159186
rect 461308 159122 461360 159128
rect 462148 159118 462176 163200
rect 458180 159112 458232 159118
rect 458180 159054 458232 159060
rect 462136 159112 462188 159118
rect 462136 159054 462188 159060
rect 456984 153128 457036 153134
rect 456984 153070 457036 153076
rect 458192 152522 458220 159054
rect 462228 158908 462280 158914
rect 462228 158850 462280 158856
rect 459652 158840 459704 158846
rect 459652 158782 459704 158788
rect 459560 158772 459612 158778
rect 459560 158714 459612 158720
rect 459468 153196 459520 153202
rect 459468 153138 459520 153144
rect 458916 152720 458968 152726
rect 458916 152662 458968 152668
rect 456984 152516 457036 152522
rect 456984 152458 457036 152464
rect 458180 152516 458232 152522
rect 458180 152458 458232 152464
rect 456892 152040 456944 152046
rect 456892 151982 456944 151988
rect 456996 150226 457024 152458
rect 457628 152380 457680 152386
rect 457628 152322 457680 152328
rect 457640 150226 457668 152322
rect 458180 152108 458232 152114
rect 458180 152050 458232 152056
rect 458192 150226 458220 152050
rect 458928 150226 458956 152662
rect 440896 150198 440970 150226
rect 441540 150198 441614 150226
rect 442184 150198 442258 150226
rect 442828 150198 442902 150226
rect 443472 150198 443546 150226
rect 444116 150198 444190 150226
rect 444760 150198 444834 150226
rect 445404 150198 445478 150226
rect 446048 150198 446122 150226
rect 446692 150198 446766 150226
rect 447336 150198 447410 150226
rect 447980 150198 448054 150226
rect 448624 150198 448698 150226
rect 449268 150198 449342 150226
rect 449912 150198 449986 150226
rect 450556 150198 450630 150226
rect 451200 150198 451274 150226
rect 451844 150198 451918 150226
rect 452488 150198 452562 150226
rect 453132 150198 453206 150226
rect 453776 150198 453850 150226
rect 454420 150198 454494 150226
rect 455064 150198 455138 150226
rect 455708 150198 455782 150226
rect 456352 150198 456426 150226
rect 456996 150198 457070 150226
rect 457640 150198 457714 150226
rect 458192 150198 458266 150226
rect 440298 149940 440326 150198
rect 440942 149940 440970 150198
rect 441586 149940 441614 150198
rect 442230 149940 442258 150198
rect 442874 149940 442902 150198
rect 443518 149940 443546 150198
rect 444162 149940 444190 150198
rect 444806 149940 444834 150198
rect 445450 149940 445478 150198
rect 446094 149940 446122 150198
rect 446738 149940 446766 150198
rect 447382 149940 447410 150198
rect 448026 149940 448054 150198
rect 448670 149940 448698 150198
rect 449314 149940 449342 150198
rect 449958 149940 449986 150198
rect 450602 149940 450630 150198
rect 451246 149940 451274 150198
rect 451890 149940 451918 150198
rect 452534 149940 452562 150198
rect 453178 149940 453206 150198
rect 453822 149940 453850 150198
rect 454466 149940 454494 150198
rect 455110 149940 455138 150198
rect 455754 149940 455782 150198
rect 456398 149940 456426 150198
rect 457042 149940 457070 150198
rect 457686 149940 457714 150198
rect 458238 149940 458266 150198
rect 458882 150198 458956 150226
rect 459480 150226 459508 153138
rect 459572 152590 459600 158714
rect 459664 152726 459692 158782
rect 462240 153202 462268 158850
rect 462976 158778 463004 163200
rect 463516 159044 463568 159050
rect 463516 158986 463568 158992
rect 462964 158772 463016 158778
rect 462964 158714 463016 158720
rect 462228 153196 462280 153202
rect 462228 153138 462280 153144
rect 463528 153134 463556 158986
rect 463608 158976 463660 158982
rect 463608 158918 463660 158924
rect 460756 153128 460808 153134
rect 460756 153070 460808 153076
rect 463516 153128 463568 153134
rect 463516 153070 463568 153076
rect 460112 152856 460164 152862
rect 460112 152798 460164 152804
rect 459652 152720 459704 152726
rect 459652 152662 459704 152668
rect 459560 152584 459612 152590
rect 459560 152526 459612 152532
rect 460124 150226 460152 152798
rect 460768 150226 460796 153070
rect 463620 153066 463648 158918
rect 463804 158846 463832 163200
rect 463884 159996 463936 160002
rect 463884 159938 463936 159944
rect 463792 158840 463844 158846
rect 463792 158782 463844 158788
rect 463608 153060 463660 153066
rect 463608 153002 463660 153008
rect 463332 152924 463384 152930
rect 463332 152866 463384 152872
rect 462688 152040 462740 152046
rect 462688 151982 462740 151988
rect 461400 151972 461452 151978
rect 461400 151914 461452 151920
rect 461412 150226 461440 151914
rect 462044 151836 462096 151842
rect 462044 151778 462096 151784
rect 462056 150226 462084 151778
rect 462700 150226 462728 151982
rect 463344 150226 463372 152866
rect 463896 151842 463924 159938
rect 464632 158982 464660 163200
rect 465080 159860 465132 159866
rect 465080 159802 465132 159808
rect 464712 159520 464764 159526
rect 464712 159462 464764 159468
rect 464620 158976 464672 158982
rect 464620 158918 464672 158924
rect 464724 152998 464752 159462
rect 464712 152992 464764 152998
rect 464712 152934 464764 152940
rect 465092 152930 465120 159802
rect 465552 159050 465580 163200
rect 465540 159044 465592 159050
rect 465540 158986 465592 158992
rect 466380 158914 466408 163200
rect 467208 159594 467236 163200
rect 468036 159866 468064 163200
rect 468024 159860 468076 159866
rect 468024 159802 468076 159808
rect 467196 159588 467248 159594
rect 467196 159530 467248 159536
rect 468864 159458 468892 163200
rect 469692 160002 469720 163200
rect 469680 159996 469732 160002
rect 469680 159938 469732 159944
rect 466460 159452 466512 159458
rect 466460 159394 466512 159400
rect 468852 159452 468904 159458
rect 468852 159394 468904 159400
rect 466368 158908 466420 158914
rect 466368 158850 466420 158856
rect 466472 153202 466500 159394
rect 470520 159390 470548 163200
rect 470508 159384 470560 159390
rect 470508 159326 470560 159332
rect 466644 159316 466696 159322
rect 466644 159258 466696 159264
rect 465908 153196 465960 153202
rect 465908 153138 465960 153144
rect 466460 153196 466512 153202
rect 466460 153138 466512 153144
rect 465080 152924 465132 152930
rect 465080 152866 465132 152872
rect 464620 152720 464672 152726
rect 464620 152662 464672 152668
rect 463976 152516 464028 152522
rect 463976 152458 464028 152464
rect 463884 151836 463936 151842
rect 463884 151778 463936 151784
rect 463988 150226 464016 152458
rect 464632 150226 464660 152662
rect 465264 152584 465316 152590
rect 465264 152526 465316 152532
rect 465276 150226 465304 152526
rect 465920 150226 465948 153138
rect 466656 153134 466684 159258
rect 467840 159180 467892 159186
rect 467840 159122 467892 159128
rect 466552 153128 466604 153134
rect 466552 153070 466604 153076
rect 466644 153128 466696 153134
rect 466644 153070 466696 153076
rect 466564 150226 466592 153070
rect 467288 153060 467340 153066
rect 467288 153002 467340 153008
rect 467300 150226 467328 153002
rect 467852 151910 467880 159122
rect 471440 159118 471468 163200
rect 472268 159186 472296 163200
rect 472256 159180 472308 159186
rect 472256 159122 472308 159128
rect 467932 159112 467984 159118
rect 467932 159054 467984 159060
rect 471428 159112 471480 159118
rect 471428 159054 471480 159060
rect 467840 151904 467892 151910
rect 467840 151846 467892 151852
rect 467944 151842 467972 159054
rect 472532 159044 472584 159050
rect 472532 158986 472584 158992
rect 471428 158976 471480 158982
rect 471428 158918 471480 158924
rect 471336 158840 471388 158846
rect 471336 158782 471388 158788
rect 469220 158772 469272 158778
rect 469220 158714 469272 158720
rect 468392 152992 468444 152998
rect 468392 152934 468444 152940
rect 467748 151836 467800 151842
rect 467932 151836 467984 151842
rect 467800 151786 467880 151814
rect 467748 151778 467800 151784
rect 459480 150198 459554 150226
rect 460124 150198 460198 150226
rect 460768 150198 460842 150226
rect 461412 150198 461486 150226
rect 462056 150198 462130 150226
rect 462700 150198 462774 150226
rect 463344 150198 463418 150226
rect 463988 150198 464062 150226
rect 464632 150198 464706 150226
rect 465276 150198 465350 150226
rect 465920 150198 465994 150226
rect 466564 150198 466638 150226
rect 458882 149940 458910 150198
rect 459526 149940 459554 150198
rect 460170 149940 460198 150198
rect 460814 149940 460842 150198
rect 461458 149940 461486 150198
rect 462102 149940 462130 150198
rect 462746 149940 462774 150198
rect 463390 149940 463418 150198
rect 464034 149940 464062 150198
rect 464678 149940 464706 150198
rect 465322 149940 465350 150198
rect 465966 149940 465994 150198
rect 466610 149940 466638 150198
rect 467254 150198 467328 150226
rect 467852 150226 467880 151786
rect 468404 151814 468432 152934
rect 469128 152924 469180 152930
rect 469128 152866 469180 152872
rect 468404 151786 468524 151814
rect 467932 151778 467984 151784
rect 468496 150226 468524 151786
rect 469140 150226 469168 152866
rect 469232 151978 469260 158714
rect 471348 153202 471376 158782
rect 469772 153196 469824 153202
rect 469772 153138 469824 153144
rect 471336 153196 471388 153202
rect 471336 153138 471388 153144
rect 469220 151972 469272 151978
rect 469220 151914 469272 151920
rect 469784 150226 469812 153138
rect 471440 153134 471468 158918
rect 472440 158908 472492 158914
rect 472440 158850 472492 158856
rect 470416 153128 470468 153134
rect 470416 153070 470468 153076
rect 471428 153128 471480 153134
rect 471428 153070 471480 153076
rect 470428 150226 470456 153070
rect 472452 153066 472480 158850
rect 472440 153060 472492 153066
rect 472440 153002 472492 153008
rect 472544 152998 472572 158986
rect 473096 158778 473124 163200
rect 473360 159588 473412 159594
rect 473360 159530 473412 159536
rect 473084 158772 473136 158778
rect 473084 158714 473136 158720
rect 473372 153202 473400 159530
rect 473924 159050 473952 163200
rect 473912 159044 473964 159050
rect 473912 158986 473964 158992
rect 474752 158846 474780 163200
rect 474832 159452 474884 159458
rect 474832 159394 474884 159400
rect 474740 158840 474792 158846
rect 474740 158782 474792 158788
rect 472992 153196 473044 153202
rect 472992 153138 473044 153144
rect 473360 153196 473412 153202
rect 473360 153138 473412 153144
rect 472532 152992 472584 152998
rect 472532 152934 472584 152940
rect 472348 151972 472400 151978
rect 472348 151914 472400 151920
rect 471060 151904 471112 151910
rect 471060 151846 471112 151852
rect 471072 150226 471100 151846
rect 471704 151836 471756 151842
rect 471704 151778 471756 151784
rect 471716 150226 471744 151778
rect 472360 150226 472388 151914
rect 473004 150226 473032 153138
rect 474844 153134 474872 159394
rect 475580 158982 475608 163200
rect 476028 159860 476080 159866
rect 476028 159802 476080 159808
rect 475568 158976 475620 158982
rect 475568 158918 475620 158924
rect 475568 153196 475620 153202
rect 475568 153138 475620 153144
rect 473636 153128 473688 153134
rect 473636 153070 473688 153076
rect 474832 153128 474884 153134
rect 474832 153070 474884 153076
rect 473648 150226 473676 153070
rect 474924 153060 474976 153066
rect 474924 153002 474976 153008
rect 474280 152992 474332 152998
rect 474280 152934 474332 152940
rect 474292 150226 474320 152934
rect 474936 150226 474964 153002
rect 475580 150226 475608 153138
rect 476040 151814 476068 159802
rect 476120 159384 476172 159390
rect 476120 159326 476172 159332
rect 476132 153202 476160 159326
rect 476408 158914 476436 163200
rect 477328 159458 477356 163200
rect 477408 159996 477460 160002
rect 477408 159938 477460 159944
rect 477316 159452 477368 159458
rect 477316 159394 477368 159400
rect 476396 158908 476448 158914
rect 476396 158850 476448 158856
rect 476120 153196 476172 153202
rect 476120 153138 476172 153144
rect 476856 153128 476908 153134
rect 476856 153070 476908 153076
rect 476040 151786 476252 151814
rect 476224 150226 476252 151786
rect 476868 150226 476896 153070
rect 477420 151814 477448 159938
rect 478156 159390 478184 163200
rect 478984 159662 479012 163200
rect 479812 159866 479840 163200
rect 480640 159934 480668 163200
rect 480628 159928 480680 159934
rect 480628 159870 480680 159876
rect 479800 159860 479852 159866
rect 479800 159802 479852 159808
rect 478972 159656 479024 159662
rect 478972 159598 479024 159604
rect 478144 159384 478196 159390
rect 478144 159326 478196 159332
rect 479432 159180 479484 159186
rect 479432 159122 479484 159128
rect 477684 159112 477736 159118
rect 477684 159054 477736 159060
rect 477420 151786 477540 151814
rect 477512 150226 477540 151786
rect 467852 150198 467926 150226
rect 468496 150198 468570 150226
rect 469140 150198 469214 150226
rect 469784 150198 469858 150226
rect 470428 150198 470502 150226
rect 471072 150198 471146 150226
rect 471716 150198 471790 150226
rect 472360 150198 472434 150226
rect 473004 150198 473078 150226
rect 473648 150198 473722 150226
rect 474292 150198 474366 150226
rect 474936 150198 475010 150226
rect 475580 150198 475654 150226
rect 476224 150198 476298 150226
rect 476868 150198 476942 150226
rect 477512 150198 477586 150226
rect 477696 150210 477724 159054
rect 478972 158772 479024 158778
rect 478972 158714 479024 158720
rect 478144 153196 478196 153202
rect 478144 153138 478196 153144
rect 478156 150226 478184 153138
rect 467254 149940 467282 150198
rect 467898 149940 467926 150198
rect 468542 149940 468570 150198
rect 469186 149940 469214 150198
rect 469830 149940 469858 150198
rect 470474 149940 470502 150198
rect 471118 149940 471146 150198
rect 471762 149940 471790 150198
rect 472406 149940 472434 150198
rect 473050 149940 473078 150198
rect 473694 149940 473722 150198
rect 474338 149940 474366 150198
rect 474982 149940 475010 150198
rect 475626 149940 475654 150198
rect 476270 149940 476298 150198
rect 476914 149940 476942 150198
rect 477558 149940 477586 150198
rect 477684 150204 477736 150210
rect 478156 150198 478230 150226
rect 478984 150210 479012 158714
rect 479444 150226 479472 159122
rect 480720 159044 480772 159050
rect 480720 158986 480772 158992
rect 480260 158840 480312 158846
rect 480260 158782 480312 158788
rect 477684 150146 477736 150152
rect 478202 149940 478230 150198
rect 478834 150204 478886 150210
rect 478834 150146 478886 150152
rect 478972 150204 479024 150210
rect 479444 150198 479518 150226
rect 480272 150210 480300 158782
rect 480732 150226 480760 158986
rect 481468 158778 481496 163200
rect 481640 158976 481692 158982
rect 481640 158918 481692 158924
rect 481456 158772 481508 158778
rect 481456 158714 481508 158720
rect 481652 151814 481680 158918
rect 482296 158846 482324 163200
rect 483216 161474 483244 163200
rect 483124 161446 483244 161474
rect 482652 158908 482704 158914
rect 482652 158850 482704 158856
rect 482284 158840 482336 158846
rect 482284 158782 482336 158788
rect 481652 151786 482048 151814
rect 482020 150226 482048 151786
rect 482664 150226 482692 158850
rect 483124 152998 483152 161446
rect 483296 159452 483348 159458
rect 483296 159394 483348 159400
rect 483204 159384 483256 159390
rect 483204 159326 483256 159332
rect 483112 152992 483164 152998
rect 483112 152934 483164 152940
rect 478972 150146 479024 150152
rect 478846 149940 478874 150146
rect 479490 149940 479518 150198
rect 480122 150204 480174 150210
rect 480122 150146 480174 150152
rect 480260 150204 480312 150210
rect 480732 150198 480806 150226
rect 480260 150146 480312 150152
rect 480134 149940 480162 150146
rect 480778 149940 480806 150198
rect 481410 150204 481462 150210
rect 482020 150198 482094 150226
rect 482664 150198 482738 150226
rect 483216 150210 483244 159326
rect 483308 150226 483336 159394
rect 484044 153202 484072 163200
rect 484032 153196 484084 153202
rect 484032 153138 484084 153144
rect 484412 153066 484440 163254
rect 484780 163146 484808 163254
rect 484858 163200 484914 164400
rect 484964 163254 485636 163282
rect 484872 163146 484900 163200
rect 484780 163118 484900 163146
rect 484584 159656 484636 159662
rect 484584 159598 484636 159604
rect 484400 153060 484452 153066
rect 484400 153002 484452 153008
rect 484596 150226 484624 159598
rect 484964 153134 484992 163254
rect 485608 163146 485636 163254
rect 485686 163200 485742 164400
rect 485792 163254 486464 163282
rect 485700 163146 485728 163200
rect 485608 163118 485728 163146
rect 485228 159860 485280 159866
rect 485228 159802 485280 159808
rect 484952 153128 485004 153134
rect 484952 153070 485004 153076
rect 485240 150226 485268 159802
rect 485792 152046 485820 163254
rect 486436 163146 486464 163254
rect 486514 163200 486570 164400
rect 487342 163200 487398 164400
rect 488170 163200 488226 164400
rect 488552 163254 489040 163282
rect 486528 163146 486556 163200
rect 486436 163118 486556 163146
rect 485964 159928 486016 159934
rect 485964 159870 486016 159876
rect 485780 152040 485832 152046
rect 485780 151982 485832 151988
rect 485976 150226 486004 159870
rect 487252 158840 487304 158846
rect 487252 158782 487304 158788
rect 486516 158772 486568 158778
rect 486516 158714 486568 158720
rect 481410 150146 481462 150152
rect 481422 149940 481450 150146
rect 482066 149940 482094 150198
rect 482710 149940 482738 150198
rect 483204 150204 483256 150210
rect 483308 150198 483382 150226
rect 483204 150146 483256 150152
rect 483354 149940 483382 150198
rect 483986 150204 484038 150210
rect 484596 150198 484670 150226
rect 485240 150198 485314 150226
rect 483986 150146 484038 150152
rect 483998 149940 484026 150146
rect 484642 149940 484670 150198
rect 485286 149940 485314 150198
rect 485930 150198 486004 150226
rect 486528 150226 486556 158714
rect 487264 150226 487292 158782
rect 487356 151978 487384 163200
rect 487804 152992 487856 152998
rect 487804 152934 487856 152940
rect 487344 151972 487396 151978
rect 487344 151914 487396 151920
rect 486528 150198 486602 150226
rect 485930 149940 485958 150198
rect 486574 149940 486602 150198
rect 487218 150198 487292 150226
rect 487816 150226 487844 152934
rect 488184 151842 488212 163200
rect 488448 153196 488500 153202
rect 488448 153138 488500 153144
rect 488172 151836 488224 151842
rect 488172 151778 488224 151784
rect 488460 150226 488488 153138
rect 488552 151910 488580 163254
rect 489012 163146 489040 163254
rect 489090 163200 489146 164400
rect 489918 163200 489974 164400
rect 490024 163254 490696 163282
rect 489104 163146 489132 163200
rect 489012 163118 489132 163146
rect 489932 153202 489960 163200
rect 489920 153196 489972 153202
rect 489920 153138 489972 153144
rect 489644 153128 489696 153134
rect 489644 153070 489696 153076
rect 489000 153060 489052 153066
rect 489000 153002 489052 153008
rect 488540 151904 488592 151910
rect 488540 151846 488592 151852
rect 489012 150226 489040 153002
rect 489656 150226 489684 153070
rect 490024 152930 490052 163254
rect 490668 163146 490696 163254
rect 490746 163200 490802 164400
rect 491312 163254 491524 163282
rect 490760 163146 490788 163200
rect 490668 163118 490788 163146
rect 491312 152998 491340 163254
rect 491496 163146 491524 163254
rect 491574 163200 491630 164400
rect 491680 163254 492352 163282
rect 491588 163146 491616 163200
rect 491496 163118 491616 163146
rect 491680 153134 491708 163254
rect 492324 163146 492352 163254
rect 492402 163200 492458 164400
rect 492692 163254 493180 163282
rect 492416 163146 492444 163200
rect 492324 163118 492444 163146
rect 491668 153128 491720 153134
rect 491668 153070 491720 153076
rect 492692 153066 492720 163254
rect 493152 163146 493180 163254
rect 493230 163200 493286 164400
rect 494058 163200 494114 164400
rect 494978 163200 495034 164400
rect 495544 163254 495756 163282
rect 493244 163146 493272 163200
rect 493152 163118 493272 163146
rect 494072 153202 494100 163200
rect 492864 153196 492916 153202
rect 492864 153138 492916 153144
rect 494060 153196 494112 153202
rect 494060 153138 494112 153144
rect 492680 153060 492732 153066
rect 492680 153002 492732 153008
rect 491300 152992 491352 152998
rect 491300 152934 491352 152940
rect 490012 152924 490064 152930
rect 490012 152866 490064 152872
rect 490288 152040 490340 152046
rect 490288 151982 490340 151988
rect 490300 150226 490328 151982
rect 490932 151972 490984 151978
rect 490932 151914 490984 151920
rect 490944 150226 490972 151914
rect 492220 151904 492272 151910
rect 492220 151846 492272 151852
rect 491576 151836 491628 151842
rect 491576 151778 491628 151784
rect 491588 150226 491616 151778
rect 492232 150226 492260 151846
rect 492876 150226 492904 153138
rect 494992 153134 495020 163200
rect 494796 153128 494848 153134
rect 494796 153070 494848 153076
rect 494980 153128 495032 153134
rect 494980 153070 495032 153076
rect 494152 152992 494204 152998
rect 494152 152934 494204 152940
rect 493508 152924 493560 152930
rect 493508 152866 493560 152872
rect 493520 150226 493548 152866
rect 494164 150226 494192 152934
rect 494808 150226 494836 153070
rect 495544 153066 495572 163254
rect 495728 163146 495756 163254
rect 495806 163200 495862 164400
rect 496634 163200 496690 164400
rect 496832 163254 497412 163282
rect 495820 163146 495848 163200
rect 495728 163118 495848 163146
rect 496648 153202 496676 163200
rect 496084 153196 496136 153202
rect 496084 153138 496136 153144
rect 496636 153196 496688 153202
rect 496636 153138 496688 153144
rect 495440 153060 495492 153066
rect 495440 153002 495492 153008
rect 495532 153060 495584 153066
rect 495532 153002 495584 153008
rect 495452 150226 495480 153002
rect 496096 150226 496124 153138
rect 496832 153134 496860 163254
rect 497384 163146 497412 163254
rect 497462 163200 497518 164400
rect 498290 163200 498346 164400
rect 499118 163200 499174 164400
rect 499946 163200 500002 164400
rect 500052 163254 500632 163282
rect 497476 163146 497504 163200
rect 497384 163118 497504 163146
rect 498304 156670 498332 163200
rect 498292 156664 498344 156670
rect 498292 156606 498344 156612
rect 498016 153196 498068 153202
rect 498016 153138 498068 153144
rect 496728 153128 496780 153134
rect 496728 153070 496780 153076
rect 496820 153128 496872 153134
rect 496820 153070 496872 153076
rect 496740 150226 496768 153070
rect 497372 153060 497424 153066
rect 497372 153002 497424 153008
rect 497384 150226 497412 153002
rect 498028 150226 498056 153138
rect 498660 153128 498712 153134
rect 498660 153070 498712 153076
rect 498672 150226 498700 153070
rect 499132 151842 499160 163200
rect 499960 163146 499988 163200
rect 500052 163146 500080 163254
rect 499960 163118 500080 163146
rect 499304 156664 499356 156670
rect 499304 156606 499356 156612
rect 499120 151836 499172 151842
rect 499120 151778 499172 151784
rect 499316 150226 499344 156606
rect 499948 151836 500000 151842
rect 499948 151778 500000 151784
rect 499960 150226 499988 151778
rect 500604 150226 500632 163254
rect 500866 163200 500922 164400
rect 501694 163200 501750 164400
rect 502522 163200 502578 164400
rect 503350 163200 503406 164400
rect 503824 163254 504128 163282
rect 500880 151814 500908 163200
rect 501708 161474 501736 163200
rect 501708 161446 501920 161474
rect 500880 151786 501276 151814
rect 501248 150226 501276 151786
rect 501892 150226 501920 161446
rect 502340 156664 502392 156670
rect 502340 156606 502392 156612
rect 487816 150198 487890 150226
rect 488460 150198 488534 150226
rect 489012 150198 489086 150226
rect 489656 150198 489730 150226
rect 490300 150198 490374 150226
rect 490944 150198 491018 150226
rect 491588 150198 491662 150226
rect 492232 150198 492306 150226
rect 492876 150198 492950 150226
rect 493520 150198 493594 150226
rect 494164 150198 494238 150226
rect 494808 150198 494882 150226
rect 495452 150198 495526 150226
rect 496096 150198 496170 150226
rect 496740 150198 496814 150226
rect 497384 150198 497458 150226
rect 498028 150198 498102 150226
rect 498672 150198 498746 150226
rect 499316 150198 499390 150226
rect 499960 150198 500034 150226
rect 500604 150198 500678 150226
rect 501248 150198 501322 150226
rect 501892 150198 501966 150226
rect 502352 150210 502380 156606
rect 502536 150226 502564 163200
rect 503364 156670 503392 163200
rect 503352 156664 503404 156670
rect 503352 156606 503404 156612
rect 503824 150226 503852 163254
rect 504100 163146 504128 163254
rect 504178 163200 504234 164400
rect 504468 163254 504956 163282
rect 504192 163146 504220 163200
rect 504100 163118 504220 163146
rect 504468 150226 504496 163254
rect 504928 163146 504956 163254
rect 505006 163200 505062 164400
rect 505112 163254 505784 163282
rect 505020 163146 505048 163200
rect 504928 163118 505048 163146
rect 505112 150226 505140 163254
rect 505756 163146 505784 163254
rect 505834 163200 505890 164400
rect 506754 163200 506810 164400
rect 507582 163200 507638 164400
rect 508410 163200 508466 164400
rect 509238 163200 509294 164400
rect 509344 163254 509556 163282
rect 505848 163146 505876 163200
rect 505756 163118 505876 163146
rect 506388 158840 506440 158846
rect 506388 158782 506440 158788
rect 505284 158772 505336 158778
rect 505284 158714 505336 158720
rect 505296 151814 505324 158714
rect 505296 151786 505784 151814
rect 505756 150226 505784 151786
rect 506400 150226 506428 158782
rect 506768 158778 506796 163200
rect 507596 158846 507624 163200
rect 508320 158908 508372 158914
rect 508320 158850 508372 158856
rect 507584 158840 507636 158846
rect 507584 158782 507636 158788
rect 506756 158772 506808 158778
rect 506756 158714 506808 158720
rect 507032 158772 507084 158778
rect 507032 158714 507084 158720
rect 507044 150226 507072 158714
rect 507768 151904 507820 151910
rect 507768 151846 507820 151852
rect 507780 150226 507808 151846
rect 487218 149940 487246 150198
rect 487862 149940 487890 150198
rect 488506 149940 488534 150198
rect 489058 149940 489086 150198
rect 489702 149940 489730 150198
rect 490346 149940 490374 150198
rect 490990 149940 491018 150198
rect 491634 149940 491662 150198
rect 492278 149940 492306 150198
rect 492922 149940 492950 150198
rect 493566 149940 493594 150198
rect 494210 149940 494238 150198
rect 494854 149940 494882 150198
rect 495498 149940 495526 150198
rect 496142 149940 496170 150198
rect 496786 149940 496814 150198
rect 497430 149940 497458 150198
rect 498074 149940 498102 150198
rect 498718 149940 498746 150198
rect 499362 149940 499390 150198
rect 500006 149940 500034 150198
rect 500650 149940 500678 150198
rect 501294 149940 501322 150198
rect 501938 149940 501966 150198
rect 502340 150204 502392 150210
rect 502536 150198 502610 150226
rect 502340 150146 502392 150152
rect 502582 149940 502610 150198
rect 503214 150204 503266 150210
rect 503824 150198 503898 150226
rect 504468 150198 504542 150226
rect 505112 150198 505186 150226
rect 505756 150198 505830 150226
rect 506400 150198 506474 150226
rect 507044 150198 507118 150226
rect 503214 150146 503266 150152
rect 503226 149940 503254 150146
rect 503870 149940 503898 150198
rect 504514 149940 504542 150198
rect 505158 149940 505186 150198
rect 505802 149940 505830 150198
rect 506446 149940 506474 150198
rect 507090 149940 507118 150198
rect 507734 150198 507808 150226
rect 508332 150226 508360 158850
rect 508424 158778 508452 163200
rect 509252 163146 509280 163200
rect 509344 163146 509372 163254
rect 509252 163118 509372 163146
rect 508412 158772 508464 158778
rect 508412 158714 508464 158720
rect 509424 158772 509476 158778
rect 509424 158714 509476 158720
rect 509056 151972 509108 151978
rect 509056 151914 509108 151920
rect 509068 150226 509096 151914
rect 509436 151814 509464 158714
rect 509528 151910 509556 163254
rect 510066 163200 510122 164400
rect 510894 163200 510950 164400
rect 511722 163200 511778 164400
rect 512012 163254 512592 163282
rect 510080 158914 510108 163200
rect 510068 158908 510120 158914
rect 510068 158850 510120 158856
rect 510344 152856 510396 152862
rect 510344 152798 510396 152804
rect 509516 151904 509568 151910
rect 509516 151846 509568 151852
rect 509436 151786 509648 151814
rect 508332 150198 508406 150226
rect 507734 149940 507762 150198
rect 508378 149940 508406 150198
rect 509022 150198 509096 150226
rect 509620 150226 509648 151786
rect 510356 150226 510384 152798
rect 510908 151978 510936 163200
rect 511736 158778 511764 163200
rect 511724 158772 511776 158778
rect 511724 158714 511776 158720
rect 510988 153128 511040 153134
rect 510988 153070 511040 153076
rect 510896 151972 510948 151978
rect 510896 151914 510948 151920
rect 511000 150226 511028 153070
rect 511632 153060 511684 153066
rect 511632 153002 511684 153008
rect 511644 150226 511672 153002
rect 512012 152862 512040 163254
rect 512564 163146 512592 163254
rect 512642 163200 512698 164400
rect 513470 163200 513526 164400
rect 514298 163200 514354 164400
rect 514864 163254 515076 163282
rect 512656 163146 512684 163200
rect 512564 163118 512684 163146
rect 512276 153196 512328 153202
rect 512276 153138 512328 153144
rect 512000 152856 512052 152862
rect 512000 152798 512052 152804
rect 512288 150226 512316 153138
rect 513484 153134 513512 163200
rect 513472 153128 513524 153134
rect 513472 153070 513524 153076
rect 513564 153128 513616 153134
rect 513564 153070 513616 153076
rect 512920 152992 512972 152998
rect 512920 152934 512972 152940
rect 512932 150226 512960 152934
rect 513576 150226 513604 153070
rect 514312 153066 514340 163200
rect 514864 153202 514892 163254
rect 515048 163146 515076 163254
rect 515126 163200 515182 164400
rect 515954 163200 516010 164400
rect 516152 163254 516732 163282
rect 515140 163146 515168 163200
rect 515048 163118 515168 163146
rect 514944 158772 514996 158778
rect 514944 158714 514996 158720
rect 514852 153196 514904 153202
rect 514852 153138 514904 153144
rect 514300 153060 514352 153066
rect 514300 153002 514352 153008
rect 514208 152924 514260 152930
rect 514208 152866 514260 152872
rect 514220 150226 514248 152866
rect 514956 151814 514984 158714
rect 515968 152998 515996 163200
rect 516152 153134 516180 163254
rect 516704 163146 516732 163254
rect 516782 163200 516838 164400
rect 517610 163200 517666 164400
rect 518530 163200 518586 164400
rect 518912 163254 519308 163282
rect 516796 163146 516824 163200
rect 516704 163118 516824 163146
rect 517624 161474 517652 163200
rect 517532 161446 517652 161474
rect 517532 158794 517560 161446
rect 517440 158766 517560 158794
rect 518544 158778 518572 163200
rect 518808 159452 518860 159458
rect 518808 159394 518860 159400
rect 518716 159384 518768 159390
rect 518716 159326 518768 159332
rect 518532 158772 518584 158778
rect 516140 153128 516192 153134
rect 516140 153070 516192 153076
rect 515956 152992 516008 152998
rect 515956 152934 516008 152940
rect 517440 152930 517468 158766
rect 518532 158714 518584 158720
rect 517428 152924 517480 152930
rect 517428 152866 517480 152872
rect 516692 152108 516744 152114
rect 516692 152050 516744 152056
rect 516048 151904 516100 151910
rect 516048 151846 516100 151852
rect 514864 151786 514984 151814
rect 515496 151836 515548 151842
rect 514864 150226 514892 151786
rect 515496 151778 515548 151784
rect 515508 150226 515536 151778
rect 509620 150198 509694 150226
rect 509022 149940 509050 150198
rect 509666 149940 509694 150198
rect 510310 150198 510384 150226
rect 510954 150198 511028 150226
rect 511598 150198 511672 150226
rect 512242 150198 512316 150226
rect 512886 150198 512960 150226
rect 513530 150198 513604 150226
rect 514174 150198 514248 150226
rect 514818 150198 514892 150226
rect 515462 150198 515536 150226
rect 516060 150226 516088 151846
rect 516704 150226 516732 152050
rect 517428 151972 517480 151978
rect 517428 151914 517480 151920
rect 517440 150226 517468 151914
rect 518728 150226 518756 159326
rect 516060 150198 516134 150226
rect 516704 150198 516778 150226
rect 510310 149940 510338 150198
rect 510954 149940 510982 150198
rect 511598 149940 511626 150198
rect 512242 149940 512270 150198
rect 512886 149940 512914 150198
rect 513530 149940 513558 150198
rect 514174 149940 514202 150198
rect 514818 149940 514846 150198
rect 515462 149940 515490 150198
rect 516106 149940 516134 150198
rect 516750 149940 516778 150198
rect 517394 150198 517468 150226
rect 518026 150204 518078 150210
rect 517394 149940 517422 150198
rect 518026 150146 518078 150152
rect 518682 150198 518756 150226
rect 518820 150210 518848 159394
rect 518912 151842 518940 163254
rect 519280 163146 519308 163254
rect 519358 163200 519414 164400
rect 519464 163254 520136 163282
rect 519372 163146 519400 163200
rect 519280 163118 519400 163146
rect 519358 154184 519414 154193
rect 519358 154119 519414 154128
rect 518900 151836 518952 151842
rect 519372 151814 519400 154119
rect 519464 151910 519492 163254
rect 519726 163160 519782 163169
rect 520108 163146 520136 163254
rect 520186 163200 520242 164400
rect 520292 163254 520964 163282
rect 520200 163146 520228 163200
rect 520108 163118 520228 163146
rect 519726 163095 519782 163104
rect 519542 161664 519598 161673
rect 519542 161599 519598 161608
rect 519452 151904 519504 151910
rect 519452 151846 519504 151852
rect 519372 151786 519492 151814
rect 518900 151778 518952 151784
rect 518808 150204 518860 150210
rect 518038 149940 518066 150146
rect 518682 149940 518710 150198
rect 518808 150146 518860 150152
rect 519464 141137 519492 151786
rect 519556 147937 519584 161599
rect 519634 160168 519690 160177
rect 519634 160103 519690 160112
rect 519542 147928 519598 147937
rect 519542 147863 519598 147872
rect 519648 146577 519676 160103
rect 519740 149297 519768 163095
rect 520186 158672 520242 158681
rect 520186 158607 520242 158616
rect 520002 157176 520058 157185
rect 520002 157111 520058 157120
rect 519818 151192 519874 151201
rect 519818 151127 519874 151136
rect 519726 149288 519782 149297
rect 519726 149223 519782 149232
rect 519726 148200 519782 148209
rect 519726 148135 519782 148144
rect 519634 146568 519690 146577
rect 519634 146503 519690 146512
rect 519634 145208 519690 145217
rect 519634 145143 519690 145152
rect 519542 142216 519598 142225
rect 519542 142151 519598 142160
rect 519450 141128 519506 141137
rect 519450 141063 519506 141072
rect 519266 140584 519322 140593
rect 519266 140519 519322 140528
rect 117240 132518 117360 132546
rect 117332 132410 117360 132518
rect 117240 132382 117360 132410
rect 117240 127945 117268 132382
rect 519280 128897 519308 140519
rect 519358 139088 519414 139097
rect 519358 139023 519414 139032
rect 519266 128888 519322 128897
rect 519266 128823 519322 128832
rect 117226 127936 117282 127945
rect 117226 127871 117282 127880
rect 519372 127537 519400 139023
rect 519450 133104 519506 133113
rect 519450 133039 519506 133048
rect 519358 127528 519414 127537
rect 519358 127463 519414 127472
rect 519358 124128 519414 124137
rect 519358 124063 519414 124072
rect 519266 122632 519322 122641
rect 519266 122567 519322 122576
rect 519280 112577 519308 122567
rect 519372 113937 519400 124063
rect 519464 122097 519492 133039
rect 519556 130257 519584 142151
rect 519648 132977 519676 145143
rect 519740 135697 519768 148135
rect 519832 138417 519860 151127
rect 519910 149696 519966 149705
rect 519910 149631 519966 149640
rect 519818 138408 519874 138417
rect 519818 138343 519874 138352
rect 519924 137057 519952 149631
rect 520016 143857 520044 157111
rect 520094 155680 520150 155689
rect 520094 155615 520150 155624
rect 520002 143848 520058 143857
rect 520002 143783 520058 143792
rect 520108 142497 520136 155615
rect 520200 145353 520228 158607
rect 520292 152114 520320 163254
rect 520936 163146 520964 163254
rect 521014 163200 521070 164400
rect 521842 163200 521898 164400
rect 522670 163200 522726 164400
rect 523498 163200 523554 164400
rect 521028 163146 521056 163200
rect 520936 163118 521056 163146
rect 521856 161474 521884 163200
rect 521672 161446 521884 161474
rect 521672 158794 521700 161446
rect 522684 159458 522712 163200
rect 522672 159452 522724 159458
rect 522672 159394 522724 159400
rect 523512 159390 523540 163200
rect 523500 159384 523552 159390
rect 523500 159326 523552 159332
rect 521580 158766 521700 158794
rect 521014 152688 521070 152697
rect 521014 152623 521070 152632
rect 520280 152108 520332 152114
rect 520280 152050 520332 152056
rect 520186 145344 520242 145353
rect 520186 145279 520242 145288
rect 520922 143712 520978 143721
rect 520922 143647 520978 143656
rect 520094 142488 520150 142497
rect 520094 142423 520150 142432
rect 520094 137592 520150 137601
rect 520094 137527 520150 137536
rect 519910 137048 519966 137057
rect 519910 136983 519966 136992
rect 519910 136096 519966 136105
rect 519910 136031 519966 136040
rect 519726 135688 519782 135697
rect 519726 135623 519782 135632
rect 519634 132968 519690 132977
rect 519634 132903 519690 132912
rect 519634 131472 519690 131481
rect 519634 131407 519690 131416
rect 519542 130248 519598 130257
rect 519542 130183 519598 130192
rect 519542 125624 519598 125633
rect 519542 125559 519598 125568
rect 519450 122088 519506 122097
rect 519450 122023 519506 122032
rect 519556 115297 519584 125559
rect 519648 120737 519676 131407
rect 519726 130112 519782 130121
rect 519726 130047 519782 130056
rect 519634 120728 519690 120737
rect 519634 120663 519690 120672
rect 519740 119377 519768 130047
rect 519818 127120 519874 127129
rect 519818 127055 519874 127064
rect 519726 119368 519782 119377
rect 519726 119303 519782 119312
rect 519832 116657 519860 127055
rect 519924 124817 519952 136031
rect 520002 128616 520058 128625
rect 520002 128551 520058 128560
rect 519910 124808 519966 124817
rect 519910 124743 519966 124752
rect 519910 121136 519966 121145
rect 519910 121071 519966 121080
rect 519818 116648 519874 116657
rect 519818 116583 519874 116592
rect 519542 115288 519598 115297
rect 519542 115223 519598 115232
rect 519818 115016 519874 115025
rect 519818 114951 519874 114960
rect 519358 113928 519414 113937
rect 519358 113863 519414 113872
rect 519726 113520 519782 113529
rect 519726 113455 519782 113464
rect 519266 112568 519322 112577
rect 519266 112503 519322 112512
rect 519542 112024 519598 112033
rect 519542 111959 519598 111968
rect 117134 104816 117190 104825
rect 117134 104751 117190 104760
rect 519556 103057 519584 111959
rect 519634 110528 519690 110537
rect 519634 110463 519690 110472
rect 519542 103048 519598 103057
rect 519542 102983 519598 102992
rect 519648 101697 519676 110463
rect 519740 104417 519768 113455
rect 519832 105777 519860 114951
rect 519924 111217 519952 121071
rect 520016 118017 520044 128551
rect 520108 126177 520136 137527
rect 520186 134600 520242 134609
rect 520186 134535 520242 134544
rect 520094 126168 520150 126177
rect 520094 126103 520150 126112
rect 520200 123457 520228 134535
rect 520936 131617 520964 143647
rect 521028 139777 521056 152623
rect 521580 151978 521608 158766
rect 521568 151972 521620 151978
rect 521568 151914 521620 151920
rect 521106 146704 521162 146713
rect 521106 146639 521162 146648
rect 521014 139768 521070 139777
rect 521014 139703 521070 139712
rect 521120 134337 521148 146639
rect 521106 134328 521162 134337
rect 521106 134263 521162 134272
rect 520922 131608 520978 131617
rect 520922 131543 520978 131552
rect 520186 123448 520242 123457
rect 520186 123383 520242 123392
rect 520094 119640 520150 119649
rect 520094 119575 520150 119584
rect 520002 118008 520058 118017
rect 520002 117943 520058 117952
rect 520002 116512 520058 116521
rect 520002 116447 520058 116456
rect 519910 111208 519966 111217
rect 519910 111143 519966 111152
rect 520016 107137 520044 116447
rect 520108 109857 520136 119575
rect 520186 118144 520242 118153
rect 520186 118079 520242 118088
rect 520094 109848 520150 109857
rect 520094 109783 520150 109792
rect 520200 108497 520228 118079
rect 520922 109032 520978 109041
rect 520922 108967 520978 108976
rect 520186 108488 520242 108497
rect 520186 108423 520242 108432
rect 520002 107128 520058 107137
rect 520002 107063 520058 107072
rect 520278 106040 520334 106049
rect 520278 105975 520334 105984
rect 519818 105768 519874 105777
rect 519818 105703 519874 105712
rect 519726 104408 519782 104417
rect 519726 104343 519782 104352
rect 519634 101688 519690 101697
rect 519634 101623 519690 101632
rect 117042 101008 117098 101017
rect 117042 100943 117098 100952
rect 116858 99104 116914 99113
rect 116858 99039 116914 99048
rect 520292 97617 520320 105975
rect 520830 104544 520886 104553
rect 520830 104479 520886 104488
rect 520738 103048 520794 103057
rect 520738 102983 520794 102992
rect 520278 97608 520334 97617
rect 520278 97543 520334 97552
rect 116766 97200 116822 97209
rect 116766 97135 116822 97144
rect 520278 95568 520334 95577
rect 520278 95503 520334 95512
rect 116674 95296 116730 95305
rect 116674 95231 116730 95240
rect 116582 93392 116638 93401
rect 116582 93327 116638 93336
rect 116124 92472 116176 92478
rect 116124 92414 116176 92420
rect 520186 92440 520242 92449
rect 116136 91361 116164 92414
rect 520186 92375 520242 92384
rect 116122 91352 116178 91361
rect 116122 91287 116178 91296
rect 520002 90944 520058 90953
rect 520002 90879 520058 90888
rect 116124 89684 116176 89690
rect 116124 89626 116176 89632
rect 116136 89457 116164 89626
rect 116122 89448 116178 89457
rect 116122 89383 116178 89392
rect 519634 89448 519690 89457
rect 519634 89383 519690 89392
rect 116032 88324 116084 88330
rect 116032 88266 116084 88272
rect 116044 87553 116072 88266
rect 116030 87544 116086 87553
rect 116030 87479 116086 87488
rect 519082 86456 519138 86465
rect 519082 86391 519138 86400
rect 115202 85640 115258 85649
rect 115202 85575 115258 85584
rect 116584 83972 116636 83978
rect 116584 83914 116636 83920
rect 116596 83745 116624 83914
rect 116582 83736 116638 83745
rect 116582 83671 116638 83680
rect 116216 82816 116268 82822
rect 116216 82758 116268 82764
rect 116228 81841 116256 82758
rect 116214 81832 116270 81841
rect 116214 81767 116270 81776
rect 115940 80028 115992 80034
rect 115940 79970 115992 79976
rect 115952 79937 115980 79970
rect 519096 79937 519124 86391
rect 519648 82657 519676 89383
rect 519910 87952 519966 87961
rect 519910 87887 519966 87896
rect 519818 84960 519874 84969
rect 519818 84895 519874 84904
rect 519634 82648 519690 82657
rect 519634 82583 519690 82592
rect 519726 81968 519782 81977
rect 519726 81903 519782 81912
rect 115938 79928 115994 79937
rect 115938 79863 115994 79872
rect 519082 79928 519138 79937
rect 519082 79863 519138 79872
rect 519634 78976 519690 78985
rect 519634 78911 519690 78920
rect 114192 78668 114244 78674
rect 114192 78610 114244 78616
rect 116124 78668 116176 78674
rect 116124 78610 116176 78616
rect 116136 78033 116164 78610
rect 116122 78024 116178 78033
rect 116122 77959 116178 77968
rect 116674 74080 116730 74089
rect 116674 74015 116730 74024
rect 116582 72176 116638 72185
rect 116582 72111 116638 72120
rect 116596 71806 116624 72111
rect 114192 71800 114244 71806
rect 114192 71742 114244 71748
rect 116584 71800 116636 71806
rect 116584 71742 116636 71748
rect 114100 69080 114152 69086
rect 114100 69022 114152 69028
rect 114008 67652 114060 67658
rect 114008 67594 114060 67600
rect 113916 66292 113968 66298
rect 113916 66234 113968 66240
rect 113364 64728 113416 64734
rect 113364 64670 113416 64676
rect 113376 64569 113404 64670
rect 113362 64560 113418 64569
rect 113362 64495 113418 64504
rect 113824 63572 113876 63578
rect 113824 63514 113876 63520
rect 112444 62144 112496 62150
rect 112444 62086 112496 62092
rect 110326 53952 110382 53961
rect 109696 53910 110326 53938
rect 109696 12434 109724 53910
rect 110326 53887 110382 53896
rect 110326 52592 110382 52601
rect 110326 52527 110382 52536
rect 110340 51218 110368 52527
rect 110340 51190 110460 51218
rect 110326 51096 110382 51105
rect 109512 12406 109724 12434
rect 109788 51054 110326 51082
rect 109512 3913 109540 12406
rect 109788 8242 109816 51054
rect 110326 51031 110382 51040
rect 110432 50946 110460 51190
rect 109604 8214 109816 8242
rect 109880 50918 110460 50946
rect 109498 3904 109554 3913
rect 109498 3839 109554 3848
rect 109498 3496 109554 3505
rect 109498 3431 109554 3440
rect 32402 2680 32458 2689
rect 36358 2680 36414 2689
rect 36018 2638 36358 2666
rect 32402 2615 32458 2624
rect 36358 2615 36414 2624
rect 62394 2680 62450 2689
rect 62394 2615 62450 2624
rect 64142 2680 64198 2689
rect 64142 2615 64198 2624
rect 65338 2680 65394 2689
rect 65338 2615 65394 2624
rect 68006 2680 68062 2689
rect 68006 2615 68062 2624
rect 68466 2680 68522 2689
rect 68466 2615 68522 2624
rect 68834 2680 68890 2689
rect 68834 2615 68890 2624
rect 69386 2680 69442 2689
rect 69386 2615 69442 2624
rect 77022 2680 77078 2689
rect 77252 2680 77308 2689
rect 77022 2615 77078 2624
rect 77128 2638 77252 2666
rect 29550 2408 29606 2417
rect 29302 2366 29550 2394
rect 29550 2343 29606 2352
rect 26054 2272 26110 2281
rect 25990 2230 26054 2258
rect 26054 2207 26110 2216
rect 22926 2136 22982 2145
rect 2700 1358 2728 2108
rect 6012 1737 6040 2108
rect 5998 1728 6054 1737
rect 5998 1663 6054 1672
rect 9324 1465 9352 2108
rect 12636 1601 12664 2108
rect 15948 1873 15976 2108
rect 19366 2094 19656 2122
rect 22678 2094 22926 2122
rect 19628 2009 19656 2094
rect 22926 2071 22982 2080
rect 19614 2000 19670 2009
rect 19614 1935 19670 1944
rect 15934 1864 15990 1873
rect 15934 1799 15990 1808
rect 12622 1592 12678 1601
rect 12622 1527 12678 1536
rect 9310 1456 9366 1465
rect 9310 1391 9366 1400
rect 2688 1352 2740 1358
rect 2688 1294 2740 1300
rect 32416 762 32444 2615
rect 33046 2544 33102 2553
rect 32706 2502 33046 2530
rect 33046 2479 33102 2488
rect 39316 1290 39344 2108
rect 42628 1494 42656 2108
rect 42616 1488 42668 1494
rect 42616 1430 42668 1436
rect 46032 1426 46060 2108
rect 46020 1420 46072 1426
rect 46020 1362 46072 1368
rect 39304 1284 39356 1290
rect 39304 1226 39356 1232
rect 49344 1222 49372 2108
rect 49332 1216 49384 1222
rect 49332 1158 49384 1164
rect 52656 1154 52684 2108
rect 52644 1148 52696 1154
rect 52644 1090 52696 1096
rect 55968 1086 55996 2108
rect 59372 1630 59400 2108
rect 62408 1902 62436 2615
rect 62396 1896 62448 1902
rect 62396 1838 62448 1844
rect 62684 1766 62712 2108
rect 64156 1834 64184 2615
rect 65352 1902 65380 2615
rect 65340 1896 65392 1902
rect 65340 1838 65392 1844
rect 64144 1828 64196 1834
rect 64144 1770 64196 1776
rect 62672 1760 62724 1766
rect 62672 1702 62724 1708
rect 59360 1624 59412 1630
rect 59360 1566 59412 1572
rect 55956 1080 56008 1086
rect 55956 1022 56008 1028
rect 65996 1018 66024 2108
rect 68020 1902 68048 2615
rect 68008 1896 68060 1902
rect 68008 1838 68060 1844
rect 68480 1630 68508 2615
rect 68848 1766 68876 2615
rect 68836 1760 68888 1766
rect 68836 1702 68888 1708
rect 69308 1698 69336 2108
rect 69400 1834 69428 2615
rect 69388 1828 69440 1834
rect 69388 1770 69440 1776
rect 69296 1692 69348 1698
rect 69296 1634 69348 1640
rect 68468 1624 68520 1630
rect 68468 1566 68520 1572
rect 72712 1562 72740 2108
rect 72700 1556 72752 1562
rect 72700 1498 72752 1504
rect 65984 1012 66036 1018
rect 65984 954 66036 960
rect 76024 950 76052 2108
rect 77036 1834 77064 2615
rect 77128 1902 77156 2638
rect 77252 2615 77308 2624
rect 77758 2680 77814 2689
rect 77758 2615 77814 2624
rect 79966 2680 80022 2689
rect 79966 2615 80022 2624
rect 80242 2680 80298 2689
rect 80242 2615 80298 2624
rect 80426 2680 80482 2689
rect 80610 2680 80666 2689
rect 80426 2615 80482 2624
rect 80532 2638 80610 2666
rect 77772 1902 77800 2615
rect 77116 1896 77168 1902
rect 77116 1838 77168 1844
rect 77760 1896 77812 1902
rect 77760 1838 77812 1844
rect 77024 1828 77076 1834
rect 77024 1770 77076 1776
rect 79336 1630 79364 2108
rect 79980 1766 80008 2615
rect 79968 1760 80020 1766
rect 79968 1702 80020 1708
rect 79324 1624 79376 1630
rect 79324 1566 79376 1572
rect 80256 1306 80284 2615
rect 80440 1494 80468 2615
rect 80428 1488 80480 1494
rect 80428 1430 80480 1436
rect 80532 1306 80560 2638
rect 80610 2615 80666 2624
rect 80794 2680 80850 2689
rect 93030 2680 93086 2689
rect 92690 2638 93030 2666
rect 80794 2615 80850 2624
rect 93030 2615 93086 2624
rect 94686 2680 94742 2689
rect 94686 2615 94742 2624
rect 96342 2680 96398 2689
rect 96342 2615 96398 2624
rect 100114 2680 100170 2689
rect 100114 2615 100170 2624
rect 101862 2680 101918 2689
rect 103426 2680 103482 2689
rect 101862 2615 101918 2624
rect 102796 2638 103426 2666
rect 80808 1766 80836 2615
rect 94318 2544 94374 2553
rect 94318 2479 94374 2488
rect 94332 2145 94360 2479
rect 94134 2136 94190 2145
rect 82648 1766 82676 2108
rect 86052 1834 86080 2108
rect 89364 1902 89392 2108
rect 94134 2071 94190 2080
rect 94318 2136 94374 2145
rect 94318 2071 94374 2080
rect 89260 1896 89312 1902
rect 89260 1838 89312 1844
rect 89352 1896 89404 1902
rect 89352 1838 89404 1844
rect 85948 1828 86000 1834
rect 85948 1770 86000 1776
rect 86040 1828 86092 1834
rect 86040 1770 86092 1776
rect 80796 1760 80848 1766
rect 80796 1702 80848 1708
rect 82636 1760 82688 1766
rect 82636 1702 82688 1708
rect 85960 1329 85988 1770
rect 80256 1278 80560 1306
rect 85946 1320 86002 1329
rect 85946 1255 86002 1264
rect 76012 944 76064 950
rect 32692 870 32812 898
rect 89272 921 89300 1838
rect 94148 1494 94176 2071
rect 94136 1488 94188 1494
rect 94136 1430 94188 1436
rect 76012 886 76064 892
rect 89258 912 89314 921
rect 32692 762 32720 870
rect 32784 800 32812 870
rect 94700 882 94728 2615
rect 95988 1057 96016 2108
rect 95974 1048 96030 1057
rect 95974 983 96030 992
rect 89258 847 89314 856
rect 94688 876 94740 882
rect 94688 818 94740 824
rect 96356 814 96384 2615
rect 96434 2544 96490 2553
rect 96434 2479 96490 2488
rect 99838 2544 99894 2553
rect 99838 2479 99894 2488
rect 96448 2145 96476 2479
rect 99852 2145 99880 2479
rect 96434 2136 96490 2145
rect 96434 2071 96490 2080
rect 96618 2136 96674 2145
rect 99654 2136 99710 2145
rect 99406 2094 99604 2122
rect 96618 2071 96674 2080
rect 96632 1494 96660 2071
rect 99576 1630 99604 2094
rect 99654 2071 99710 2080
rect 99838 2136 99894 2145
rect 99838 2071 99894 2080
rect 99668 1902 99696 2071
rect 99656 1896 99708 1902
rect 99656 1838 99708 1844
rect 99472 1624 99524 1630
rect 99472 1566 99524 1572
rect 99564 1624 99616 1630
rect 99564 1566 99616 1572
rect 96620 1488 96672 1494
rect 99484 1476 99512 1566
rect 99656 1488 99708 1494
rect 99484 1448 99656 1476
rect 96620 1430 96672 1436
rect 99656 1430 99708 1436
rect 98274 1320 98330 1329
rect 98274 1255 98330 1264
rect 96344 808 96396 814
rect 32416 734 32720 762
rect 32770 -400 32826 800
rect 98288 800 98316 1255
rect 100128 882 100156 2615
rect 101494 2544 101550 2553
rect 101494 2479 101550 2488
rect 100850 2408 100906 2417
rect 101402 2408 101458 2417
rect 100850 2343 100906 2352
rect 101140 2366 101402 2394
rect 100864 2258 100892 2343
rect 101140 2258 101168 2366
rect 101402 2343 101458 2352
rect 100864 2230 101168 2258
rect 100758 2000 100814 2009
rect 101218 2000 101274 2009
rect 100814 1958 101218 1986
rect 100758 1935 100814 1944
rect 101218 1935 101274 1944
rect 101508 921 101536 2479
rect 101494 912 101550 921
rect 100116 876 100168 882
rect 101494 847 101550 856
rect 100116 818 100168 824
rect 101876 814 101904 2615
rect 102704 1698 102732 2108
rect 102600 1692 102652 1698
rect 102600 1634 102652 1640
rect 102692 1692 102744 1698
rect 102692 1634 102744 1640
rect 102612 1578 102640 1634
rect 102796 1578 102824 2638
rect 103426 2615 103482 2624
rect 103610 2680 103666 2689
rect 103610 2615 103666 2624
rect 102612 1550 102824 1578
rect 103624 1476 103652 2615
rect 104162 2544 104218 2553
rect 104162 2479 104218 2488
rect 104176 2145 104204 2479
rect 104162 2136 104218 2145
rect 104162 2071 104218 2080
rect 104346 2136 104402 2145
rect 106030 2094 106228 2122
rect 104346 2071 104402 2080
rect 104360 1902 104388 2071
rect 104348 1896 104400 1902
rect 104532 1896 104584 1902
rect 104348 1838 104400 1844
rect 104452 1856 104532 1884
rect 104072 1760 104124 1766
rect 104452 1714 104480 1856
rect 104532 1838 104584 1844
rect 105728 1896 105780 1902
rect 105728 1838 105780 1844
rect 105820 1896 105872 1902
rect 105820 1838 105872 1844
rect 105912 1896 105964 1902
rect 105912 1838 105964 1844
rect 104124 1708 104480 1714
rect 104072 1702 104480 1708
rect 104084 1686 104480 1702
rect 103348 1448 103652 1476
rect 105740 1476 105768 1838
rect 105832 1698 105860 1838
rect 105820 1692 105872 1698
rect 105820 1634 105872 1640
rect 105924 1630 105952 1838
rect 106200 1698 106228 2094
rect 109328 1902 109356 2108
rect 109224 1896 109276 1902
rect 109224 1838 109276 1844
rect 109316 1896 109368 1902
rect 109316 1838 109368 1844
rect 106188 1692 106240 1698
rect 106188 1634 106240 1640
rect 105912 1624 105964 1630
rect 105912 1566 105964 1572
rect 106004 1624 106056 1630
rect 106004 1566 106056 1572
rect 106016 1476 106044 1566
rect 105740 1448 106044 1476
rect 108212 1488 108264 1494
rect 103348 1329 103376 1448
rect 108212 1430 108264 1436
rect 108304 1488 108356 1494
rect 108304 1430 108356 1436
rect 103440 1366 103928 1394
rect 103334 1320 103390 1329
rect 103334 1255 103390 1264
rect 103440 1193 103468 1366
rect 103900 1193 103928 1366
rect 108224 1329 108252 1430
rect 108210 1320 108266 1329
rect 108210 1255 108266 1264
rect 108316 1193 108344 1430
rect 103426 1184 103482 1193
rect 103426 1119 103482 1128
rect 103886 1184 103942 1193
rect 103886 1119 103942 1128
rect 108302 1184 108358 1193
rect 109236 1170 109264 1838
rect 109512 1737 109540 3431
rect 109604 1834 109632 8214
rect 109880 7970 109908 50918
rect 110326 48376 110382 48385
rect 109696 7942 109908 7970
rect 109972 48334 110326 48362
rect 109696 3641 109724 7942
rect 109682 3632 109738 3641
rect 109682 3567 109738 3576
rect 109866 2816 109922 2825
rect 109866 2751 109922 2760
rect 109592 1828 109644 1834
rect 109592 1770 109644 1776
rect 109498 1728 109554 1737
rect 109498 1663 109554 1672
rect 109880 1442 109908 2751
rect 109972 1766 110000 48334
rect 110326 48311 110382 48320
rect 110326 47152 110382 47161
rect 110326 47087 110382 47096
rect 110340 45554 110368 47087
rect 110064 45526 110368 45554
rect 110064 7562 110092 45526
rect 110326 44296 110382 44305
rect 110156 44254 110326 44282
rect 110156 8242 110184 44254
rect 110326 44231 110382 44240
rect 110326 41440 110382 41449
rect 110326 41375 110382 41384
rect 110340 35894 110368 41375
rect 110248 35866 110368 35894
rect 110248 8378 110276 35866
rect 110326 34640 110382 34649
rect 110326 34575 110382 34584
rect 110340 8514 110368 34575
rect 110340 8486 110736 8514
rect 110326 8392 110382 8401
rect 110248 8350 110326 8378
rect 110326 8327 110382 8336
rect 110510 8392 110566 8401
rect 110510 8327 110566 8336
rect 110156 8214 110368 8242
rect 110064 7534 110184 7562
rect 110156 7426 110184 7534
rect 110156 7398 110276 7426
rect 110248 4026 110276 7398
rect 110340 7290 110368 8214
rect 110340 7262 110460 7290
rect 110156 3998 110276 4026
rect 110050 3904 110106 3913
rect 110050 3839 110106 3848
rect 109960 1760 110012 1766
rect 109960 1702 110012 1708
rect 109788 1414 109908 1442
rect 109788 1306 109816 1414
rect 109604 1278 109816 1306
rect 109604 1170 109632 1278
rect 109236 1142 109632 1170
rect 108302 1119 108358 1128
rect 110064 1057 110092 3839
rect 110156 1630 110184 3998
rect 110234 3904 110290 3913
rect 110234 3839 110290 3848
rect 110248 3505 110276 3839
rect 110234 3496 110290 3505
rect 110234 3431 110290 3440
rect 110144 1624 110196 1630
rect 110144 1566 110196 1572
rect 110432 1329 110460 7262
rect 110524 1562 110552 8327
rect 110602 5672 110658 5681
rect 110602 5607 110658 5616
rect 110616 2825 110644 5607
rect 110708 3233 110736 8486
rect 111062 7984 111118 7993
rect 111062 7919 111118 7928
rect 110694 3224 110750 3233
rect 110694 3159 110750 3168
rect 110602 2816 110658 2825
rect 110602 2751 110658 2760
rect 111076 1970 111104 7919
rect 111706 2952 111762 2961
rect 111706 2887 111708 2896
rect 111760 2887 111762 2896
rect 111708 2858 111760 2864
rect 111800 2848 111852 2854
rect 111800 2790 111852 2796
rect 111064 1964 111116 1970
rect 111064 1906 111116 1912
rect 110512 1556 110564 1562
rect 110512 1498 110564 1504
rect 110418 1320 110474 1329
rect 110418 1255 110474 1264
rect 111812 1086 111840 2790
rect 112456 1766 112484 62086
rect 112536 42832 112588 42838
rect 112536 42774 112588 42780
rect 112444 1760 112496 1766
rect 112444 1702 112496 1708
rect 111800 1080 111852 1086
rect 110050 1048 110106 1057
rect 111800 1022 111852 1028
rect 110050 983 110106 992
rect 112548 950 112576 42774
rect 113836 7721 113864 63514
rect 113928 19009 113956 66234
rect 114020 30433 114048 67594
rect 114112 41857 114140 69022
rect 114204 53145 114232 71742
rect 116306 70272 116362 70281
rect 116306 70207 116362 70216
rect 116320 69086 116348 70207
rect 116308 69080 116360 69086
rect 116308 69022 116360 69028
rect 116122 68368 116178 68377
rect 116122 68303 116178 68312
rect 116136 67658 116164 68303
rect 116124 67652 116176 67658
rect 116124 67594 116176 67600
rect 116582 66464 116638 66473
rect 116582 66399 116638 66408
rect 116596 66298 116624 66399
rect 116584 66292 116636 66298
rect 116584 66234 116636 66240
rect 116688 64874 116716 74015
rect 519648 73273 519676 78911
rect 519740 75993 519768 81903
rect 519832 78577 519860 84895
rect 519924 81297 519952 87887
rect 520016 84017 520044 90879
rect 520200 85377 520228 92375
rect 520292 88097 520320 95503
rect 520752 94897 520780 102983
rect 520844 96257 520872 104479
rect 520936 100337 520964 108967
rect 521106 107536 521162 107545
rect 521106 107471 521162 107480
rect 521014 101552 521070 101561
rect 521014 101487 521070 101496
rect 520922 100328 520978 100337
rect 520922 100263 520978 100272
rect 520922 98560 520978 98569
rect 520922 98495 520978 98504
rect 520830 96248 520886 96257
rect 520830 96183 520886 96192
rect 520738 94888 520794 94897
rect 520738 94823 520794 94832
rect 520936 90817 520964 98495
rect 521028 93537 521056 101487
rect 521120 98977 521148 107471
rect 521198 100056 521254 100065
rect 521198 99991 521254 100000
rect 521106 98968 521162 98977
rect 521106 98903 521162 98912
rect 521106 93936 521162 93945
rect 521106 93871 521162 93880
rect 521014 93528 521070 93537
rect 521014 93463 521070 93472
rect 520922 90808 520978 90817
rect 520922 90743 520978 90752
rect 520278 88088 520334 88097
rect 520278 88023 520334 88032
rect 521120 86737 521148 93871
rect 521212 92177 521240 99991
rect 521382 97064 521438 97073
rect 521382 96999 521438 97008
rect 521198 92168 521254 92177
rect 521198 92103 521254 92112
rect 521396 89593 521424 96999
rect 521382 89584 521438 89593
rect 521382 89519 521438 89528
rect 521106 86728 521162 86737
rect 521106 86663 521162 86672
rect 520186 85368 520242 85377
rect 520186 85303 520242 85312
rect 520002 84008 520058 84017
rect 520002 83943 520058 83952
rect 520186 83464 520242 83473
rect 520186 83399 520242 83408
rect 519910 81288 519966 81297
rect 519910 81223 519966 81232
rect 520002 80472 520058 80481
rect 520002 80407 520058 80416
rect 519818 78568 519874 78577
rect 519818 78503 519874 78512
rect 519910 77480 519966 77489
rect 519910 77415 519966 77424
rect 519726 75984 519782 75993
rect 519726 75919 519782 75928
rect 519634 73264 519690 73273
rect 519634 73199 519690 73208
rect 519924 71913 519952 77415
rect 520016 74633 520044 80407
rect 520200 77217 520228 83399
rect 520186 77208 520242 77217
rect 520186 77143 520242 77152
rect 520186 75984 520242 75993
rect 520186 75919 520242 75928
rect 520002 74624 520058 74633
rect 520002 74559 520058 74568
rect 519910 71904 519966 71913
rect 519910 71839 519966 71848
rect 520200 70553 520228 75919
rect 521014 74488 521070 74497
rect 521014 74423 521070 74432
rect 520922 72992 520978 73001
rect 520922 72927 520978 72936
rect 520186 70544 520242 70553
rect 520186 70479 520242 70488
rect 520936 67833 520964 72927
rect 521028 69193 521056 74423
rect 521198 71496 521254 71505
rect 521198 71431 521254 71440
rect 521106 69864 521162 69873
rect 521106 69799 521162 69808
rect 521014 69184 521070 69193
rect 521014 69119 521070 69128
rect 521014 68368 521070 68377
rect 521014 68303 521070 68312
rect 520922 67824 520978 67833
rect 520922 67759 520978 67768
rect 520462 66872 520518 66881
rect 520462 66807 520518 66816
rect 520370 65376 520426 65385
rect 520370 65311 520426 65320
rect 116596 64846 116716 64874
rect 116596 64734 116624 64846
rect 116584 64728 116636 64734
rect 116584 64670 116636 64676
rect 116214 64560 116270 64569
rect 116214 64495 116270 64504
rect 116228 63578 116256 64495
rect 116216 63572 116268 63578
rect 116216 63514 116268 63520
rect 116122 62656 116178 62665
rect 116122 62591 116178 62600
rect 116136 62150 116164 62591
rect 116124 62144 116176 62150
rect 116124 62086 116176 62092
rect 520384 61033 520412 65311
rect 520476 62393 520504 66807
rect 521028 63753 521056 68303
rect 521120 65113 521148 69799
rect 521212 66473 521240 71431
rect 521198 66464 521254 66473
rect 521198 66399 521254 66408
rect 521106 65104 521162 65113
rect 521106 65039 521162 65048
rect 521106 63880 521162 63889
rect 521106 63815 521162 63824
rect 521014 63744 521070 63753
rect 521014 63679 521070 63688
rect 520462 62384 520518 62393
rect 520462 62319 520518 62328
rect 521014 62384 521070 62393
rect 521014 62319 521070 62328
rect 520370 61024 520426 61033
rect 520370 60959 520426 60968
rect 520738 60888 520794 60897
rect 520738 60823 520794 60832
rect 116582 60616 116638 60625
rect 116582 60551 116638 60560
rect 114190 53136 114246 53145
rect 114190 53071 114246 53080
rect 116122 43344 116178 43353
rect 116122 43279 116178 43288
rect 116136 42838 116164 43279
rect 116124 42832 116176 42838
rect 116124 42774 116176 42780
rect 114098 41848 114154 41857
rect 114098 41783 114154 41792
rect 114006 30424 114062 30433
rect 114006 30359 114062 30368
rect 116490 27976 116546 27985
rect 116490 27911 116546 27920
rect 116306 26072 116362 26081
rect 116306 26007 116362 26016
rect 116214 22264 116270 22273
rect 116214 22199 116270 22208
rect 116030 20360 116086 20369
rect 116030 20295 116086 20304
rect 113914 19000 113970 19009
rect 113914 18935 113970 18944
rect 115938 16416 115994 16425
rect 115938 16351 115994 16360
rect 113822 7712 113878 7721
rect 113822 7647 113878 7656
rect 115952 2281 115980 16351
rect 116044 2553 116072 20295
rect 116122 18456 116178 18465
rect 116122 18391 116178 18400
rect 116030 2544 116086 2553
rect 116030 2479 116086 2488
rect 116136 2417 116164 18391
rect 116228 2689 116256 22199
rect 116320 3641 116348 26007
rect 116398 24168 116454 24177
rect 116398 24103 116454 24112
rect 116306 3632 116362 3641
rect 116306 3567 116362 3576
rect 116306 3088 116362 3097
rect 116306 3023 116362 3032
rect 116214 2680 116270 2689
rect 116214 2615 116270 2624
rect 116122 2408 116178 2417
rect 116122 2343 116178 2352
rect 115938 2272 115994 2281
rect 115938 2207 115994 2216
rect 116320 1358 116348 3023
rect 116308 1352 116360 1358
rect 116308 1294 116360 1300
rect 116412 1290 116440 24103
rect 116504 1426 116532 27911
rect 116596 1698 116624 60551
rect 116766 58712 116822 58721
rect 116766 58647 116822 58656
rect 116674 56808 116730 56817
rect 116674 56743 116730 56752
rect 116688 7954 116716 56743
rect 116780 7993 116808 58647
rect 519910 57896 519966 57905
rect 519910 57831 519966 57840
rect 519818 56400 519874 56409
rect 519818 56335 519874 56344
rect 519082 53408 519138 53417
rect 519082 53343 519138 53352
rect 519096 50153 519124 53343
rect 519832 52873 519860 56335
rect 519924 54233 519952 57831
rect 520752 56953 520780 60823
rect 521028 58313 521056 62319
rect 521120 59673 521148 63815
rect 521106 59664 521162 59673
rect 521106 59599 521162 59608
rect 521106 59392 521162 59401
rect 521106 59327 521162 59336
rect 521014 58304 521070 58313
rect 521014 58239 521070 58248
rect 520738 56944 520794 56953
rect 520738 56879 520794 56888
rect 521120 55593 521148 59327
rect 521106 55584 521162 55593
rect 521106 55519 521162 55528
rect 520186 54904 520242 54913
rect 520186 54839 520242 54848
rect 519910 54224 519966 54233
rect 519910 54159 519966 54168
rect 519818 52864 519874 52873
rect 519818 52799 519874 52808
rect 520094 51912 520150 51921
rect 520094 51847 520150 51856
rect 519082 50144 519138 50153
rect 519082 50079 519138 50088
rect 519082 48920 519138 48929
rect 519082 48855 519138 48864
rect 519096 46073 519124 48855
rect 520108 48793 520136 51847
rect 520200 51513 520228 54839
rect 520186 51504 520242 51513
rect 520186 51439 520242 51448
rect 520186 50416 520242 50425
rect 520186 50351 520242 50360
rect 520094 48784 520150 48793
rect 520094 48719 520150 48728
rect 520200 47433 520228 50351
rect 520186 47424 520242 47433
rect 520186 47359 520242 47368
rect 519910 47288 519966 47297
rect 519910 47223 519966 47232
rect 519082 46064 519138 46073
rect 519082 45999 519138 46008
rect 519726 45792 519782 45801
rect 519726 45727 519782 45736
rect 519740 43353 519768 45727
rect 519924 44713 519952 47223
rect 519910 44704 519966 44713
rect 519910 44639 519966 44648
rect 520186 44296 520242 44305
rect 520186 44231 520242 44240
rect 519726 43344 519782 43353
rect 519726 43279 519782 43288
rect 520200 41993 520228 44231
rect 520738 42800 520794 42809
rect 520738 42735 520794 42744
rect 520186 41984 520242 41993
rect 520186 41919 520242 41928
rect 520752 41313 520780 42735
rect 520738 41304 520794 41313
rect 520738 41239 520794 41248
rect 520922 41304 520978 41313
rect 520922 41239 520978 41248
rect 520936 39953 520964 41239
rect 520922 39944 520978 39953
rect 520922 39879 520978 39888
rect 520922 39808 520978 39817
rect 520922 39743 520978 39752
rect 116950 39536 117006 39545
rect 116950 39471 117006 39480
rect 116858 37632 116914 37641
rect 116858 37567 116914 37576
rect 116766 7984 116822 7993
rect 116676 7948 116728 7954
rect 116872 7954 116900 37567
rect 116766 7919 116822 7928
rect 116860 7948 116912 7954
rect 116676 7890 116728 7896
rect 116860 7890 116912 7896
rect 116964 7834 116992 39471
rect 520936 37913 520964 39743
rect 521106 38312 521162 38321
rect 521106 38247 521162 38256
rect 520922 37904 520978 37913
rect 520922 37839 520978 37848
rect 521120 37233 521148 38247
rect 521106 37224 521162 37233
rect 521106 37159 521162 37168
rect 521566 36816 521622 36825
rect 521566 36751 521622 36760
rect 521580 36009 521608 36751
rect 521566 36000 521622 36009
rect 521566 35935 521622 35944
rect 520922 35320 520978 35329
rect 520922 35255 520978 35264
rect 520936 34513 520964 35255
rect 520922 34504 520978 34513
rect 520922 34439 520978 34448
rect 117134 33824 117190 33833
rect 117134 33759 117190 33768
rect 521106 33824 521162 33833
rect 521106 33759 521162 33768
rect 117042 31784 117098 31793
rect 117042 31719 117098 31728
rect 116688 7806 116992 7834
rect 117056 7818 117084 31719
rect 117044 7812 117096 7818
rect 116688 3233 116716 7806
rect 117044 7754 117096 7760
rect 116860 7744 116912 7750
rect 117148 7698 117176 33759
rect 521120 33153 521148 33759
rect 521106 33144 521162 33153
rect 521106 33079 521162 33088
rect 521106 32328 521162 32337
rect 521106 32263 521162 32272
rect 521120 31657 521148 32263
rect 521106 31648 521162 31657
rect 521106 31583 521162 31592
rect 117226 29880 117282 29889
rect 117226 29815 117282 29824
rect 116860 7686 116912 7692
rect 116768 7676 116820 7682
rect 116768 7618 116820 7624
rect 116674 3224 116730 3233
rect 116674 3159 116730 3168
rect 116584 1692 116636 1698
rect 116584 1634 116636 1640
rect 116492 1420 116544 1426
rect 116492 1362 116544 1368
rect 116400 1284 116452 1290
rect 116400 1226 116452 1232
rect 116780 1222 116808 7618
rect 116768 1216 116820 1222
rect 116768 1158 116820 1164
rect 116872 1018 116900 7686
rect 116964 7670 117176 7698
rect 117240 7682 117268 29815
rect 520922 29336 520978 29345
rect 520922 29271 520978 29280
rect 520936 28393 520964 29271
rect 520922 28384 520978 28393
rect 520922 28319 520978 28328
rect 521106 24848 521162 24857
rect 521106 24783 521162 24792
rect 521120 23633 521148 24783
rect 521106 23624 521162 23633
rect 521106 23559 521162 23568
rect 520370 23216 520426 23225
rect 520370 23151 520426 23160
rect 520384 22273 520412 23151
rect 520370 22264 520426 22273
rect 520370 22199 520426 22208
rect 520922 21720 520978 21729
rect 520922 21655 520978 21664
rect 520936 20913 520964 21655
rect 520922 20904 520978 20913
rect 520922 20839 520978 20848
rect 521106 20224 521162 20233
rect 521106 20159 521162 20168
rect 521120 19553 521148 20159
rect 521106 19544 521162 19553
rect 521106 19479 521162 19488
rect 521106 9344 521162 9353
rect 521106 9279 521162 9288
rect 521120 8265 521148 9279
rect 521106 8256 521162 8265
rect 521106 8191 521162 8200
rect 520370 7984 520426 7993
rect 520370 7919 520426 7928
rect 117320 7812 117372 7818
rect 117320 7754 117372 7760
rect 117228 7676 117280 7682
rect 116964 3369 116992 7670
rect 117228 7618 117280 7624
rect 117332 7562 117360 7754
rect 117240 7534 117360 7562
rect 117044 7472 117096 7478
rect 117044 7414 117096 7420
rect 117056 5681 117084 7414
rect 117134 6896 117190 6905
rect 117134 6831 117190 6840
rect 117042 5672 117098 5681
rect 117042 5607 117098 5616
rect 116950 3360 117006 3369
rect 116950 3295 117006 3304
rect 117148 1465 117176 6831
rect 117134 1456 117190 1465
rect 117134 1391 117190 1400
rect 117240 1154 117268 7534
rect 520384 6769 520412 7919
rect 520370 6760 520426 6769
rect 520370 6695 520426 6704
rect 521106 6624 521162 6633
rect 521106 6559 521162 6568
rect 521120 5273 521148 6559
rect 520922 5264 520978 5273
rect 520922 5199 520978 5208
rect 521106 5264 521162 5273
rect 521106 5199 521162 5208
rect 520936 3777 520964 5199
rect 521014 3904 521070 3913
rect 521014 3839 521070 3848
rect 520922 3768 520978 3777
rect 520922 3703 520978 3712
rect 193600 2514 193936 2530
rect 443656 2514 443992 2530
rect 170312 2508 170364 2514
rect 170312 2450 170364 2456
rect 193588 2508 193936 2514
rect 193640 2502 193936 2508
rect 294788 2508 294840 2514
rect 193588 2450 193640 2456
rect 294788 2450 294840 2456
rect 425796 2508 425848 2514
rect 425796 2450 425848 2456
rect 443644 2508 443992 2514
rect 443696 2502 443992 2508
rect 443644 2450 443696 2456
rect 170324 2378 170352 2450
rect 170312 2372 170364 2378
rect 170312 2314 170364 2320
rect 143644 2094 143980 2122
rect 243648 2094 243984 2122
rect 293604 2094 293940 2122
rect 143644 1494 143672 2094
rect 229282 1592 229338 1601
rect 229282 1527 229338 1536
rect 143632 1488 143684 1494
rect 143632 1430 143684 1436
rect 163778 1456 163834 1465
rect 163778 1391 163834 1400
rect 117228 1148 117280 1154
rect 117228 1090 117280 1096
rect 116860 1012 116912 1018
rect 116860 954 116912 960
rect 112536 944 112588 950
rect 112536 886 112588 892
rect 101864 808 101916 814
rect 96344 750 96396 756
rect 98274 -400 98330 800
rect 163792 800 163820 1391
rect 229296 800 229324 1527
rect 243648 1465 243676 2094
rect 293604 1601 293632 2094
rect 293590 1592 293646 1601
rect 293590 1527 293646 1536
rect 243634 1456 243690 1465
rect 294800 1426 294828 2450
rect 343652 2094 343988 2122
rect 393608 2094 393944 2122
rect 343652 1426 343680 2094
rect 393608 1465 393636 2094
rect 360290 1456 360346 1465
rect 243634 1391 243690 1400
rect 294788 1420 294840 1426
rect 294788 1362 294840 1368
rect 343640 1420 343692 1426
rect 360290 1391 360346 1400
rect 393594 1456 393650 1465
rect 393594 1391 393650 1400
rect 343640 1362 343692 1368
rect 294800 800 294828 1362
rect 360304 800 360332 1391
rect 425808 800 425836 2450
rect 521028 2281 521056 3839
rect 521106 2680 521162 2689
rect 521106 2615 521162 2624
rect 521014 2272 521070 2281
rect 521014 2207 521070 2216
rect 493612 2094 493948 2122
rect 493612 1426 493640 2094
rect 491300 1420 491352 1426
rect 491300 1362 491352 1368
rect 493600 1420 493652 1426
rect 493600 1362 493652 1368
rect 491312 800 491340 1362
rect 101864 750 101916 756
rect 163778 -400 163834 800
rect 229282 -400 229338 800
rect 294786 -400 294842 800
rect 360290 -400 360346 800
rect 425794 -400 425850 800
rect 491298 -400 491354 800
rect 521120 785 521148 2615
rect 521106 776 521162 785
rect 521106 711 521162 720
<< via2 >>
rect 2962 153720 3018 153776
rect 16302 159296 16358 159352
rect 16578 153856 16634 153912
rect 19890 153992 19946 154048
rect 23018 159432 23074 159488
rect 12438 152496 12494 152552
rect 8850 152360 8906 152416
rect 6090 150592 6146 150648
rect 2686 150456 2742 150512
rect 28078 156576 28134 156632
rect 29826 159568 29882 159624
rect 31482 156712 31538 156768
rect 30378 154128 30434 154184
rect 33966 157936 34022 157992
rect 40682 158208 40738 158264
rect 44086 158072 44142 158128
rect 57518 158344 57574 158400
rect 55862 156848 55918 156904
rect 54298 154264 54354 154320
rect 65982 155488 66038 155544
rect 62578 155352 62634 155408
rect 72698 156984 72754 157040
rect 68466 155216 68522 155272
rect 76010 155760 76066 155816
rect 78586 155624 78642 155680
rect 85302 155896 85358 155952
rect 85578 154400 85634 154456
rect 104622 158480 104678 158536
rect 82818 149640 82874 149696
rect 109590 148008 109646 148064
rect 115570 157120 115626 157176
rect 111062 150456 111118 150512
rect 110970 147872 111026 147928
rect 110326 146376 110382 146432
rect 110326 106256 110382 106312
rect 111338 150592 111394 150648
rect 111338 147872 111394 147928
rect 113822 144200 113878 144256
rect 116122 145152 116178 145208
rect 116030 143248 116086 143304
rect 115294 141344 115350 141400
rect 116122 139440 116178 139496
rect 116122 137536 116178 137592
rect 115202 135496 115258 135552
rect 116030 133592 116086 133648
rect 114190 132776 114246 132832
rect 113914 121352 113970 121408
rect 114006 110064 114062 110120
rect 114098 98640 114154 98696
rect 114190 87216 114246 87272
rect 116122 131688 116178 131744
rect 116582 149640 116638 149696
rect 116490 129784 116546 129840
rect 116122 125976 116178 126032
rect 116122 124108 116124 124128
rect 116124 124108 116176 124128
rect 116176 124108 116178 124128
rect 116122 124072 116178 124108
rect 115938 122168 115994 122224
rect 116122 120128 116178 120184
rect 116122 118224 116178 118280
rect 116122 116320 116178 116376
rect 116122 114452 116124 114472
rect 116124 114452 116176 114472
rect 116176 114452 116178 114472
rect 116122 114416 116178 114452
rect 115938 112512 115994 112568
rect 116122 110608 116178 110664
rect 116122 108704 116178 108760
rect 116950 102856 117006 102912
rect 121734 153720 121790 153776
rect 121918 153720 121974 153776
rect 126242 152360 126298 152416
rect 126794 152360 126850 152416
rect 128818 152496 128874 152552
rect 131026 159296 131082 159352
rect 133602 159432 133658 159488
rect 132038 153856 132094 153912
rect 133602 153040 133658 153096
rect 134614 153992 134670 154048
rect 136546 153040 136602 153096
rect 138018 159568 138074 159624
rect 140410 156576 140466 156632
rect 143078 156712 143134 156768
rect 142342 154128 142398 154184
rect 142618 154128 142674 154184
rect 142434 153892 142436 153912
rect 142436 153892 142488 153912
rect 142488 153892 142490 153912
rect 142434 153856 142490 153892
rect 142986 153892 142988 153912
rect 142988 153892 143040 153912
rect 143040 153892 143042 153912
rect 142986 153856 143042 153892
rect 142710 153332 142766 153368
rect 142710 153312 142712 153332
rect 142712 153312 142764 153332
rect 142764 153312 142766 153332
rect 143446 154148 143502 154184
rect 143446 154128 143448 154148
rect 143448 154128 143500 154148
rect 143500 154128 143502 154148
rect 143354 153312 143410 153368
rect 144918 157936 144974 157992
rect 143630 152360 143686 152416
rect 147586 154164 147588 154184
rect 147588 154164 147640 154184
rect 147640 154164 147642 154184
rect 147586 154128 147642 154164
rect 148138 154128 148194 154184
rect 149610 158208 149666 158264
rect 152554 158072 152610 158128
rect 161570 156848 161626 156904
rect 160926 154264 160982 154320
rect 162858 158344 162914 158400
rect 166722 155352 166778 155408
rect 168470 155488 168526 155544
rect 169666 158380 169668 158400
rect 169668 158380 169720 158400
rect 169720 158380 169722 158400
rect 169666 158344 169722 158380
rect 171230 155216 171286 155272
rect 173162 158380 173164 158400
rect 173164 158380 173216 158400
rect 173216 158380 173218 158400
rect 173162 158344 173218 158380
rect 174450 156984 174506 157040
rect 177026 155760 177082 155816
rect 178958 155624 179014 155680
rect 184018 155896 184074 155952
rect 184662 154400 184718 154456
rect 186318 155080 186374 155136
rect 187238 155080 187294 155136
rect 186870 154128 186926 154184
rect 189814 154128 189870 154184
rect 192390 153720 192446 153776
rect 195886 153584 195942 153640
rect 196070 153620 196072 153640
rect 196072 153620 196124 153640
rect 196124 153620 196126 153640
rect 196070 153584 196126 153620
rect 198738 158480 198794 158536
rect 204718 159296 204774 159352
rect 207202 157120 207258 157176
rect 209778 156712 209834 156768
rect 210606 156712 210662 156768
rect 211526 153720 211582 153776
rect 227442 152360 227498 152416
rect 274546 159432 274602 159488
rect 275190 159296 275246 159352
rect 280986 153720 281042 153776
rect 292578 152360 292634 152416
rect 313370 152360 313426 152416
rect 328550 159432 328606 159488
rect 357438 152360 357494 152416
rect 407670 152360 407726 152416
rect 430578 152360 430634 152416
rect 431866 152496 431922 152552
rect 448610 152496 448666 152552
rect 519358 154128 519414 154184
rect 519726 163104 519782 163160
rect 519542 161608 519598 161664
rect 519634 160112 519690 160168
rect 519542 147872 519598 147928
rect 520186 158616 520242 158672
rect 520002 157120 520058 157176
rect 519818 151136 519874 151192
rect 519726 149232 519782 149288
rect 519726 148144 519782 148200
rect 519634 146512 519690 146568
rect 519634 145152 519690 145208
rect 519542 142160 519598 142216
rect 519450 141072 519506 141128
rect 519266 140528 519322 140584
rect 519358 139032 519414 139088
rect 519266 128832 519322 128888
rect 117226 127880 117282 127936
rect 519450 133048 519506 133104
rect 519358 127472 519414 127528
rect 519358 124072 519414 124128
rect 519266 122576 519322 122632
rect 519910 149640 519966 149696
rect 519818 138352 519874 138408
rect 520094 155624 520150 155680
rect 520002 143792 520058 143848
rect 521014 152632 521070 152688
rect 520186 145288 520242 145344
rect 520922 143656 520978 143712
rect 520094 142432 520150 142488
rect 520094 137536 520150 137592
rect 519910 136992 519966 137048
rect 519910 136040 519966 136096
rect 519726 135632 519782 135688
rect 519634 132912 519690 132968
rect 519634 131416 519690 131472
rect 519542 130192 519598 130248
rect 519542 125568 519598 125624
rect 519450 122032 519506 122088
rect 519726 130056 519782 130112
rect 519634 120672 519690 120728
rect 519818 127064 519874 127120
rect 519726 119312 519782 119368
rect 520002 128560 520058 128616
rect 519910 124752 519966 124808
rect 519910 121080 519966 121136
rect 519818 116592 519874 116648
rect 519542 115232 519598 115288
rect 519818 114960 519874 115016
rect 519358 113872 519414 113928
rect 519726 113464 519782 113520
rect 519266 112512 519322 112568
rect 519542 111968 519598 112024
rect 117134 104760 117190 104816
rect 519634 110472 519690 110528
rect 519542 102992 519598 103048
rect 520186 134544 520242 134600
rect 520094 126112 520150 126168
rect 521106 146648 521162 146704
rect 521014 139712 521070 139768
rect 521106 134272 521162 134328
rect 520922 131552 520978 131608
rect 520186 123392 520242 123448
rect 520094 119584 520150 119640
rect 520002 117952 520058 118008
rect 520002 116456 520058 116512
rect 519910 111152 519966 111208
rect 520186 118088 520242 118144
rect 520094 109792 520150 109848
rect 520922 108976 520978 109032
rect 520186 108432 520242 108488
rect 520002 107072 520058 107128
rect 520278 105984 520334 106040
rect 519818 105712 519874 105768
rect 519726 104352 519782 104408
rect 519634 101632 519690 101688
rect 117042 100952 117098 101008
rect 116858 99048 116914 99104
rect 520830 104488 520886 104544
rect 520738 102992 520794 103048
rect 520278 97552 520334 97608
rect 116766 97144 116822 97200
rect 520278 95512 520334 95568
rect 116674 95240 116730 95296
rect 116582 93336 116638 93392
rect 520186 92384 520242 92440
rect 116122 91296 116178 91352
rect 520002 90888 520058 90944
rect 116122 89392 116178 89448
rect 519634 89392 519690 89448
rect 116030 87488 116086 87544
rect 519082 86400 519138 86456
rect 115202 85584 115258 85640
rect 116582 83680 116638 83736
rect 116214 81776 116270 81832
rect 519910 87896 519966 87952
rect 519818 84904 519874 84960
rect 519634 82592 519690 82648
rect 519726 81912 519782 81968
rect 115938 79872 115994 79928
rect 519082 79872 519138 79928
rect 519634 78920 519690 78976
rect 116122 77968 116178 78024
rect 116674 74024 116730 74080
rect 116582 72120 116638 72176
rect 113362 64504 113418 64560
rect 110326 53896 110382 53952
rect 110326 52536 110382 52592
rect 110326 51040 110382 51096
rect 109498 3848 109554 3904
rect 109498 3440 109554 3496
rect 32402 2624 32458 2680
rect 36358 2624 36414 2680
rect 62394 2624 62450 2680
rect 64142 2624 64198 2680
rect 65338 2624 65394 2680
rect 68006 2624 68062 2680
rect 68466 2624 68522 2680
rect 68834 2624 68890 2680
rect 69386 2624 69442 2680
rect 77022 2624 77078 2680
rect 29550 2352 29606 2408
rect 26054 2216 26110 2272
rect 5998 1672 6054 1728
rect 22926 2080 22982 2136
rect 19614 1944 19670 2000
rect 15934 1808 15990 1864
rect 12622 1536 12678 1592
rect 9310 1400 9366 1456
rect 33046 2488 33102 2544
rect 77252 2624 77308 2680
rect 77758 2624 77814 2680
rect 79966 2624 80022 2680
rect 80242 2624 80298 2680
rect 80426 2624 80482 2680
rect 80610 2624 80666 2680
rect 80794 2624 80850 2680
rect 93030 2624 93086 2680
rect 94686 2624 94742 2680
rect 96342 2624 96398 2680
rect 100114 2624 100170 2680
rect 101862 2624 101918 2680
rect 94318 2488 94374 2544
rect 94134 2080 94190 2136
rect 94318 2080 94374 2136
rect 85946 1264 86002 1320
rect 89258 856 89314 912
rect 95974 992 96030 1048
rect 96434 2488 96490 2544
rect 99838 2488 99894 2544
rect 96434 2080 96490 2136
rect 96618 2080 96674 2136
rect 99654 2080 99710 2136
rect 99838 2080 99894 2136
rect 98274 1264 98330 1320
rect 101494 2488 101550 2544
rect 100850 2352 100906 2408
rect 101402 2352 101458 2408
rect 100758 1944 100814 2000
rect 101218 1944 101274 2000
rect 101494 856 101550 912
rect 103426 2624 103482 2680
rect 103610 2624 103666 2680
rect 104162 2488 104218 2544
rect 104162 2080 104218 2136
rect 104346 2080 104402 2136
rect 103334 1264 103390 1320
rect 108210 1264 108266 1320
rect 103426 1128 103482 1184
rect 103886 1128 103942 1184
rect 108302 1128 108358 1184
rect 109682 3576 109738 3632
rect 109866 2760 109922 2816
rect 109498 1672 109554 1728
rect 110326 48320 110382 48376
rect 110326 47096 110382 47152
rect 110326 44240 110382 44296
rect 110326 41384 110382 41440
rect 110326 34584 110382 34640
rect 110326 8336 110382 8392
rect 110510 8336 110566 8392
rect 110050 3848 110106 3904
rect 110234 3848 110290 3904
rect 110234 3440 110290 3496
rect 110602 5616 110658 5672
rect 111062 7928 111118 7984
rect 110694 3168 110750 3224
rect 110602 2760 110658 2816
rect 111706 2916 111762 2952
rect 111706 2896 111708 2916
rect 111708 2896 111760 2916
rect 111760 2896 111762 2916
rect 110418 1264 110474 1320
rect 110050 992 110106 1048
rect 116306 70216 116362 70272
rect 116122 68312 116178 68368
rect 116582 66408 116638 66464
rect 521106 107480 521162 107536
rect 521014 101496 521070 101552
rect 520922 100272 520978 100328
rect 520922 98504 520978 98560
rect 520830 96192 520886 96248
rect 520738 94832 520794 94888
rect 521198 100000 521254 100056
rect 521106 98912 521162 98968
rect 521106 93880 521162 93936
rect 521014 93472 521070 93528
rect 520922 90752 520978 90808
rect 520278 88032 520334 88088
rect 521382 97008 521438 97064
rect 521198 92112 521254 92168
rect 521382 89528 521438 89584
rect 521106 86672 521162 86728
rect 520186 85312 520242 85368
rect 520002 83952 520058 84008
rect 520186 83408 520242 83464
rect 519910 81232 519966 81288
rect 520002 80416 520058 80472
rect 519818 78512 519874 78568
rect 519910 77424 519966 77480
rect 519726 75928 519782 75984
rect 519634 73208 519690 73264
rect 520186 77152 520242 77208
rect 520186 75928 520242 75984
rect 520002 74568 520058 74624
rect 519910 71848 519966 71904
rect 521014 74432 521070 74488
rect 520922 72936 520978 72992
rect 520186 70488 520242 70544
rect 521198 71440 521254 71496
rect 521106 69808 521162 69864
rect 521014 69128 521070 69184
rect 521014 68312 521070 68368
rect 520922 67768 520978 67824
rect 520462 66816 520518 66872
rect 520370 65320 520426 65376
rect 116214 64504 116270 64560
rect 116122 62600 116178 62656
rect 521198 66408 521254 66464
rect 521106 65048 521162 65104
rect 521106 63824 521162 63880
rect 521014 63688 521070 63744
rect 520462 62328 520518 62384
rect 521014 62328 521070 62384
rect 520370 60968 520426 61024
rect 520738 60832 520794 60888
rect 116582 60560 116638 60616
rect 114190 53080 114246 53136
rect 116122 43288 116178 43344
rect 114098 41792 114154 41848
rect 114006 30368 114062 30424
rect 116490 27920 116546 27976
rect 116306 26016 116362 26072
rect 116214 22208 116270 22264
rect 116030 20304 116086 20360
rect 113914 18944 113970 19000
rect 115938 16360 115994 16416
rect 113822 7656 113878 7712
rect 116122 18400 116178 18456
rect 116030 2488 116086 2544
rect 116398 24112 116454 24168
rect 116306 3576 116362 3632
rect 116306 3032 116362 3088
rect 116214 2624 116270 2680
rect 116122 2352 116178 2408
rect 115938 2216 115994 2272
rect 116766 58656 116822 58712
rect 116674 56752 116730 56808
rect 519910 57840 519966 57896
rect 519818 56344 519874 56400
rect 519082 53352 519138 53408
rect 521106 59608 521162 59664
rect 521106 59336 521162 59392
rect 521014 58248 521070 58304
rect 520738 56888 520794 56944
rect 521106 55528 521162 55584
rect 520186 54848 520242 54904
rect 519910 54168 519966 54224
rect 519818 52808 519874 52864
rect 520094 51856 520150 51912
rect 519082 50088 519138 50144
rect 519082 48864 519138 48920
rect 520186 51448 520242 51504
rect 520186 50360 520242 50416
rect 520094 48728 520150 48784
rect 520186 47368 520242 47424
rect 519910 47232 519966 47288
rect 519082 46008 519138 46064
rect 519726 45736 519782 45792
rect 519910 44648 519966 44704
rect 520186 44240 520242 44296
rect 519726 43288 519782 43344
rect 520738 42744 520794 42800
rect 520186 41928 520242 41984
rect 520738 41248 520794 41304
rect 520922 41248 520978 41304
rect 520922 39888 520978 39944
rect 520922 39752 520978 39808
rect 116950 39480 117006 39536
rect 116858 37576 116914 37632
rect 116766 7928 116822 7984
rect 521106 38256 521162 38312
rect 520922 37848 520978 37904
rect 521106 37168 521162 37224
rect 521566 36760 521622 36816
rect 521566 35944 521622 36000
rect 520922 35264 520978 35320
rect 520922 34448 520978 34504
rect 117134 33768 117190 33824
rect 521106 33768 521162 33824
rect 117042 31728 117098 31784
rect 521106 33088 521162 33144
rect 521106 32272 521162 32328
rect 521106 31592 521162 31648
rect 117226 29824 117282 29880
rect 116674 3168 116730 3224
rect 520922 29280 520978 29336
rect 520922 28328 520978 28384
rect 521106 24792 521162 24848
rect 521106 23568 521162 23624
rect 520370 23160 520426 23216
rect 520370 22208 520426 22264
rect 520922 21664 520978 21720
rect 520922 20848 520978 20904
rect 521106 20168 521162 20224
rect 521106 19488 521162 19544
rect 521106 9288 521162 9344
rect 521106 8200 521162 8256
rect 520370 7928 520426 7984
rect 117134 6840 117190 6896
rect 117042 5616 117098 5672
rect 116950 3304 117006 3360
rect 117134 1400 117190 1456
rect 520370 6704 520426 6760
rect 521106 6568 521162 6624
rect 520922 5208 520978 5264
rect 521106 5208 521162 5264
rect 521014 3848 521070 3904
rect 520922 3712 520978 3768
rect 229282 1536 229338 1592
rect 163778 1400 163834 1456
rect 293590 1536 293646 1592
rect 243634 1400 243690 1456
rect 360290 1400 360346 1456
rect 393594 1400 393650 1456
rect 521106 2624 521162 2680
rect 521014 2216 521070 2272
rect 521106 720 521162 776
<< metal3 >>
rect 519721 163162 519787 163165
rect 523200 163162 524400 163192
rect 519721 163160 524400 163162
rect 519721 163104 519726 163160
rect 519782 163104 524400 163160
rect 519721 163102 524400 163104
rect 519721 163099 519787 163102
rect 523200 163072 524400 163102
rect 519537 161666 519603 161669
rect 523200 161666 524400 161696
rect 519537 161664 524400 161666
rect 519537 161608 519542 161664
rect 519598 161608 524400 161664
rect 519537 161606 524400 161608
rect 519537 161603 519603 161606
rect 523200 161576 524400 161606
rect 519629 160170 519695 160173
rect 523200 160170 524400 160200
rect 519629 160168 524400 160170
rect 519629 160112 519634 160168
rect 519690 160112 524400 160168
rect 519629 160110 524400 160112
rect 519629 160107 519695 160110
rect 523200 160080 524400 160110
rect 29821 159626 29887 159629
rect 138013 159626 138079 159629
rect 29821 159624 138079 159626
rect 29821 159568 29826 159624
rect 29882 159568 138018 159624
rect 138074 159568 138079 159624
rect 29821 159566 138079 159568
rect 29821 159563 29887 159566
rect 138013 159563 138079 159566
rect 23013 159490 23079 159493
rect 133597 159490 133663 159493
rect 23013 159488 133663 159490
rect 23013 159432 23018 159488
rect 23074 159432 133602 159488
rect 133658 159432 133663 159488
rect 23013 159430 133663 159432
rect 23013 159427 23079 159430
rect 133597 159427 133663 159430
rect 274541 159490 274607 159493
rect 328545 159490 328611 159493
rect 274541 159488 328611 159490
rect 274541 159432 274546 159488
rect 274602 159432 328550 159488
rect 328606 159432 328611 159488
rect 274541 159430 328611 159432
rect 274541 159427 274607 159430
rect 328545 159427 328611 159430
rect 16297 159354 16363 159357
rect 131021 159354 131087 159357
rect 16297 159352 131087 159354
rect 16297 159296 16302 159352
rect 16358 159296 131026 159352
rect 131082 159296 131087 159352
rect 16297 159294 131087 159296
rect 16297 159291 16363 159294
rect 131021 159291 131087 159294
rect 204713 159354 204779 159357
rect 275185 159354 275251 159357
rect 204713 159352 275251 159354
rect 204713 159296 204718 159352
rect 204774 159296 275190 159352
rect 275246 159296 275251 159352
rect 204713 159294 275251 159296
rect 204713 159291 204779 159294
rect 275185 159291 275251 159294
rect 520181 158674 520247 158677
rect 523200 158674 524400 158704
rect 520181 158672 524400 158674
rect 520181 158616 520186 158672
rect 520242 158616 524400 158672
rect 520181 158614 524400 158616
rect 520181 158611 520247 158614
rect 523200 158584 524400 158614
rect 104617 158538 104683 158541
rect 198733 158538 198799 158541
rect 104617 158536 198799 158538
rect 104617 158480 104622 158536
rect 104678 158480 198738 158536
rect 198794 158480 198799 158536
rect 104617 158478 198799 158480
rect 104617 158475 104683 158478
rect 198733 158475 198799 158478
rect 57513 158402 57579 158405
rect 162853 158402 162919 158405
rect 57513 158400 162919 158402
rect 57513 158344 57518 158400
rect 57574 158344 162858 158400
rect 162914 158344 162919 158400
rect 57513 158342 162919 158344
rect 57513 158339 57579 158342
rect 162853 158339 162919 158342
rect 169661 158402 169727 158405
rect 173157 158402 173223 158405
rect 169661 158400 173223 158402
rect 169661 158344 169666 158400
rect 169722 158344 173162 158400
rect 173218 158344 173223 158400
rect 169661 158342 173223 158344
rect 169661 158339 169727 158342
rect 173157 158339 173223 158342
rect 40677 158266 40743 158269
rect 149605 158266 149671 158269
rect 40677 158264 149671 158266
rect 40677 158208 40682 158264
rect 40738 158208 149610 158264
rect 149666 158208 149671 158264
rect 40677 158206 149671 158208
rect 40677 158203 40743 158206
rect 149605 158203 149671 158206
rect 44081 158130 44147 158133
rect 152549 158130 152615 158133
rect 44081 158128 152615 158130
rect 44081 158072 44086 158128
rect 44142 158072 152554 158128
rect 152610 158072 152615 158128
rect 44081 158070 152615 158072
rect 44081 158067 44147 158070
rect 152549 158067 152615 158070
rect 33961 157994 34027 157997
rect 144913 157994 144979 157997
rect 33961 157992 144979 157994
rect 33961 157936 33966 157992
rect 34022 157936 144918 157992
rect 144974 157936 144979 157992
rect 33961 157934 144979 157936
rect 33961 157931 34027 157934
rect 144913 157931 144979 157934
rect 115565 157178 115631 157181
rect 207197 157178 207263 157181
rect 115565 157176 207263 157178
rect 115565 157120 115570 157176
rect 115626 157120 207202 157176
rect 207258 157120 207263 157176
rect 115565 157118 207263 157120
rect 115565 157115 115631 157118
rect 207197 157115 207263 157118
rect 519997 157178 520063 157181
rect 523200 157178 524400 157208
rect 519997 157176 524400 157178
rect 519997 157120 520002 157176
rect 520058 157120 524400 157176
rect 519997 157118 524400 157120
rect 519997 157115 520063 157118
rect 523200 157088 524400 157118
rect 72693 157042 72759 157045
rect 174445 157042 174511 157045
rect 72693 157040 174511 157042
rect 72693 156984 72698 157040
rect 72754 156984 174450 157040
rect 174506 156984 174511 157040
rect 72693 156982 174511 156984
rect 72693 156979 72759 156982
rect 174445 156979 174511 156982
rect 55857 156906 55923 156909
rect 161565 156906 161631 156909
rect 55857 156904 161631 156906
rect 55857 156848 55862 156904
rect 55918 156848 161570 156904
rect 161626 156848 161631 156904
rect 55857 156846 161631 156848
rect 55857 156843 55923 156846
rect 161565 156843 161631 156846
rect 31477 156770 31543 156773
rect 143073 156770 143139 156773
rect 31477 156768 143139 156770
rect 31477 156712 31482 156768
rect 31538 156712 143078 156768
rect 143134 156712 143139 156768
rect 31477 156710 143139 156712
rect 31477 156707 31543 156710
rect 143073 156707 143139 156710
rect 209773 156770 209839 156773
rect 210601 156770 210667 156773
rect 209773 156768 210667 156770
rect 209773 156712 209778 156768
rect 209834 156712 210606 156768
rect 210662 156712 210667 156768
rect 209773 156710 210667 156712
rect 209773 156707 209839 156710
rect 210601 156707 210667 156710
rect 28073 156634 28139 156637
rect 140405 156634 140471 156637
rect 28073 156632 140471 156634
rect 28073 156576 28078 156632
rect 28134 156576 140410 156632
rect 140466 156576 140471 156632
rect 28073 156574 140471 156576
rect 28073 156571 28139 156574
rect 140405 156571 140471 156574
rect 85297 155954 85363 155957
rect 184013 155954 184079 155957
rect 85297 155952 184079 155954
rect 85297 155896 85302 155952
rect 85358 155896 184018 155952
rect 184074 155896 184079 155952
rect 85297 155894 184079 155896
rect 85297 155891 85363 155894
rect 184013 155891 184079 155894
rect 76005 155818 76071 155821
rect 177021 155818 177087 155821
rect 76005 155816 177087 155818
rect 76005 155760 76010 155816
rect 76066 155760 177026 155816
rect 177082 155760 177087 155816
rect 76005 155758 177087 155760
rect 76005 155755 76071 155758
rect 177021 155755 177087 155758
rect 78581 155682 78647 155685
rect 178953 155682 179019 155685
rect 78581 155680 179019 155682
rect 78581 155624 78586 155680
rect 78642 155624 178958 155680
rect 179014 155624 179019 155680
rect 78581 155622 179019 155624
rect 78581 155619 78647 155622
rect 178953 155619 179019 155622
rect 520089 155682 520155 155685
rect 523200 155682 524400 155712
rect 520089 155680 524400 155682
rect 520089 155624 520094 155680
rect 520150 155624 524400 155680
rect 520089 155622 524400 155624
rect 520089 155619 520155 155622
rect 523200 155592 524400 155622
rect 65977 155546 66043 155549
rect 168465 155546 168531 155549
rect 65977 155544 168531 155546
rect 65977 155488 65982 155544
rect 66038 155488 168470 155544
rect 168526 155488 168531 155544
rect 65977 155486 168531 155488
rect 65977 155483 66043 155486
rect 168465 155483 168531 155486
rect 62573 155410 62639 155413
rect 166717 155410 166783 155413
rect 62573 155408 166783 155410
rect 62573 155352 62578 155408
rect 62634 155352 166722 155408
rect 166778 155352 166783 155408
rect 62573 155350 166783 155352
rect 62573 155347 62639 155350
rect 166717 155347 166783 155350
rect 68461 155274 68527 155277
rect 171225 155274 171291 155277
rect 68461 155272 171291 155274
rect 68461 155216 68466 155272
rect 68522 155216 171230 155272
rect 171286 155216 171291 155272
rect 68461 155214 171291 155216
rect 68461 155211 68527 155214
rect 171225 155211 171291 155214
rect 186313 155138 186379 155141
rect 187233 155138 187299 155141
rect 186313 155136 187299 155138
rect 186313 155080 186318 155136
rect 186374 155080 187238 155136
rect 187294 155080 187299 155136
rect 186313 155078 187299 155080
rect 186313 155075 186379 155078
rect 187233 155075 187299 155078
rect 85573 154458 85639 154461
rect 184657 154458 184723 154461
rect 85573 154456 184723 154458
rect 85573 154400 85578 154456
rect 85634 154400 184662 154456
rect 184718 154400 184723 154456
rect 85573 154398 184723 154400
rect 85573 154395 85639 154398
rect 184657 154395 184723 154398
rect 54293 154322 54359 154325
rect 160921 154322 160987 154325
rect 54293 154320 160987 154322
rect 54293 154264 54298 154320
rect 54354 154264 160926 154320
rect 160982 154264 160987 154320
rect 54293 154262 160987 154264
rect 54293 154259 54359 154262
rect 160921 154259 160987 154262
rect 30373 154186 30439 154189
rect 142337 154186 142403 154189
rect 30373 154184 142403 154186
rect 30373 154128 30378 154184
rect 30434 154128 142342 154184
rect 142398 154128 142403 154184
rect 30373 154126 142403 154128
rect 30373 154123 30439 154126
rect 142337 154123 142403 154126
rect 142613 154186 142679 154189
rect 143441 154186 143507 154189
rect 142613 154184 143507 154186
rect 142613 154128 142618 154184
rect 142674 154128 143446 154184
rect 143502 154128 143507 154184
rect 142613 154126 143507 154128
rect 142613 154123 142679 154126
rect 143441 154123 143507 154126
rect 147581 154186 147647 154189
rect 148133 154186 148199 154189
rect 147581 154184 148199 154186
rect 147581 154128 147586 154184
rect 147642 154128 148138 154184
rect 148194 154128 148199 154184
rect 147581 154126 148199 154128
rect 147581 154123 147647 154126
rect 148133 154123 148199 154126
rect 186865 154186 186931 154189
rect 189809 154186 189875 154189
rect 186865 154184 189875 154186
rect 186865 154128 186870 154184
rect 186926 154128 189814 154184
rect 189870 154128 189875 154184
rect 186865 154126 189875 154128
rect 186865 154123 186931 154126
rect 189809 154123 189875 154126
rect 519353 154186 519419 154189
rect 523200 154186 524400 154216
rect 519353 154184 524400 154186
rect 519353 154128 519358 154184
rect 519414 154128 524400 154184
rect 519353 154126 524400 154128
rect 519353 154123 519419 154126
rect 523200 154096 524400 154126
rect 19885 154050 19951 154053
rect 134609 154050 134675 154053
rect 19885 154048 134675 154050
rect 19885 153992 19890 154048
rect 19946 153992 134614 154048
rect 134670 153992 134675 154048
rect 19885 153990 134675 153992
rect 19885 153987 19951 153990
rect 134609 153987 134675 153990
rect 16573 153914 16639 153917
rect 132033 153914 132099 153917
rect 16573 153912 132099 153914
rect 16573 153856 16578 153912
rect 16634 153856 132038 153912
rect 132094 153856 132099 153912
rect 16573 153854 132099 153856
rect 16573 153851 16639 153854
rect 132033 153851 132099 153854
rect 142429 153914 142495 153917
rect 142981 153914 143047 153917
rect 142429 153912 143047 153914
rect 142429 153856 142434 153912
rect 142490 153856 142986 153912
rect 143042 153856 143047 153912
rect 142429 153854 143047 153856
rect 142429 153851 142495 153854
rect 142981 153851 143047 153854
rect 2957 153778 3023 153781
rect 121729 153778 121795 153781
rect 2957 153776 121795 153778
rect 2957 153720 2962 153776
rect 3018 153720 121734 153776
rect 121790 153720 121795 153776
rect 2957 153718 121795 153720
rect 2957 153715 3023 153718
rect 121729 153715 121795 153718
rect 121913 153778 121979 153781
rect 192385 153778 192451 153781
rect 121913 153776 192451 153778
rect 121913 153720 121918 153776
rect 121974 153720 192390 153776
rect 192446 153720 192451 153776
rect 121913 153718 192451 153720
rect 121913 153715 121979 153718
rect 192385 153715 192451 153718
rect 211521 153778 211587 153781
rect 280981 153778 281047 153781
rect 211521 153776 281047 153778
rect 211521 153720 211526 153776
rect 211582 153720 280986 153776
rect 281042 153720 281047 153776
rect 211521 153718 281047 153720
rect 211521 153715 211587 153718
rect 280981 153715 281047 153718
rect 195881 153642 195947 153645
rect 196065 153642 196131 153645
rect 195881 153640 196131 153642
rect 195881 153584 195886 153640
rect 195942 153584 196070 153640
rect 196126 153584 196131 153640
rect 195881 153582 196131 153584
rect 195881 153579 195947 153582
rect 196065 153579 196131 153582
rect 142705 153370 142771 153373
rect 143349 153370 143415 153373
rect 142705 153368 143415 153370
rect 142705 153312 142710 153368
rect 142766 153312 143354 153368
rect 143410 153312 143415 153368
rect 142705 153310 143415 153312
rect 142705 153307 142771 153310
rect 143349 153307 143415 153310
rect 133597 153098 133663 153101
rect 136541 153098 136607 153101
rect 133597 153096 136607 153098
rect 133597 153040 133602 153096
rect 133658 153040 136546 153096
rect 136602 153040 136607 153096
rect 133597 153038 136607 153040
rect 133597 153035 133663 153038
rect 136541 153035 136607 153038
rect 521009 152690 521075 152693
rect 523200 152690 524400 152720
rect 521009 152688 524400 152690
rect 521009 152632 521014 152688
rect 521070 152632 524400 152688
rect 521009 152630 524400 152632
rect 521009 152627 521075 152630
rect 523200 152600 524400 152630
rect 12433 152554 12499 152557
rect 128813 152554 128879 152557
rect 12433 152552 128879 152554
rect 12433 152496 12438 152552
rect 12494 152496 128818 152552
rect 128874 152496 128879 152552
rect 12433 152494 128879 152496
rect 12433 152491 12499 152494
rect 128813 152491 128879 152494
rect 431861 152554 431927 152557
rect 448605 152554 448671 152557
rect 431861 152552 448671 152554
rect 431861 152496 431866 152552
rect 431922 152496 448610 152552
rect 448666 152496 448671 152552
rect 431861 152494 448671 152496
rect 431861 152491 431927 152494
rect 448605 152491 448671 152494
rect 8845 152418 8911 152421
rect 126237 152418 126303 152421
rect 8845 152416 126303 152418
rect 8845 152360 8850 152416
rect 8906 152360 126242 152416
rect 126298 152360 126303 152416
rect 8845 152358 126303 152360
rect 8845 152355 8911 152358
rect 126237 152355 126303 152358
rect 126789 152418 126855 152421
rect 143625 152418 143691 152421
rect 126789 152416 143691 152418
rect 126789 152360 126794 152416
rect 126850 152360 143630 152416
rect 143686 152360 143691 152416
rect 126789 152358 143691 152360
rect 126789 152355 126855 152358
rect 143625 152355 143691 152358
rect 227437 152418 227503 152421
rect 292573 152418 292639 152421
rect 227437 152416 292639 152418
rect 227437 152360 227442 152416
rect 227498 152360 292578 152416
rect 292634 152360 292639 152416
rect 227437 152358 292639 152360
rect 227437 152355 227503 152358
rect 292573 152355 292639 152358
rect 313365 152418 313431 152421
rect 357433 152418 357499 152421
rect 313365 152416 357499 152418
rect 313365 152360 313370 152416
rect 313426 152360 357438 152416
rect 357494 152360 357499 152416
rect 313365 152358 357499 152360
rect 313365 152355 313431 152358
rect 357433 152355 357499 152358
rect 407665 152418 407731 152421
rect 430573 152418 430639 152421
rect 407665 152416 430639 152418
rect 407665 152360 407670 152416
rect 407726 152360 430578 152416
rect 430634 152360 430639 152416
rect 407665 152358 430639 152360
rect 407665 152355 407731 152358
rect 430573 152355 430639 152358
rect 519813 151194 519879 151197
rect 523200 151194 524400 151224
rect 519813 151192 524400 151194
rect 519813 151136 519818 151192
rect 519874 151136 524400 151192
rect 519813 151134 524400 151136
rect 519813 151131 519879 151134
rect 523200 151104 524400 151134
rect 6085 150650 6151 150653
rect 111333 150650 111399 150653
rect 6085 150648 111399 150650
rect 6085 150592 6090 150648
rect 6146 150592 111338 150648
rect 111394 150592 111399 150648
rect 6085 150590 111399 150592
rect 6085 150587 6151 150590
rect 111333 150587 111399 150590
rect 2681 150514 2747 150517
rect 111057 150514 111123 150517
rect 2681 150512 111123 150514
rect 2681 150456 2686 150512
rect 2742 150456 111062 150512
rect 111118 150456 111123 150512
rect 2681 150454 111123 150456
rect 2681 150451 2747 150454
rect 111057 150451 111123 150454
rect 82813 149698 82879 149701
rect 116577 149698 116643 149701
rect 82813 149696 116643 149698
rect 82813 149640 82818 149696
rect 82874 149640 116582 149696
rect 116638 149640 116643 149696
rect 82813 149638 116643 149640
rect 82813 149635 82879 149638
rect 116577 149635 116643 149638
rect 519905 149698 519971 149701
rect 523200 149698 524400 149728
rect 519905 149696 524400 149698
rect 519905 149640 519910 149696
rect 519966 149640 524400 149696
rect 519905 149638 524400 149640
rect 519905 149635 519971 149638
rect 523200 149608 524400 149638
rect 519721 149290 519787 149293
rect 518788 149288 519787 149290
rect 518788 149232 519726 149288
rect 519782 149232 519787 149288
rect 518788 149230 519787 149232
rect 519721 149227 519787 149230
rect 109585 148066 109651 148069
rect 119110 148066 119170 148988
rect 519721 148202 519787 148205
rect 523200 148202 524400 148232
rect 519721 148200 524400 148202
rect 519721 148144 519726 148200
rect 519782 148144 524400 148200
rect 519721 148142 524400 148144
rect 519721 148139 519787 148142
rect 523200 148112 524400 148142
rect 109585 148064 119170 148066
rect 109585 148008 109590 148064
rect 109646 148008 119170 148064
rect 109585 148006 119170 148008
rect 109585 148003 109651 148006
rect 110965 147930 111031 147933
rect 111333 147930 111399 147933
rect 519537 147930 519603 147933
rect 110965 147928 111399 147930
rect 110965 147872 110970 147928
rect 111026 147872 111338 147928
rect 111394 147872 111399 147928
rect 110965 147870 111399 147872
rect 518788 147928 519603 147930
rect 518788 147872 519542 147928
rect 519598 147872 519603 147928
rect 518788 147870 519603 147872
rect 110965 147867 111031 147870
rect 111333 147867 111399 147870
rect 519537 147867 519603 147870
rect 110321 146434 110387 146437
rect 119110 146434 119170 147084
rect 521101 146706 521167 146709
rect 523200 146706 524400 146736
rect 521101 146704 524400 146706
rect 521101 146648 521106 146704
rect 521162 146648 524400 146704
rect 521101 146646 524400 146648
rect 521101 146643 521167 146646
rect 523200 146616 524400 146646
rect 519629 146570 519695 146573
rect 518788 146568 519695 146570
rect 518788 146512 519634 146568
rect 519690 146512 519695 146568
rect 518788 146510 519695 146512
rect 519629 146507 519695 146510
rect 110321 146432 119170 146434
rect 110321 146376 110326 146432
rect 110382 146376 119170 146432
rect 110321 146374 119170 146376
rect 110321 146371 110387 146374
rect 520181 145346 520247 145349
rect 518758 145344 520247 145346
rect 518758 145288 520186 145344
rect 520242 145288 520247 145344
rect 518758 145286 520247 145288
rect 116117 145210 116183 145213
rect 116117 145208 119140 145210
rect 116117 145152 116122 145208
rect 116178 145152 119140 145208
rect 518758 145180 518818 145286
rect 520181 145283 520247 145286
rect 519629 145210 519695 145213
rect 523200 145210 524400 145240
rect 519629 145208 524400 145210
rect 116117 145150 119140 145152
rect 519629 145152 519634 145208
rect 519690 145152 524400 145208
rect 519629 145150 524400 145152
rect 116117 145147 116183 145150
rect 519629 145147 519695 145150
rect 523200 145120 524400 145150
rect 113817 144258 113883 144261
rect 110860 144256 113883 144258
rect 110860 144200 113822 144256
rect 113878 144200 113883 144256
rect 110860 144198 113883 144200
rect 113817 144195 113883 144198
rect 519997 143850 520063 143853
rect 518788 143848 520063 143850
rect 518788 143792 520002 143848
rect 520058 143792 520063 143848
rect 518788 143790 520063 143792
rect 519997 143787 520063 143790
rect 520917 143714 520983 143717
rect 523200 143714 524400 143744
rect 520917 143712 524400 143714
rect 520917 143656 520922 143712
rect 520978 143656 524400 143712
rect 520917 143654 524400 143656
rect 520917 143651 520983 143654
rect 523200 143624 524400 143654
rect 116025 143306 116091 143309
rect 116025 143304 119140 143306
rect 116025 143248 116030 143304
rect 116086 143248 119140 143304
rect 116025 143246 119140 143248
rect 116025 143243 116091 143246
rect 520089 142490 520155 142493
rect 518788 142488 520155 142490
rect 518788 142432 520094 142488
rect 520150 142432 520155 142488
rect 518788 142430 520155 142432
rect 520089 142427 520155 142430
rect 519537 142218 519603 142221
rect 523200 142218 524400 142248
rect 519537 142216 524400 142218
rect 519537 142160 519542 142216
rect 519598 142160 524400 142216
rect 519537 142158 524400 142160
rect 519537 142155 519603 142158
rect 523200 142128 524400 142158
rect 115289 141402 115355 141405
rect 115289 141400 119140 141402
rect 115289 141344 115294 141400
rect 115350 141344 119140 141400
rect 115289 141342 119140 141344
rect 115289 141339 115355 141342
rect 519445 141130 519511 141133
rect 518788 141128 519511 141130
rect 518788 141072 519450 141128
rect 519506 141072 519511 141128
rect 518788 141070 519511 141072
rect 519445 141067 519511 141070
rect 519261 140586 519327 140589
rect 523200 140586 524400 140616
rect 519261 140584 524400 140586
rect 519261 140528 519266 140584
rect 519322 140528 524400 140584
rect 519261 140526 524400 140528
rect 519261 140523 519327 140526
rect 523200 140496 524400 140526
rect 521009 139770 521075 139773
rect 518788 139768 521075 139770
rect 518788 139712 521014 139768
rect 521070 139712 521075 139768
rect 518788 139710 521075 139712
rect 521009 139707 521075 139710
rect 116117 139498 116183 139501
rect 116117 139496 119140 139498
rect 116117 139440 116122 139496
rect 116178 139440 119140 139496
rect 116117 139438 119140 139440
rect 116117 139435 116183 139438
rect 519353 139090 519419 139093
rect 523200 139090 524400 139120
rect 519353 139088 524400 139090
rect 519353 139032 519358 139088
rect 519414 139032 524400 139088
rect 519353 139030 524400 139032
rect 519353 139027 519419 139030
rect 523200 139000 524400 139030
rect 519813 138410 519879 138413
rect 518788 138408 519879 138410
rect 518788 138352 519818 138408
rect 519874 138352 519879 138408
rect 518788 138350 519879 138352
rect 519813 138347 519879 138350
rect 116117 137594 116183 137597
rect 520089 137594 520155 137597
rect 523200 137594 524400 137624
rect 116117 137592 119140 137594
rect 116117 137536 116122 137592
rect 116178 137536 119140 137592
rect 116117 137534 119140 137536
rect 520089 137592 524400 137594
rect 520089 137536 520094 137592
rect 520150 137536 524400 137592
rect 520089 137534 524400 137536
rect 116117 137531 116183 137534
rect 520089 137531 520155 137534
rect 523200 137504 524400 137534
rect 519905 137050 519971 137053
rect 518788 137048 519971 137050
rect 518788 136992 519910 137048
rect 519966 136992 519971 137048
rect 518788 136990 519971 136992
rect 519905 136987 519971 136990
rect 519905 136098 519971 136101
rect 523200 136098 524400 136128
rect 519905 136096 524400 136098
rect 519905 136040 519910 136096
rect 519966 136040 524400 136096
rect 519905 136038 524400 136040
rect 519905 136035 519971 136038
rect 523200 136008 524400 136038
rect 519721 135690 519787 135693
rect 518788 135688 519787 135690
rect 518788 135632 519726 135688
rect 519782 135632 519787 135688
rect 518788 135630 519787 135632
rect 519721 135627 519787 135630
rect 115197 135554 115263 135557
rect 115197 135552 119140 135554
rect 115197 135496 115202 135552
rect 115258 135496 119140 135552
rect 115197 135494 119140 135496
rect 115197 135491 115263 135494
rect 520181 134602 520247 134605
rect 523200 134602 524400 134632
rect 520181 134600 524400 134602
rect 520181 134544 520186 134600
rect 520242 134544 524400 134600
rect 520181 134542 524400 134544
rect 520181 134539 520247 134542
rect 523200 134512 524400 134542
rect 521101 134330 521167 134333
rect 518788 134328 521167 134330
rect 518788 134272 521106 134328
rect 521162 134272 521167 134328
rect 518788 134270 521167 134272
rect 521101 134267 521167 134270
rect 116025 133650 116091 133653
rect 116025 133648 119140 133650
rect 116025 133592 116030 133648
rect 116086 133592 119140 133648
rect 116025 133590 119140 133592
rect 116025 133587 116091 133590
rect 519445 133106 519511 133109
rect 523200 133106 524400 133136
rect 519445 133104 524400 133106
rect 519445 133048 519450 133104
rect 519506 133048 524400 133104
rect 519445 133046 524400 133048
rect 519445 133043 519511 133046
rect 523200 133016 524400 133046
rect 519629 132970 519695 132973
rect 518788 132968 519695 132970
rect 518788 132912 519634 132968
rect 519690 132912 519695 132968
rect 518788 132910 519695 132912
rect 519629 132907 519695 132910
rect 114185 132834 114251 132837
rect 110860 132832 114251 132834
rect 110860 132776 114190 132832
rect 114246 132776 114251 132832
rect 110860 132774 114251 132776
rect 114185 132771 114251 132774
rect 116117 131746 116183 131749
rect 116117 131744 119140 131746
rect 116117 131688 116122 131744
rect 116178 131688 119140 131744
rect 116117 131686 119140 131688
rect 116117 131683 116183 131686
rect 520917 131610 520983 131613
rect 523200 131610 524400 131640
rect 518788 131608 520983 131610
rect 518788 131552 520922 131608
rect 520978 131552 520983 131608
rect 518788 131550 520983 131552
rect 520917 131547 520983 131550
rect 521518 131550 524400 131610
rect 519629 131474 519695 131477
rect 521518 131474 521578 131550
rect 523200 131520 524400 131550
rect 519629 131472 521578 131474
rect 519629 131416 519634 131472
rect 519690 131416 521578 131472
rect 519629 131414 521578 131416
rect 519629 131411 519695 131414
rect 519537 130250 519603 130253
rect 518788 130248 519603 130250
rect 518788 130192 519542 130248
rect 519598 130192 519603 130248
rect 518788 130190 519603 130192
rect 519537 130187 519603 130190
rect 519721 130114 519787 130117
rect 523200 130114 524400 130144
rect 519721 130112 524400 130114
rect 519721 130056 519726 130112
rect 519782 130056 524400 130112
rect 519721 130054 524400 130056
rect 519721 130051 519787 130054
rect 523200 130024 524400 130054
rect 116485 129842 116551 129845
rect 116485 129840 119140 129842
rect 116485 129784 116490 129840
rect 116546 129784 119140 129840
rect 116485 129782 119140 129784
rect 116485 129779 116551 129782
rect 519261 128890 519327 128893
rect 518788 128888 519327 128890
rect 518788 128832 519266 128888
rect 519322 128832 519327 128888
rect 518788 128830 519327 128832
rect 519261 128827 519327 128830
rect 519997 128618 520063 128621
rect 523200 128618 524400 128648
rect 519997 128616 524400 128618
rect 519997 128560 520002 128616
rect 520058 128560 524400 128616
rect 519997 128558 524400 128560
rect 519997 128555 520063 128558
rect 523200 128528 524400 128558
rect 117221 127938 117287 127941
rect 117221 127936 119140 127938
rect 117221 127880 117226 127936
rect 117282 127880 119140 127936
rect 117221 127878 119140 127880
rect 117221 127875 117287 127878
rect 519353 127530 519419 127533
rect 518788 127528 519419 127530
rect 518788 127472 519358 127528
rect 519414 127472 519419 127528
rect 518788 127470 519419 127472
rect 519353 127467 519419 127470
rect 519813 127122 519879 127125
rect 523200 127122 524400 127152
rect 519813 127120 524400 127122
rect 519813 127064 519818 127120
rect 519874 127064 524400 127120
rect 519813 127062 524400 127064
rect 519813 127059 519879 127062
rect 523200 127032 524400 127062
rect 520089 126170 520155 126173
rect 518788 126168 520155 126170
rect 518788 126112 520094 126168
rect 520150 126112 520155 126168
rect 518788 126110 520155 126112
rect 520089 126107 520155 126110
rect 116117 126034 116183 126037
rect 116117 126032 119140 126034
rect 116117 125976 116122 126032
rect 116178 125976 119140 126032
rect 116117 125974 119140 125976
rect 116117 125971 116183 125974
rect 519537 125626 519603 125629
rect 523200 125626 524400 125656
rect 519537 125624 524400 125626
rect 519537 125568 519542 125624
rect 519598 125568 524400 125624
rect 519537 125566 524400 125568
rect 519537 125563 519603 125566
rect 523200 125536 524400 125566
rect 519905 124810 519971 124813
rect 518788 124808 519971 124810
rect 518788 124752 519910 124808
rect 519966 124752 519971 124808
rect 518788 124750 519971 124752
rect 519905 124747 519971 124750
rect 116117 124130 116183 124133
rect 519353 124130 519419 124133
rect 523200 124130 524400 124160
rect 116117 124128 119140 124130
rect 116117 124072 116122 124128
rect 116178 124072 119140 124128
rect 116117 124070 119140 124072
rect 519353 124128 524400 124130
rect 519353 124072 519358 124128
rect 519414 124072 524400 124128
rect 519353 124070 524400 124072
rect 116117 124067 116183 124070
rect 519353 124067 519419 124070
rect 523200 124040 524400 124070
rect 520181 123450 520247 123453
rect 518788 123448 520247 123450
rect 518788 123392 520186 123448
rect 520242 123392 520247 123448
rect 518788 123390 520247 123392
rect 520181 123387 520247 123390
rect 519261 122634 519327 122637
rect 523200 122634 524400 122664
rect 519261 122632 524400 122634
rect 519261 122576 519266 122632
rect 519322 122576 524400 122632
rect 519261 122574 524400 122576
rect 519261 122571 519327 122574
rect 523200 122544 524400 122574
rect 115933 122226 115999 122229
rect 115933 122224 119140 122226
rect 115933 122168 115938 122224
rect 115994 122168 119140 122224
rect 115933 122166 119140 122168
rect 115933 122163 115999 122166
rect 519445 122090 519511 122093
rect 518788 122088 519511 122090
rect 518788 122032 519450 122088
rect 519506 122032 519511 122088
rect 518788 122030 519511 122032
rect 519445 122027 519511 122030
rect 113909 121410 113975 121413
rect 110860 121408 113975 121410
rect 110860 121352 113914 121408
rect 113970 121352 113975 121408
rect 110860 121350 113975 121352
rect 113909 121347 113975 121350
rect 519905 121138 519971 121141
rect 523200 121138 524400 121168
rect 519905 121136 524400 121138
rect 519905 121080 519910 121136
rect 519966 121080 524400 121136
rect 519905 121078 524400 121080
rect 519905 121075 519971 121078
rect 523200 121048 524400 121078
rect 519629 120730 519695 120733
rect 518788 120728 519695 120730
rect 518788 120672 519634 120728
rect 519690 120672 519695 120728
rect 518788 120670 519695 120672
rect 519629 120667 519695 120670
rect 116117 120186 116183 120189
rect 116117 120184 119140 120186
rect 116117 120128 116122 120184
rect 116178 120128 119140 120184
rect 116117 120126 119140 120128
rect 116117 120123 116183 120126
rect 520089 119642 520155 119645
rect 523200 119642 524400 119672
rect 520089 119640 524400 119642
rect 520089 119584 520094 119640
rect 520150 119584 524400 119640
rect 520089 119582 524400 119584
rect 520089 119579 520155 119582
rect 523200 119552 524400 119582
rect 519721 119370 519787 119373
rect 518788 119368 519787 119370
rect 518788 119312 519726 119368
rect 519782 119312 519787 119368
rect 518788 119310 519787 119312
rect 519721 119307 519787 119310
rect 116117 118282 116183 118285
rect 116117 118280 119140 118282
rect 116117 118224 116122 118280
rect 116178 118224 119140 118280
rect 116117 118222 119140 118224
rect 116117 118219 116183 118222
rect 520181 118146 520247 118149
rect 523200 118146 524400 118176
rect 520181 118144 524400 118146
rect 520181 118088 520186 118144
rect 520242 118088 524400 118144
rect 520181 118086 524400 118088
rect 520181 118083 520247 118086
rect 523200 118056 524400 118086
rect 519997 118010 520063 118013
rect 518788 118008 520063 118010
rect 518788 117952 520002 118008
rect 520058 117952 520063 118008
rect 518788 117950 520063 117952
rect 519997 117947 520063 117950
rect 519813 116650 519879 116653
rect 518788 116648 519879 116650
rect 518788 116592 519818 116648
rect 519874 116592 519879 116648
rect 518788 116590 519879 116592
rect 519813 116587 519879 116590
rect 519997 116514 520063 116517
rect 523200 116514 524400 116544
rect 519997 116512 524400 116514
rect 519997 116456 520002 116512
rect 520058 116456 524400 116512
rect 519997 116454 524400 116456
rect 519997 116451 520063 116454
rect 523200 116424 524400 116454
rect 116117 116378 116183 116381
rect 116117 116376 119140 116378
rect 116117 116320 116122 116376
rect 116178 116320 119140 116376
rect 116117 116318 119140 116320
rect 116117 116315 116183 116318
rect 519537 115290 519603 115293
rect 518788 115288 519603 115290
rect 518788 115232 519542 115288
rect 519598 115232 519603 115288
rect 518788 115230 519603 115232
rect 519537 115227 519603 115230
rect 519813 115018 519879 115021
rect 523200 115018 524400 115048
rect 519813 115016 524400 115018
rect 519813 114960 519818 115016
rect 519874 114960 524400 115016
rect 519813 114958 524400 114960
rect 519813 114955 519879 114958
rect 523200 114928 524400 114958
rect 116117 114474 116183 114477
rect 116117 114472 119140 114474
rect 116117 114416 116122 114472
rect 116178 114416 119140 114472
rect 116117 114414 119140 114416
rect 116117 114411 116183 114414
rect 519353 113930 519419 113933
rect 518788 113928 519419 113930
rect 518788 113872 519358 113928
rect 519414 113872 519419 113928
rect 518788 113870 519419 113872
rect 519353 113867 519419 113870
rect 519721 113522 519787 113525
rect 523200 113522 524400 113552
rect 519721 113520 524400 113522
rect 519721 113464 519726 113520
rect 519782 113464 524400 113520
rect 519721 113462 524400 113464
rect 519721 113459 519787 113462
rect 523200 113432 524400 113462
rect 115933 112570 115999 112573
rect 519261 112570 519327 112573
rect 115933 112568 119140 112570
rect 115933 112512 115938 112568
rect 115994 112512 119140 112568
rect 115933 112510 119140 112512
rect 518788 112568 519327 112570
rect 518788 112512 519266 112568
rect 519322 112512 519327 112568
rect 518788 112510 519327 112512
rect 115933 112507 115999 112510
rect 519261 112507 519327 112510
rect 519537 112026 519603 112029
rect 523200 112026 524400 112056
rect 519537 112024 524400 112026
rect 519537 111968 519542 112024
rect 519598 111968 524400 112024
rect 519537 111966 524400 111968
rect 519537 111963 519603 111966
rect 523200 111936 524400 111966
rect 519905 111210 519971 111213
rect 518788 111208 519971 111210
rect 518788 111152 519910 111208
rect 519966 111152 519971 111208
rect 518788 111150 519971 111152
rect 519905 111147 519971 111150
rect 116117 110666 116183 110669
rect 116117 110664 119140 110666
rect 116117 110608 116122 110664
rect 116178 110608 119140 110664
rect 116117 110606 119140 110608
rect 116117 110603 116183 110606
rect 519629 110530 519695 110533
rect 523200 110530 524400 110560
rect 519629 110528 524400 110530
rect 519629 110472 519634 110528
rect 519690 110472 524400 110528
rect 519629 110470 524400 110472
rect 519629 110467 519695 110470
rect 523200 110440 524400 110470
rect 114001 110122 114067 110125
rect 110860 110120 114067 110122
rect 110860 110064 114006 110120
rect 114062 110064 114067 110120
rect 110860 110062 114067 110064
rect 114001 110059 114067 110062
rect 520089 109850 520155 109853
rect 518788 109848 520155 109850
rect 518788 109792 520094 109848
rect 520150 109792 520155 109848
rect 518788 109790 520155 109792
rect 520089 109787 520155 109790
rect 520917 109034 520983 109037
rect 523200 109034 524400 109064
rect 520917 109032 524400 109034
rect 520917 108976 520922 109032
rect 520978 108976 524400 109032
rect 520917 108974 524400 108976
rect 520917 108971 520983 108974
rect 523200 108944 524400 108974
rect 116117 108762 116183 108765
rect 116117 108760 119140 108762
rect 116117 108704 116122 108760
rect 116178 108704 119140 108760
rect 116117 108702 119140 108704
rect 116117 108699 116183 108702
rect 520181 108490 520247 108493
rect 518788 108488 520247 108490
rect 518788 108432 520186 108488
rect 520242 108432 520247 108488
rect 518788 108430 520247 108432
rect 520181 108427 520247 108430
rect 521101 107538 521167 107541
rect 523200 107538 524400 107568
rect 521101 107536 524400 107538
rect 521101 107480 521106 107536
rect 521162 107480 524400 107536
rect 521101 107478 524400 107480
rect 521101 107475 521167 107478
rect 523200 107448 524400 107478
rect 519997 107130 520063 107133
rect 518788 107128 520063 107130
rect 518788 107072 520002 107128
rect 520058 107072 520063 107128
rect 518788 107070 520063 107072
rect 519997 107067 520063 107070
rect 110321 106314 110387 106317
rect 119110 106314 119170 106828
rect 110321 106312 119170 106314
rect 110321 106256 110326 106312
rect 110382 106256 119170 106312
rect 110321 106254 119170 106256
rect 110321 106251 110387 106254
rect 520273 106042 520339 106045
rect 523200 106042 524400 106072
rect 520273 106040 524400 106042
rect 520273 105984 520278 106040
rect 520334 105984 524400 106040
rect 520273 105982 524400 105984
rect 520273 105979 520339 105982
rect 523200 105952 524400 105982
rect 519813 105770 519879 105773
rect 518788 105768 519879 105770
rect 518788 105712 519818 105768
rect 519874 105712 519879 105768
rect 518788 105710 519879 105712
rect 519813 105707 519879 105710
rect 117129 104818 117195 104821
rect 117129 104816 119140 104818
rect 117129 104760 117134 104816
rect 117190 104760 119140 104816
rect 117129 104758 119140 104760
rect 117129 104755 117195 104758
rect 520825 104546 520891 104549
rect 523200 104546 524400 104576
rect 520825 104544 524400 104546
rect 520825 104488 520830 104544
rect 520886 104488 524400 104544
rect 520825 104486 524400 104488
rect 520825 104483 520891 104486
rect 523200 104456 524400 104486
rect 519721 104410 519787 104413
rect 518788 104408 519787 104410
rect 518788 104352 519726 104408
rect 519782 104352 519787 104408
rect 518788 104350 519787 104352
rect 519721 104347 519787 104350
rect 519537 103050 519603 103053
rect 518788 103048 519603 103050
rect 518788 102992 519542 103048
rect 519598 102992 519603 103048
rect 518788 102990 519603 102992
rect 519537 102987 519603 102990
rect 520733 103050 520799 103053
rect 523200 103050 524400 103080
rect 520733 103048 524400 103050
rect 520733 102992 520738 103048
rect 520794 102992 524400 103048
rect 520733 102990 524400 102992
rect 520733 102987 520799 102990
rect 523200 102960 524400 102990
rect 116945 102914 117011 102917
rect 116945 102912 119140 102914
rect 116945 102856 116950 102912
rect 117006 102856 119140 102912
rect 116945 102854 119140 102856
rect 116945 102851 117011 102854
rect 519629 101690 519695 101693
rect 518788 101688 519695 101690
rect 518788 101632 519634 101688
rect 519690 101632 519695 101688
rect 518788 101630 519695 101632
rect 519629 101627 519695 101630
rect 521009 101554 521075 101557
rect 523200 101554 524400 101584
rect 521009 101552 524400 101554
rect 521009 101496 521014 101552
rect 521070 101496 524400 101552
rect 521009 101494 524400 101496
rect 521009 101491 521075 101494
rect 523200 101464 524400 101494
rect 117037 101010 117103 101013
rect 117037 101008 119140 101010
rect 117037 100952 117042 101008
rect 117098 100952 119140 101008
rect 117037 100950 119140 100952
rect 117037 100947 117103 100950
rect 520917 100330 520983 100333
rect 518788 100328 520983 100330
rect 518788 100272 520922 100328
rect 520978 100272 520983 100328
rect 518788 100270 520983 100272
rect 520917 100267 520983 100270
rect 521193 100058 521259 100061
rect 523200 100058 524400 100088
rect 521193 100056 524400 100058
rect 521193 100000 521198 100056
rect 521254 100000 524400 100056
rect 521193 99998 524400 100000
rect 521193 99995 521259 99998
rect 523200 99968 524400 99998
rect 116853 99106 116919 99109
rect 116853 99104 119140 99106
rect 116853 99048 116858 99104
rect 116914 99048 119140 99104
rect 116853 99046 119140 99048
rect 116853 99043 116919 99046
rect 521101 98970 521167 98973
rect 518788 98968 521167 98970
rect 518788 98912 521106 98968
rect 521162 98912 521167 98968
rect 518788 98910 521167 98912
rect 521101 98907 521167 98910
rect 114093 98698 114159 98701
rect 110860 98696 114159 98698
rect 110860 98640 114098 98696
rect 114154 98640 114159 98696
rect 110860 98638 114159 98640
rect 114093 98635 114159 98638
rect 520917 98562 520983 98565
rect 523200 98562 524400 98592
rect 520917 98560 524400 98562
rect 520917 98504 520922 98560
rect 520978 98504 524400 98560
rect 520917 98502 524400 98504
rect 520917 98499 520983 98502
rect 523200 98472 524400 98502
rect 520273 97610 520339 97613
rect 518788 97608 520339 97610
rect 518788 97552 520278 97608
rect 520334 97552 520339 97608
rect 518788 97550 520339 97552
rect 520273 97547 520339 97550
rect 116761 97202 116827 97205
rect 116761 97200 119140 97202
rect 116761 97144 116766 97200
rect 116822 97144 119140 97200
rect 116761 97142 119140 97144
rect 116761 97139 116827 97142
rect 521377 97066 521443 97069
rect 523200 97066 524400 97096
rect 521377 97064 524400 97066
rect 521377 97008 521382 97064
rect 521438 97008 524400 97064
rect 521377 97006 524400 97008
rect 521377 97003 521443 97006
rect 523200 96976 524400 97006
rect 520825 96250 520891 96253
rect 518788 96248 520891 96250
rect 518788 96192 520830 96248
rect 520886 96192 520891 96248
rect 518788 96190 520891 96192
rect 520825 96187 520891 96190
rect 520273 95570 520339 95573
rect 523200 95570 524400 95600
rect 520273 95568 524400 95570
rect 520273 95512 520278 95568
rect 520334 95512 524400 95568
rect 520273 95510 524400 95512
rect 520273 95507 520339 95510
rect 523200 95480 524400 95510
rect 116669 95298 116735 95301
rect 116669 95296 119140 95298
rect 116669 95240 116674 95296
rect 116730 95240 119140 95296
rect 116669 95238 119140 95240
rect 116669 95235 116735 95238
rect 520733 94890 520799 94893
rect 518788 94888 520799 94890
rect 518788 94832 520738 94888
rect 520794 94832 520799 94888
rect 518788 94830 520799 94832
rect 520733 94827 520799 94830
rect 521101 93938 521167 93941
rect 523200 93938 524400 93968
rect 521101 93936 524400 93938
rect 521101 93880 521106 93936
rect 521162 93880 524400 93936
rect 521101 93878 524400 93880
rect 521101 93875 521167 93878
rect 523200 93848 524400 93878
rect 521009 93530 521075 93533
rect 518788 93528 521075 93530
rect 518788 93472 521014 93528
rect 521070 93472 521075 93528
rect 518788 93470 521075 93472
rect 521009 93467 521075 93470
rect 116577 93394 116643 93397
rect 116577 93392 119140 93394
rect 116577 93336 116582 93392
rect 116638 93336 119140 93392
rect 116577 93334 119140 93336
rect 116577 93331 116643 93334
rect 520181 92442 520247 92445
rect 523200 92442 524400 92472
rect 520181 92440 524400 92442
rect 520181 92384 520186 92440
rect 520242 92384 524400 92440
rect 520181 92382 524400 92384
rect 520181 92379 520247 92382
rect 523200 92352 524400 92382
rect 521193 92170 521259 92173
rect 518788 92168 521259 92170
rect 518788 92112 521198 92168
rect 521254 92112 521259 92168
rect 518788 92110 521259 92112
rect 521193 92107 521259 92110
rect 116117 91354 116183 91357
rect 116117 91352 119140 91354
rect 116117 91296 116122 91352
rect 116178 91296 119140 91352
rect 116117 91294 119140 91296
rect 116117 91291 116183 91294
rect 519997 90946 520063 90949
rect 523200 90946 524400 90976
rect 519997 90944 524400 90946
rect 519997 90888 520002 90944
rect 520058 90888 524400 90944
rect 519997 90886 524400 90888
rect 519997 90883 520063 90886
rect 523200 90856 524400 90886
rect 520917 90810 520983 90813
rect 518788 90808 520983 90810
rect 518788 90752 520922 90808
rect 520978 90752 520983 90808
rect 518788 90750 520983 90752
rect 520917 90747 520983 90750
rect 521377 89586 521443 89589
rect 518758 89584 521443 89586
rect 518758 89528 521382 89584
rect 521438 89528 521443 89584
rect 518758 89526 521443 89528
rect 116117 89450 116183 89453
rect 116117 89448 119140 89450
rect 116117 89392 116122 89448
rect 116178 89392 119140 89448
rect 518758 89420 518818 89526
rect 521377 89523 521443 89526
rect 519629 89450 519695 89453
rect 523200 89450 524400 89480
rect 519629 89448 524400 89450
rect 116117 89390 119140 89392
rect 519629 89392 519634 89448
rect 519690 89392 524400 89448
rect 519629 89390 524400 89392
rect 116117 89387 116183 89390
rect 519629 89387 519695 89390
rect 523200 89360 524400 89390
rect 520273 88090 520339 88093
rect 518788 88088 520339 88090
rect 518788 88032 520278 88088
rect 520334 88032 520339 88088
rect 518788 88030 520339 88032
rect 520273 88027 520339 88030
rect 519905 87954 519971 87957
rect 523200 87954 524400 87984
rect 519905 87952 524400 87954
rect 519905 87896 519910 87952
rect 519966 87896 524400 87952
rect 519905 87894 524400 87896
rect 519905 87891 519971 87894
rect 523200 87864 524400 87894
rect 116025 87546 116091 87549
rect 116025 87544 119140 87546
rect 116025 87488 116030 87544
rect 116086 87488 119140 87544
rect 116025 87486 119140 87488
rect 116025 87483 116091 87486
rect 114185 87274 114251 87277
rect 110860 87272 114251 87274
rect 110860 87216 114190 87272
rect 114246 87216 114251 87272
rect 110860 87214 114251 87216
rect 114185 87211 114251 87214
rect 521101 86730 521167 86733
rect 518788 86728 521167 86730
rect 518788 86672 521106 86728
rect 521162 86672 521167 86728
rect 518788 86670 521167 86672
rect 521101 86667 521167 86670
rect 519077 86458 519143 86461
rect 523200 86458 524400 86488
rect 519077 86456 524400 86458
rect 519077 86400 519082 86456
rect 519138 86400 524400 86456
rect 519077 86398 524400 86400
rect 519077 86395 519143 86398
rect 523200 86368 524400 86398
rect 115197 85642 115263 85645
rect 115197 85640 119140 85642
rect 115197 85584 115202 85640
rect 115258 85584 119140 85640
rect 115197 85582 119140 85584
rect 115197 85579 115263 85582
rect 520181 85370 520247 85373
rect 518788 85368 520247 85370
rect 518788 85312 520186 85368
rect 520242 85312 520247 85368
rect 518788 85310 520247 85312
rect 520181 85307 520247 85310
rect 519813 84962 519879 84965
rect 523200 84962 524400 84992
rect 519813 84960 524400 84962
rect 519813 84904 519818 84960
rect 519874 84904 524400 84960
rect 519813 84902 524400 84904
rect 519813 84899 519879 84902
rect 523200 84872 524400 84902
rect 519997 84010 520063 84013
rect 518788 84008 520063 84010
rect 518788 83952 520002 84008
rect 520058 83952 520063 84008
rect 518788 83950 520063 83952
rect 519997 83947 520063 83950
rect 116577 83738 116643 83741
rect 116577 83736 119140 83738
rect 116577 83680 116582 83736
rect 116638 83680 119140 83736
rect 116577 83678 119140 83680
rect 116577 83675 116643 83678
rect 520181 83466 520247 83469
rect 523200 83466 524400 83496
rect 520181 83464 524400 83466
rect 520181 83408 520186 83464
rect 520242 83408 524400 83464
rect 520181 83406 524400 83408
rect 520181 83403 520247 83406
rect 523200 83376 524400 83406
rect 519629 82650 519695 82653
rect 518788 82648 519695 82650
rect 518788 82592 519634 82648
rect 519690 82592 519695 82648
rect 518788 82590 519695 82592
rect 519629 82587 519695 82590
rect 519721 81970 519787 81973
rect 523200 81970 524400 82000
rect 519721 81968 524400 81970
rect 519721 81912 519726 81968
rect 519782 81912 524400 81968
rect 519721 81910 524400 81912
rect 519721 81907 519787 81910
rect 523200 81880 524400 81910
rect 116209 81834 116275 81837
rect 116209 81832 119140 81834
rect 116209 81776 116214 81832
rect 116270 81776 119140 81832
rect 116209 81774 119140 81776
rect 116209 81771 116275 81774
rect 519905 81290 519971 81293
rect 518788 81288 519971 81290
rect 518788 81232 519910 81288
rect 519966 81232 519971 81288
rect 518788 81230 519971 81232
rect 519905 81227 519971 81230
rect 519997 80474 520063 80477
rect 523200 80474 524400 80504
rect 519997 80472 524400 80474
rect 519997 80416 520002 80472
rect 520058 80416 524400 80472
rect 519997 80414 524400 80416
rect 519997 80411 520063 80414
rect 523200 80384 524400 80414
rect 115933 79930 115999 79933
rect 519077 79930 519143 79933
rect 115933 79928 119140 79930
rect 115933 79872 115938 79928
rect 115994 79872 119140 79928
rect 115933 79870 119140 79872
rect 518788 79928 519143 79930
rect 518788 79872 519082 79928
rect 519138 79872 519143 79928
rect 518788 79870 519143 79872
rect 115933 79867 115999 79870
rect 519077 79867 519143 79870
rect 519629 78978 519695 78981
rect 523200 78978 524400 79008
rect 519629 78976 524400 78978
rect 519629 78920 519634 78976
rect 519690 78920 524400 78976
rect 519629 78918 524400 78920
rect 519629 78915 519695 78918
rect 523200 78888 524400 78918
rect 519813 78570 519879 78573
rect 518788 78568 519879 78570
rect 518788 78512 519818 78568
rect 519874 78512 519879 78568
rect 518788 78510 519879 78512
rect 519813 78507 519879 78510
rect 116117 78026 116183 78029
rect 116117 78024 119140 78026
rect 116117 77968 116122 78024
rect 116178 77968 119140 78024
rect 116117 77966 119140 77968
rect 116117 77963 116183 77966
rect 519905 77482 519971 77485
rect 523200 77482 524400 77512
rect 519905 77480 524400 77482
rect 519905 77424 519910 77480
rect 519966 77424 524400 77480
rect 519905 77422 524400 77424
rect 519905 77419 519971 77422
rect 523200 77392 524400 77422
rect 520181 77210 520247 77213
rect 518788 77208 520247 77210
rect 518788 77152 520186 77208
rect 520242 77152 520247 77208
rect 518788 77150 520247 77152
rect 520181 77147 520247 77150
rect 519721 75986 519787 75989
rect 110860 75926 119140 75986
rect 518788 75984 519787 75986
rect 518788 75928 519726 75984
rect 519782 75928 519787 75984
rect 518788 75926 519787 75928
rect 519721 75923 519787 75926
rect 520181 75986 520247 75989
rect 523200 75986 524400 76016
rect 520181 75984 524400 75986
rect 520181 75928 520186 75984
rect 520242 75928 524400 75984
rect 520181 75926 524400 75928
rect 520181 75923 520247 75926
rect 523200 75896 524400 75926
rect 519997 74626 520063 74629
rect 518788 74624 520063 74626
rect 518788 74568 520002 74624
rect 520058 74568 520063 74624
rect 518788 74566 520063 74568
rect 519997 74563 520063 74566
rect 521009 74490 521075 74493
rect 523200 74490 524400 74520
rect 521009 74488 524400 74490
rect 521009 74432 521014 74488
rect 521070 74432 524400 74488
rect 521009 74430 524400 74432
rect 521009 74427 521075 74430
rect 523200 74400 524400 74430
rect 116669 74082 116735 74085
rect 116669 74080 119140 74082
rect 116669 74024 116674 74080
rect 116730 74024 119140 74080
rect 116669 74022 119140 74024
rect 116669 74019 116735 74022
rect 519629 73266 519695 73269
rect 518788 73264 519695 73266
rect 518788 73208 519634 73264
rect 519690 73208 519695 73264
rect 518788 73206 519695 73208
rect 519629 73203 519695 73206
rect 520917 72994 520983 72997
rect 523200 72994 524400 73024
rect 520917 72992 524400 72994
rect 520917 72936 520922 72992
rect 520978 72936 524400 72992
rect 520917 72934 524400 72936
rect 520917 72931 520983 72934
rect 523200 72904 524400 72934
rect 116577 72178 116643 72181
rect 116577 72176 119140 72178
rect 116577 72120 116582 72176
rect 116638 72120 119140 72176
rect 116577 72118 119140 72120
rect 116577 72115 116643 72118
rect 519905 71906 519971 71909
rect 518788 71904 519971 71906
rect 518788 71848 519910 71904
rect 519966 71848 519971 71904
rect 518788 71846 519971 71848
rect 519905 71843 519971 71846
rect 521193 71498 521259 71501
rect 523200 71498 524400 71528
rect 521193 71496 524400 71498
rect 521193 71440 521198 71496
rect 521254 71440 524400 71496
rect 521193 71438 524400 71440
rect 521193 71435 521259 71438
rect 523200 71408 524400 71438
rect 520181 70546 520247 70549
rect 518788 70544 520247 70546
rect 518788 70488 520186 70544
rect 520242 70488 520247 70544
rect 518788 70486 520247 70488
rect 520181 70483 520247 70486
rect 116301 70274 116367 70277
rect 116301 70272 119140 70274
rect 116301 70216 116306 70272
rect 116362 70216 119140 70272
rect 116301 70214 119140 70216
rect 116301 70211 116367 70214
rect 521101 69866 521167 69869
rect 523200 69866 524400 69896
rect 521101 69864 524400 69866
rect 521101 69808 521106 69864
rect 521162 69808 524400 69864
rect 521101 69806 524400 69808
rect 521101 69803 521167 69806
rect 523200 69776 524400 69806
rect 521009 69186 521075 69189
rect 518788 69184 521075 69186
rect 518788 69128 521014 69184
rect 521070 69128 521075 69184
rect 518788 69126 521075 69128
rect 521009 69123 521075 69126
rect 116117 68370 116183 68373
rect 521009 68370 521075 68373
rect 523200 68370 524400 68400
rect 116117 68368 119140 68370
rect 116117 68312 116122 68368
rect 116178 68312 119140 68368
rect 116117 68310 119140 68312
rect 521009 68368 524400 68370
rect 521009 68312 521014 68368
rect 521070 68312 524400 68368
rect 521009 68310 524400 68312
rect 116117 68307 116183 68310
rect 521009 68307 521075 68310
rect 523200 68280 524400 68310
rect 520917 67826 520983 67829
rect 518788 67824 520983 67826
rect 518788 67768 520922 67824
rect 520978 67768 520983 67824
rect 518788 67766 520983 67768
rect 520917 67763 520983 67766
rect 520457 66874 520523 66877
rect 523200 66874 524400 66904
rect 520457 66872 524400 66874
rect 520457 66816 520462 66872
rect 520518 66816 524400 66872
rect 520457 66814 524400 66816
rect 520457 66811 520523 66814
rect 523200 66784 524400 66814
rect 116577 66466 116643 66469
rect 521193 66466 521259 66469
rect 116577 66464 119140 66466
rect 116577 66408 116582 66464
rect 116638 66408 119140 66464
rect 116577 66406 119140 66408
rect 518788 66464 521259 66466
rect 518788 66408 521198 66464
rect 521254 66408 521259 66464
rect 518788 66406 521259 66408
rect 116577 66403 116643 66406
rect 521193 66403 521259 66406
rect 520365 65378 520431 65381
rect 523200 65378 524400 65408
rect 520365 65376 524400 65378
rect 520365 65320 520370 65376
rect 520426 65320 524400 65376
rect 520365 65318 524400 65320
rect 520365 65315 520431 65318
rect 523200 65288 524400 65318
rect 521101 65106 521167 65109
rect 518788 65104 521167 65106
rect 518788 65048 521106 65104
rect 521162 65048 521167 65104
rect 518788 65046 521167 65048
rect 521101 65043 521167 65046
rect 113357 64562 113423 64565
rect 110860 64560 113423 64562
rect 110860 64504 113362 64560
rect 113418 64504 113423 64560
rect 110860 64502 113423 64504
rect 113357 64499 113423 64502
rect 116209 64562 116275 64565
rect 116209 64560 119140 64562
rect 116209 64504 116214 64560
rect 116270 64504 119140 64560
rect 116209 64502 119140 64504
rect 116209 64499 116275 64502
rect 521101 63882 521167 63885
rect 523200 63882 524400 63912
rect 521101 63880 524400 63882
rect 521101 63824 521106 63880
rect 521162 63824 524400 63880
rect 521101 63822 524400 63824
rect 521101 63819 521167 63822
rect 523200 63792 524400 63822
rect 521009 63746 521075 63749
rect 518788 63744 521075 63746
rect 518788 63688 521014 63744
rect 521070 63688 521075 63744
rect 518788 63686 521075 63688
rect 521009 63683 521075 63686
rect 116117 62658 116183 62661
rect 116117 62656 119140 62658
rect 116117 62600 116122 62656
rect 116178 62600 119140 62656
rect 116117 62598 119140 62600
rect 116117 62595 116183 62598
rect 520457 62386 520523 62389
rect 518788 62384 520523 62386
rect 518788 62328 520462 62384
rect 520518 62328 520523 62384
rect 518788 62326 520523 62328
rect 520457 62323 520523 62326
rect 521009 62386 521075 62389
rect 523200 62386 524400 62416
rect 521009 62384 524400 62386
rect 521009 62328 521014 62384
rect 521070 62328 524400 62384
rect 521009 62326 524400 62328
rect 521009 62323 521075 62326
rect 523200 62296 524400 62326
rect 520365 61026 520431 61029
rect 518788 61024 520431 61026
rect 518788 60968 520370 61024
rect 520426 60968 520431 61024
rect 518788 60966 520431 60968
rect 520365 60963 520431 60966
rect 520733 60890 520799 60893
rect 523200 60890 524400 60920
rect 520733 60888 524400 60890
rect 520733 60832 520738 60888
rect 520794 60832 524400 60888
rect 520733 60830 524400 60832
rect 520733 60827 520799 60830
rect 523200 60800 524400 60830
rect 116577 60618 116643 60621
rect 116577 60616 119140 60618
rect 116577 60560 116582 60616
rect 116638 60560 119140 60616
rect 116577 60558 119140 60560
rect 116577 60555 116643 60558
rect 521101 59666 521167 59669
rect 518788 59664 521167 59666
rect 518788 59608 521106 59664
rect 521162 59608 521167 59664
rect 518788 59606 521167 59608
rect 521101 59603 521167 59606
rect 521101 59394 521167 59397
rect 523200 59394 524400 59424
rect 521101 59392 524400 59394
rect 521101 59336 521106 59392
rect 521162 59336 524400 59392
rect 521101 59334 524400 59336
rect 521101 59331 521167 59334
rect 523200 59304 524400 59334
rect 116761 58714 116827 58717
rect 116761 58712 119140 58714
rect 116761 58656 116766 58712
rect 116822 58656 119140 58712
rect 116761 58654 119140 58656
rect 116761 58651 116827 58654
rect 521009 58306 521075 58309
rect 518788 58304 521075 58306
rect 518788 58248 521014 58304
rect 521070 58248 521075 58304
rect 518788 58246 521075 58248
rect 521009 58243 521075 58246
rect 519905 57898 519971 57901
rect 523200 57898 524400 57928
rect 519905 57896 524400 57898
rect 519905 57840 519910 57896
rect 519966 57840 524400 57896
rect 519905 57838 524400 57840
rect 519905 57835 519971 57838
rect 523200 57808 524400 57838
rect 520733 56946 520799 56949
rect 518788 56944 520799 56946
rect 518788 56888 520738 56944
rect 520794 56888 520799 56944
rect 518788 56886 520799 56888
rect 520733 56883 520799 56886
rect 116669 56810 116735 56813
rect 116669 56808 119140 56810
rect 116669 56752 116674 56808
rect 116730 56752 119140 56808
rect 116669 56750 119140 56752
rect 116669 56747 116735 56750
rect 519813 56402 519879 56405
rect 523200 56402 524400 56432
rect 519813 56400 524400 56402
rect 519813 56344 519818 56400
rect 519874 56344 524400 56400
rect 519813 56342 524400 56344
rect 519813 56339 519879 56342
rect 523200 56312 524400 56342
rect 521101 55586 521167 55589
rect 518788 55584 521167 55586
rect 518788 55528 521106 55584
rect 521162 55528 521167 55584
rect 518788 55526 521167 55528
rect 521101 55523 521167 55526
rect 520181 54906 520247 54909
rect 523200 54906 524400 54936
rect 520181 54904 524400 54906
rect 110321 53954 110387 53957
rect 119110 53954 119170 54876
rect 520181 54848 520186 54904
rect 520242 54848 524400 54904
rect 520181 54846 524400 54848
rect 520181 54843 520247 54846
rect 523200 54816 524400 54846
rect 519905 54226 519971 54229
rect 518788 54224 519971 54226
rect 518788 54168 519910 54224
rect 519966 54168 519971 54224
rect 518788 54166 519971 54168
rect 519905 54163 519971 54166
rect 110321 53952 119170 53954
rect 110321 53896 110326 53952
rect 110382 53896 119170 53952
rect 110321 53894 119170 53896
rect 110321 53891 110387 53894
rect 519077 53410 519143 53413
rect 523200 53410 524400 53440
rect 519077 53408 524400 53410
rect 519077 53352 519082 53408
rect 519138 53352 524400 53408
rect 519077 53350 524400 53352
rect 519077 53347 519143 53350
rect 523200 53320 524400 53350
rect 114185 53138 114251 53141
rect 110860 53136 114251 53138
rect 110860 53080 114190 53136
rect 114246 53080 114251 53136
rect 110860 53078 114251 53080
rect 114185 53075 114251 53078
rect 110321 52594 110387 52597
rect 119110 52594 119170 52972
rect 519813 52866 519879 52869
rect 518788 52864 519879 52866
rect 518788 52808 519818 52864
rect 519874 52808 519879 52864
rect 518788 52806 519879 52808
rect 519813 52803 519879 52806
rect 110321 52592 119170 52594
rect 110321 52536 110326 52592
rect 110382 52536 119170 52592
rect 110321 52534 119170 52536
rect 110321 52531 110387 52534
rect 520089 51914 520155 51917
rect 523200 51914 524400 51944
rect 520089 51912 524400 51914
rect 520089 51856 520094 51912
rect 520150 51856 524400 51912
rect 520089 51854 524400 51856
rect 520089 51851 520155 51854
rect 523200 51824 524400 51854
rect 520181 51506 520247 51509
rect 518788 51504 520247 51506
rect 518788 51448 520186 51504
rect 520242 51448 520247 51504
rect 518788 51446 520247 51448
rect 520181 51443 520247 51446
rect 110321 51098 110387 51101
rect 110321 51096 119140 51098
rect 110321 51040 110326 51096
rect 110382 51040 119140 51096
rect 110321 51038 119140 51040
rect 110321 51035 110387 51038
rect 520181 50418 520247 50421
rect 523200 50418 524400 50448
rect 520181 50416 524400 50418
rect 520181 50360 520186 50416
rect 520242 50360 524400 50416
rect 520181 50358 524400 50360
rect 520181 50355 520247 50358
rect 523200 50328 524400 50358
rect 519077 50146 519143 50149
rect 518788 50144 519143 50146
rect 518788 50088 519082 50144
rect 519138 50088 519143 50144
rect 518788 50086 519143 50088
rect 519077 50083 519143 50086
rect 110321 48378 110387 48381
rect 119110 48378 119170 49164
rect 519077 48922 519143 48925
rect 523200 48922 524400 48952
rect 519077 48920 524400 48922
rect 519077 48864 519082 48920
rect 519138 48864 524400 48920
rect 519077 48862 524400 48864
rect 519077 48859 519143 48862
rect 523200 48832 524400 48862
rect 520089 48786 520155 48789
rect 518788 48784 520155 48786
rect 518788 48728 520094 48784
rect 520150 48728 520155 48784
rect 518788 48726 520155 48728
rect 520089 48723 520155 48726
rect 110321 48376 119170 48378
rect 110321 48320 110326 48376
rect 110382 48320 119170 48376
rect 110321 48318 119170 48320
rect 110321 48315 110387 48318
rect 520181 47426 520247 47429
rect 518788 47424 520247 47426
rect 518788 47368 520186 47424
rect 520242 47368 520247 47424
rect 518788 47366 520247 47368
rect 520181 47363 520247 47366
rect 519905 47290 519971 47293
rect 523200 47290 524400 47320
rect 519905 47288 524400 47290
rect 519905 47232 519910 47288
rect 519966 47232 524400 47288
rect 519905 47230 524400 47232
rect 519905 47227 519971 47230
rect 523200 47200 524400 47230
rect 110321 47154 110387 47157
rect 110321 47152 119140 47154
rect 110321 47096 110326 47152
rect 110382 47096 119140 47152
rect 110321 47094 119140 47096
rect 110321 47091 110387 47094
rect 519077 46066 519143 46069
rect 518788 46064 519143 46066
rect 518788 46008 519082 46064
rect 519138 46008 519143 46064
rect 518788 46006 519143 46008
rect 519077 46003 519143 46006
rect 519721 45794 519787 45797
rect 523200 45794 524400 45824
rect 519721 45792 524400 45794
rect 519721 45736 519726 45792
rect 519782 45736 524400 45792
rect 519721 45734 524400 45736
rect 519721 45731 519787 45734
rect 523200 45704 524400 45734
rect 110321 44298 110387 44301
rect 119110 44298 119170 45220
rect 519905 44706 519971 44709
rect 518788 44704 519971 44706
rect 518788 44648 519910 44704
rect 519966 44648 519971 44704
rect 518788 44646 519971 44648
rect 519905 44643 519971 44646
rect 110321 44296 119170 44298
rect 110321 44240 110326 44296
rect 110382 44240 119170 44296
rect 110321 44238 119170 44240
rect 520181 44298 520247 44301
rect 523200 44298 524400 44328
rect 520181 44296 524400 44298
rect 520181 44240 520186 44296
rect 520242 44240 524400 44296
rect 520181 44238 524400 44240
rect 110321 44235 110387 44238
rect 520181 44235 520247 44238
rect 523200 44208 524400 44238
rect 116117 43346 116183 43349
rect 519721 43346 519787 43349
rect 116117 43344 119140 43346
rect 116117 43288 116122 43344
rect 116178 43288 119140 43344
rect 116117 43286 119140 43288
rect 518788 43344 519787 43346
rect 518788 43288 519726 43344
rect 519782 43288 519787 43344
rect 518788 43286 519787 43288
rect 116117 43283 116183 43286
rect 519721 43283 519787 43286
rect 520733 42802 520799 42805
rect 523200 42802 524400 42832
rect 520733 42800 524400 42802
rect 520733 42744 520738 42800
rect 520794 42744 524400 42800
rect 520733 42742 524400 42744
rect 520733 42739 520799 42742
rect 523200 42712 524400 42742
rect 520181 41986 520247 41989
rect 518788 41984 520247 41986
rect 518788 41928 520186 41984
rect 520242 41928 520247 41984
rect 518788 41926 520247 41928
rect 520181 41923 520247 41926
rect 114093 41850 114159 41853
rect 110860 41848 114159 41850
rect 110860 41792 114098 41848
rect 114154 41792 114159 41848
rect 110860 41790 114159 41792
rect 114093 41787 114159 41790
rect 110321 41442 110387 41445
rect 110321 41440 119140 41442
rect 110321 41384 110326 41440
rect 110382 41384 119140 41440
rect 110321 41382 119140 41384
rect 110321 41379 110387 41382
rect 520733 41306 520799 41309
rect 518758 41304 520799 41306
rect 518758 41248 520738 41304
rect 520794 41248 520799 41304
rect 518758 41246 520799 41248
rect 518758 40596 518818 41246
rect 520733 41243 520799 41246
rect 520917 41306 520983 41309
rect 523200 41306 524400 41336
rect 520917 41304 524400 41306
rect 520917 41248 520922 41304
rect 520978 41248 524400 41304
rect 520917 41246 524400 41248
rect 520917 41243 520983 41246
rect 523200 41216 524400 41246
rect 520917 39946 520983 39949
rect 518758 39944 520983 39946
rect 518758 39888 520922 39944
rect 520978 39888 520983 39944
rect 518758 39886 520983 39888
rect 116945 39538 117011 39541
rect 116945 39536 119140 39538
rect 116945 39480 116950 39536
rect 117006 39480 119140 39536
rect 116945 39478 119140 39480
rect 116945 39475 117011 39478
rect 518758 39236 518818 39886
rect 520917 39883 520983 39886
rect 520917 39810 520983 39813
rect 523200 39810 524400 39840
rect 520917 39808 524400 39810
rect 520917 39752 520922 39808
rect 520978 39752 524400 39808
rect 520917 39750 524400 39752
rect 520917 39747 520983 39750
rect 523200 39720 524400 39750
rect 521101 38314 521167 38317
rect 523200 38314 524400 38344
rect 521101 38312 524400 38314
rect 521101 38256 521106 38312
rect 521162 38256 524400 38312
rect 521101 38254 524400 38256
rect 521101 38251 521167 38254
rect 523200 38224 524400 38254
rect 520917 37906 520983 37909
rect 518788 37904 520983 37906
rect 518788 37848 520922 37904
rect 520978 37848 520983 37904
rect 518788 37846 520983 37848
rect 520917 37843 520983 37846
rect 116853 37634 116919 37637
rect 116853 37632 119140 37634
rect 116853 37576 116858 37632
rect 116914 37576 119140 37632
rect 116853 37574 119140 37576
rect 116853 37571 116919 37574
rect 521101 37226 521167 37229
rect 518758 37224 521167 37226
rect 518758 37168 521106 37224
rect 521162 37168 521167 37224
rect 518758 37166 521167 37168
rect 518758 36516 518818 37166
rect 521101 37163 521167 37166
rect 521561 36818 521627 36821
rect 523200 36818 524400 36848
rect 521561 36816 524400 36818
rect 521561 36760 521566 36816
rect 521622 36760 524400 36816
rect 521561 36758 524400 36760
rect 521561 36755 521627 36758
rect 523200 36728 524400 36758
rect 521561 36002 521627 36005
rect 521561 36000 521670 36002
rect 521561 35944 521566 36000
rect 521622 35944 521670 36000
rect 521561 35939 521670 35944
rect 521610 35866 521670 35939
rect 518758 35806 521670 35866
rect 110321 34642 110387 34645
rect 119110 34642 119170 35700
rect 518758 35156 518818 35806
rect 520917 35322 520983 35325
rect 523200 35322 524400 35352
rect 520917 35320 524400 35322
rect 520917 35264 520922 35320
rect 520978 35264 524400 35320
rect 520917 35262 524400 35264
rect 520917 35259 520983 35262
rect 523200 35232 524400 35262
rect 110321 34640 119170 34642
rect 110321 34584 110326 34640
rect 110382 34584 119170 34640
rect 110321 34582 119170 34584
rect 110321 34579 110387 34582
rect 520917 34506 520983 34509
rect 518758 34504 520983 34506
rect 518758 34448 520922 34504
rect 520978 34448 520983 34504
rect 518758 34446 520983 34448
rect 117129 33826 117195 33829
rect 117129 33824 119140 33826
rect 117129 33768 117134 33824
rect 117190 33768 119140 33824
rect 518758 33796 518818 34446
rect 520917 34443 520983 34446
rect 521101 33826 521167 33829
rect 523200 33826 524400 33856
rect 521101 33824 524400 33826
rect 117129 33766 119140 33768
rect 521101 33768 521106 33824
rect 521162 33768 524400 33824
rect 521101 33766 524400 33768
rect 117129 33763 117195 33766
rect 521101 33763 521167 33766
rect 523200 33736 524400 33766
rect 521101 33146 521167 33149
rect 518758 33144 521167 33146
rect 518758 33088 521106 33144
rect 521162 33088 521167 33144
rect 518758 33086 521167 33088
rect 518758 32436 518818 33086
rect 521101 33083 521167 33086
rect 521101 32330 521167 32333
rect 523200 32330 524400 32360
rect 521101 32328 524400 32330
rect 521101 32272 521106 32328
rect 521162 32272 524400 32328
rect 521101 32270 524400 32272
rect 521101 32267 521167 32270
rect 523200 32240 524400 32270
rect 117037 31786 117103 31789
rect 117037 31784 119140 31786
rect 117037 31728 117042 31784
rect 117098 31728 119140 31784
rect 117037 31726 119140 31728
rect 117037 31723 117103 31726
rect 521101 31650 521167 31653
rect 518758 31648 521167 31650
rect 518758 31592 521106 31648
rect 521162 31592 521167 31648
rect 518758 31590 521167 31592
rect 518758 31076 518818 31590
rect 521101 31587 521167 31590
rect 523200 30834 524400 30864
rect 518850 30774 524400 30834
rect 114001 30426 114067 30429
rect 110860 30424 114067 30426
rect 110860 30368 114006 30424
rect 114062 30368 114067 30424
rect 110860 30366 114067 30368
rect 114001 30363 114067 30366
rect 518850 30290 518910 30774
rect 523200 30744 524400 30774
rect 518758 30230 518910 30290
rect 117221 29882 117287 29885
rect 117221 29880 119140 29882
rect 117221 29824 117226 29880
rect 117282 29824 119140 29880
rect 117221 29822 119140 29824
rect 117221 29819 117287 29822
rect 518758 29716 518818 30230
rect 520917 29338 520983 29341
rect 523200 29338 524400 29368
rect 520917 29336 524400 29338
rect 520917 29280 520922 29336
rect 520978 29280 524400 29336
rect 520917 29278 524400 29280
rect 520917 29275 520983 29278
rect 523200 29248 524400 29278
rect 520917 28386 520983 28389
rect 518788 28384 520983 28386
rect 518788 28328 520922 28384
rect 520978 28328 520983 28384
rect 518788 28326 520983 28328
rect 520917 28323 520983 28326
rect 116485 27978 116551 27981
rect 116485 27976 119140 27978
rect 116485 27920 116490 27976
rect 116546 27920 119140 27976
rect 116485 27918 119140 27920
rect 116485 27915 116551 27918
rect 523200 27842 524400 27872
rect 518850 27782 524400 27842
rect 518850 27570 518910 27782
rect 523200 27752 524400 27782
rect 518758 27510 518910 27570
rect 518758 26996 518818 27510
rect 523200 26346 524400 26376
rect 521610 26286 524400 26346
rect 521610 26210 521670 26286
rect 523200 26256 524400 26286
rect 518758 26150 521670 26210
rect 116301 26074 116367 26077
rect 116301 26072 119140 26074
rect 116301 26016 116306 26072
rect 116362 26016 119140 26072
rect 116301 26014 119140 26016
rect 116301 26011 116367 26014
rect 518758 25636 518818 26150
rect 521101 24850 521167 24853
rect 523200 24850 524400 24880
rect 521101 24848 524400 24850
rect 521101 24792 521106 24848
rect 521162 24792 524400 24848
rect 521101 24790 524400 24792
rect 521101 24787 521167 24790
rect 523200 24760 524400 24790
rect 116393 24170 116459 24173
rect 116393 24168 119140 24170
rect 116393 24112 116398 24168
rect 116454 24112 119140 24168
rect 116393 24110 119140 24112
rect 116393 24107 116459 24110
rect 518758 23626 518818 24276
rect 521101 23626 521167 23629
rect 518758 23624 521167 23626
rect 518758 23568 521106 23624
rect 521162 23568 521167 23624
rect 518758 23566 521167 23568
rect 521101 23563 521167 23566
rect 520365 23218 520431 23221
rect 523200 23218 524400 23248
rect 520365 23216 524400 23218
rect 520365 23160 520370 23216
rect 520426 23160 524400 23216
rect 520365 23158 524400 23160
rect 520365 23155 520431 23158
rect 523200 23128 524400 23158
rect 116209 22266 116275 22269
rect 518758 22266 518818 22916
rect 520365 22266 520431 22269
rect 116209 22264 119140 22266
rect 116209 22208 116214 22264
rect 116270 22208 119140 22264
rect 116209 22206 119140 22208
rect 518758 22264 520431 22266
rect 518758 22208 520370 22264
rect 520426 22208 520431 22264
rect 518758 22206 520431 22208
rect 116209 22203 116275 22206
rect 520365 22203 520431 22206
rect 520917 21722 520983 21725
rect 523200 21722 524400 21752
rect 520917 21720 524400 21722
rect 520917 21664 520922 21720
rect 520978 21664 524400 21720
rect 520917 21662 524400 21664
rect 520917 21659 520983 21662
rect 523200 21632 524400 21662
rect 518758 20906 518818 21556
rect 520917 20906 520983 20909
rect 518758 20904 520983 20906
rect 518758 20848 520922 20904
rect 520978 20848 520983 20904
rect 518758 20846 520983 20848
rect 520917 20843 520983 20846
rect 116025 20362 116091 20365
rect 116025 20360 119140 20362
rect 116025 20304 116030 20360
rect 116086 20304 119140 20360
rect 116025 20302 119140 20304
rect 116025 20299 116091 20302
rect 521101 20226 521167 20229
rect 523200 20226 524400 20256
rect 521101 20224 524400 20226
rect 518758 19546 518818 20196
rect 521101 20168 521106 20224
rect 521162 20168 524400 20224
rect 521101 20166 524400 20168
rect 521101 20163 521167 20166
rect 523200 20136 524400 20166
rect 521101 19546 521167 19549
rect 518758 19544 521167 19546
rect 518758 19488 521106 19544
rect 521162 19488 521167 19544
rect 518758 19486 521167 19488
rect 521101 19483 521167 19486
rect 113909 19002 113975 19005
rect 110860 19000 113975 19002
rect 110860 18944 113914 19000
rect 113970 18944 113975 19000
rect 110860 18942 113975 18944
rect 113909 18939 113975 18942
rect 116117 18458 116183 18461
rect 116117 18456 119140 18458
rect 116117 18400 116122 18456
rect 116178 18400 119140 18456
rect 116117 18398 119140 18400
rect 116117 18395 116183 18398
rect 518758 18186 518818 18836
rect 523200 18730 524400 18760
rect 521150 18670 524400 18730
rect 521150 18186 521210 18670
rect 523200 18640 524400 18670
rect 518758 18126 521210 18186
rect 518758 16826 518818 17476
rect 523200 17234 524400 17264
rect 521150 17174 524400 17234
rect 521150 16826 521210 17174
rect 523200 17144 524400 17174
rect 518758 16766 521210 16826
rect 115933 16418 115999 16421
rect 115933 16416 119140 16418
rect 115933 16360 115938 16416
rect 115994 16360 119140 16416
rect 115933 16358 119140 16360
rect 115933 16355 115999 16358
rect 518758 15466 518818 16116
rect 523200 15738 524400 15768
rect 521104 15678 524400 15738
rect 521104 15466 521164 15678
rect 523200 15648 524400 15678
rect 518758 15406 521164 15466
rect 116526 14452 116532 14516
rect 116596 14514 116602 14516
rect 116596 14454 119140 14514
rect 116596 14452 116602 14454
rect 518758 14106 518818 14756
rect 523200 14242 524400 14272
rect 521104 14182 524400 14242
rect 521104 14106 521164 14182
rect 523200 14152 524400 14182
rect 518758 14046 521164 14106
rect 518758 12746 518818 13396
rect 523200 12746 524400 12776
rect 518758 12686 524400 12746
rect 523200 12656 524400 12686
rect 116710 12548 116716 12612
rect 116780 12610 116786 12612
rect 116780 12550 119140 12610
rect 116780 12548 116786 12550
rect 518758 11386 518818 12036
rect 518758 11326 518910 11386
rect 518850 11250 518910 11326
rect 523200 11250 524400 11280
rect 518850 11190 524400 11250
rect 523200 11160 524400 11190
rect 116894 10644 116900 10708
rect 116964 10706 116970 10708
rect 116964 10646 119140 10706
rect 116964 10644 116970 10646
rect 518758 10026 518818 10676
rect 518758 9966 518910 10026
rect 518850 9754 518910 9966
rect 523200 9754 524400 9784
rect 518850 9694 524400 9754
rect 523200 9664 524400 9694
rect 521101 9346 521167 9349
rect 518788 9344 521167 9346
rect 518788 9288 521106 9344
rect 521162 9288 521167 9344
rect 518788 9286 521167 9288
rect 521101 9283 521167 9286
rect 117262 8740 117268 8804
rect 117332 8802 117338 8804
rect 117332 8742 119140 8802
rect 117332 8740 117338 8742
rect 110321 8394 110387 8397
rect 110505 8394 110571 8397
rect 110321 8392 110571 8394
rect 110321 8336 110326 8392
rect 110382 8336 110510 8392
rect 110566 8336 110571 8392
rect 110321 8334 110571 8336
rect 110321 8331 110387 8334
rect 110505 8331 110571 8334
rect 521101 8258 521167 8261
rect 523200 8258 524400 8288
rect 521101 8256 524400 8258
rect 521101 8200 521106 8256
rect 521162 8200 524400 8256
rect 521101 8198 524400 8200
rect 521101 8195 521167 8198
rect 523200 8168 524400 8198
rect 111057 7986 111123 7989
rect 116761 7986 116827 7989
rect 520365 7986 520431 7989
rect 111057 7984 116827 7986
rect 111057 7928 111062 7984
rect 111118 7928 116766 7984
rect 116822 7928 116827 7984
rect 111057 7926 116827 7928
rect 518788 7984 520431 7986
rect 518788 7928 520370 7984
rect 520426 7928 520431 7984
rect 518788 7926 520431 7928
rect 111057 7923 111123 7926
rect 116761 7923 116827 7926
rect 520365 7923 520431 7926
rect 113817 7714 113883 7717
rect 110860 7712 113883 7714
rect 110860 7656 113822 7712
rect 113878 7656 113883 7712
rect 110860 7654 113883 7656
rect 113817 7651 113883 7654
rect 117129 6898 117195 6901
rect 117129 6896 119140 6898
rect 117129 6840 117134 6896
rect 117190 6840 119140 6896
rect 117129 6838 119140 6840
rect 117129 6835 117195 6838
rect 520365 6762 520431 6765
rect 523200 6762 524400 6792
rect 520365 6760 524400 6762
rect 520365 6704 520370 6760
rect 520426 6704 524400 6760
rect 520365 6702 524400 6704
rect 520365 6699 520431 6702
rect 523200 6672 524400 6702
rect 521101 6626 521167 6629
rect 518788 6624 521167 6626
rect 518788 6568 521106 6624
rect 521162 6568 521167 6624
rect 518788 6566 521167 6568
rect 521101 6563 521167 6566
rect 110597 5674 110663 5677
rect 117037 5674 117103 5677
rect 110597 5672 117103 5674
rect 110597 5616 110602 5672
rect 110658 5616 117042 5672
rect 117098 5616 117103 5672
rect 110597 5614 117103 5616
rect 110597 5611 110663 5614
rect 117037 5611 117103 5614
rect 520917 5266 520983 5269
rect 518788 5264 520983 5266
rect 518788 5208 520922 5264
rect 520978 5208 520983 5264
rect 518788 5206 520983 5208
rect 520917 5203 520983 5206
rect 521101 5266 521167 5269
rect 523200 5266 524400 5296
rect 521101 5264 524400 5266
rect 521101 5208 521106 5264
rect 521162 5208 524400 5264
rect 521101 5206 524400 5208
rect 521101 5203 521167 5206
rect 523200 5176 524400 5206
rect 119110 4178 119170 4964
rect 110462 4118 119170 4178
rect 88290 3982 89730 4042
rect 88290 3906 88350 3982
rect 86910 3846 88350 3906
rect 89670 3906 89730 3982
rect 93810 3982 98194 4042
rect 93810 3906 93870 3982
rect 89670 3846 93870 3906
rect 96570 3846 98010 3906
rect 86910 3770 86970 3846
rect 74490 3710 80162 3770
rect 74490 3498 74550 3710
rect 55170 3438 59370 3498
rect 55170 3090 55230 3438
rect 45510 3030 55230 3090
rect 45510 2818 45570 3030
rect 32446 2758 45570 2818
rect 59310 2818 59370 3438
rect 68464 3438 74550 3498
rect 59310 2758 63234 2818
rect 32446 2685 32506 2758
rect 32397 2680 32506 2685
rect 32397 2624 32402 2680
rect 32458 2624 32506 2680
rect 32397 2622 32506 2624
rect 36353 2682 36419 2685
rect 62389 2682 62455 2685
rect 36353 2680 62455 2682
rect 36353 2624 36358 2680
rect 36414 2624 62394 2680
rect 62450 2624 62455 2680
rect 36353 2622 62455 2624
rect 63174 2682 63234 2758
rect 68464 2685 68524 3438
rect 68832 2758 78874 2818
rect 68832 2685 68892 2758
rect 64137 2682 64203 2685
rect 63174 2680 64203 2682
rect 63174 2624 64142 2680
rect 64198 2624 64203 2680
rect 63174 2622 64203 2624
rect 32397 2619 32463 2622
rect 36353 2619 36419 2622
rect 62389 2619 62455 2622
rect 64137 2619 64203 2622
rect 65333 2682 65399 2685
rect 68001 2682 68067 2685
rect 65333 2680 68067 2682
rect 65333 2624 65338 2680
rect 65394 2624 68006 2680
rect 68062 2624 68067 2680
rect 65333 2622 68067 2624
rect 65333 2619 65399 2622
rect 68001 2619 68067 2622
rect 68461 2680 68527 2685
rect 68461 2624 68466 2680
rect 68522 2624 68527 2680
rect 68461 2619 68527 2624
rect 68829 2680 68895 2685
rect 68829 2624 68834 2680
rect 68890 2624 68895 2680
rect 68829 2619 68895 2624
rect 69381 2682 69447 2685
rect 77017 2682 77083 2685
rect 69381 2680 77083 2682
rect 69381 2624 69386 2680
rect 69442 2624 77022 2680
rect 77078 2624 77083 2680
rect 69381 2622 77083 2624
rect 69381 2619 69447 2622
rect 77017 2619 77083 2622
rect 77247 2682 77313 2685
rect 77753 2682 77819 2685
rect 77247 2680 77819 2682
rect 77247 2624 77252 2680
rect 77308 2624 77758 2680
rect 77814 2624 77819 2680
rect 77247 2622 77819 2624
rect 78814 2682 78874 2758
rect 79961 2682 80027 2685
rect 78814 2680 80027 2682
rect 78814 2624 79966 2680
rect 80022 2624 80027 2680
rect 78814 2622 80027 2624
rect 80102 2682 80162 3710
rect 80470 3710 86970 3770
rect 80470 2685 80530 3710
rect 96570 3634 96630 3846
rect 95190 3574 96630 3634
rect 95190 3498 95250 3574
rect 88290 3438 89730 3498
rect 88290 3362 88350 3438
rect 86910 3302 88350 3362
rect 89670 3362 89730 3438
rect 92430 3438 95250 3498
rect 92430 3362 92490 3438
rect 89670 3302 92490 3362
rect 86910 3226 86970 3302
rect 80608 3166 86970 3226
rect 80608 2685 80668 3166
rect 84150 2894 95066 2954
rect 80237 2682 80303 2685
rect 80102 2680 80303 2682
rect 80102 2624 80242 2680
rect 80298 2624 80303 2680
rect 80102 2622 80303 2624
rect 77247 2619 77313 2622
rect 77753 2619 77819 2622
rect 79961 2619 80027 2622
rect 80237 2619 80303 2622
rect 80421 2680 80530 2685
rect 80421 2624 80426 2680
rect 80482 2624 80530 2680
rect 80421 2622 80530 2624
rect 80605 2680 80671 2685
rect 80605 2624 80610 2680
rect 80666 2624 80671 2680
rect 80421 2619 80487 2622
rect 80605 2619 80671 2624
rect 80789 2682 80855 2685
rect 84150 2682 84210 2894
rect 80789 2680 84210 2682
rect 80789 2624 80794 2680
rect 80850 2624 84210 2680
rect 80789 2622 84210 2624
rect 93025 2682 93091 2685
rect 94681 2682 94747 2685
rect 93025 2680 94747 2682
rect 93025 2624 93030 2680
rect 93086 2624 94686 2680
rect 94742 2624 94747 2680
rect 93025 2622 94747 2624
rect 95006 2682 95066 2894
rect 96337 2682 96403 2685
rect 95006 2680 96403 2682
rect 95006 2624 96342 2680
rect 96398 2624 96403 2680
rect 95006 2622 96403 2624
rect 97950 2682 98010 3846
rect 98134 3770 98194 3982
rect 100526 3982 100770 4042
rect 100526 3906 100586 3982
rect 98502 3846 100586 3906
rect 100710 3906 100770 3982
rect 109493 3906 109559 3909
rect 110045 3906 110111 3909
rect 100710 3846 102426 3906
rect 98502 3770 98562 3846
rect 98134 3710 98562 3770
rect 102366 3770 102426 3846
rect 109493 3904 110111 3906
rect 109493 3848 109498 3904
rect 109554 3848 110050 3904
rect 110106 3848 110111 3904
rect 109493 3846 110111 3848
rect 109493 3843 109559 3846
rect 110045 3843 110111 3846
rect 110229 3906 110295 3909
rect 110462 3906 110522 4118
rect 521009 3906 521075 3909
rect 110229 3904 110522 3906
rect 110229 3848 110234 3904
rect 110290 3848 110522 3904
rect 110229 3846 110522 3848
rect 518788 3904 521075 3906
rect 518788 3848 521014 3904
rect 521070 3848 521075 3904
rect 518788 3846 521075 3848
rect 110229 3843 110295 3846
rect 521009 3843 521075 3846
rect 520917 3770 520983 3773
rect 523200 3770 524400 3800
rect 102366 3710 110430 3770
rect 109677 3634 109743 3637
rect 101814 3632 109743 3634
rect 101814 3576 109682 3632
rect 109738 3576 109743 3632
rect 101814 3574 109743 3576
rect 110370 3634 110430 3710
rect 520917 3768 524400 3770
rect 520917 3712 520922 3768
rect 520978 3712 524400 3768
rect 520917 3710 524400 3712
rect 520917 3707 520983 3710
rect 523200 3680 524400 3710
rect 116301 3634 116367 3637
rect 110370 3632 116367 3634
rect 110370 3576 116306 3632
rect 116362 3576 116367 3632
rect 110370 3574 116367 3576
rect 101814 3498 101874 3574
rect 109677 3571 109743 3574
rect 116301 3571 116367 3574
rect 109493 3498 109559 3501
rect 110229 3498 110295 3501
rect 100710 3438 101874 3498
rect 102090 3438 102610 3498
rect 100109 2682 100175 2685
rect 100710 2682 100770 3438
rect 102090 3362 102150 3438
rect 101400 3302 102150 3362
rect 102550 3362 102610 3438
rect 109493 3496 110295 3498
rect 109493 3440 109498 3496
rect 109554 3440 110234 3496
rect 110290 3440 110295 3496
rect 109493 3438 110295 3440
rect 109493 3435 109559 3438
rect 110229 3435 110295 3438
rect 116945 3362 117011 3365
rect 102550 3360 117011 3362
rect 102550 3304 116950 3360
rect 117006 3304 117011 3360
rect 102550 3302 117011 3304
rect 101400 2818 101460 3302
rect 116945 3299 117011 3302
rect 110689 3226 110755 3229
rect 116669 3226 116735 3229
rect 102090 3224 110755 3226
rect 102090 3168 110694 3224
rect 110750 3168 110755 3224
rect 102090 3166 110755 3168
rect 102090 2954 102150 3166
rect 110689 3163 110755 3166
rect 113038 3224 116735 3226
rect 113038 3168 116674 3224
rect 116730 3168 116735 3224
rect 113038 3166 116735 3168
rect 113038 3090 113098 3166
rect 116669 3163 116735 3166
rect 97950 2622 100034 2682
rect 80789 2619 80855 2622
rect 93025 2619 93091 2622
rect 94681 2619 94747 2622
rect 96337 2619 96403 2622
rect 33041 2546 33107 2549
rect 94313 2546 94379 2549
rect 33041 2544 94379 2546
rect 33041 2488 33046 2544
rect 33102 2488 94318 2544
rect 94374 2488 94379 2544
rect 33041 2486 94379 2488
rect 33041 2483 33107 2486
rect 94313 2483 94379 2486
rect 96429 2546 96495 2549
rect 99833 2546 99899 2549
rect 96429 2544 99899 2546
rect 96429 2488 96434 2544
rect 96490 2488 99838 2544
rect 99894 2488 99899 2544
rect 96429 2486 99899 2488
rect 99974 2546 100034 2622
rect 100109 2680 100770 2682
rect 100109 2624 100114 2680
rect 100170 2624 100770 2680
rect 100109 2622 100770 2624
rect 101032 2758 101460 2818
rect 101998 2894 102150 2954
rect 103470 3030 113098 3090
rect 116301 3090 116367 3093
rect 116301 3088 119140 3090
rect 116301 3032 116306 3088
rect 116362 3032 119140 3088
rect 116301 3030 119140 3032
rect 100109 2619 100175 2622
rect 101032 2546 101092 2758
rect 101857 2682 101923 2685
rect 101998 2682 102058 2894
rect 103470 2685 103530 3030
rect 116301 3027 116367 3030
rect 111701 2954 111767 2957
rect 107610 2952 111767 2954
rect 107610 2896 111706 2952
rect 111762 2896 111767 2952
rect 107610 2894 111767 2896
rect 107610 2818 107670 2894
rect 111701 2891 111767 2894
rect 103838 2758 107670 2818
rect 109861 2818 109927 2821
rect 110597 2818 110663 2821
rect 109861 2816 110663 2818
rect 109861 2760 109866 2816
rect 109922 2760 110602 2816
rect 110658 2760 110663 2816
rect 109861 2758 110663 2760
rect 101857 2680 102058 2682
rect 101857 2624 101862 2680
rect 101918 2624 102058 2680
rect 101857 2622 102058 2624
rect 103421 2680 103530 2685
rect 103421 2624 103426 2680
rect 103482 2624 103530 2680
rect 103421 2622 103530 2624
rect 103605 2682 103671 2685
rect 103838 2682 103898 2758
rect 109861 2755 109927 2758
rect 110597 2755 110663 2758
rect 116209 2682 116275 2685
rect 521101 2682 521167 2685
rect 103605 2680 103898 2682
rect 103605 2624 103610 2680
rect 103666 2624 103898 2680
rect 103605 2622 103898 2624
rect 104022 2680 116275 2682
rect 104022 2624 116214 2680
rect 116270 2624 116275 2680
rect 104022 2622 116275 2624
rect 518788 2680 521167 2682
rect 518788 2624 521106 2680
rect 521162 2624 521167 2680
rect 518788 2622 521167 2624
rect 101857 2619 101923 2622
rect 103421 2619 103487 2622
rect 103605 2619 103671 2622
rect 99974 2486 101092 2546
rect 101489 2546 101555 2549
rect 104022 2546 104082 2622
rect 116209 2619 116275 2622
rect 521101 2619 521167 2622
rect 101489 2544 104082 2546
rect 101489 2488 101494 2544
rect 101550 2488 104082 2544
rect 101489 2486 104082 2488
rect 104157 2546 104223 2549
rect 116025 2546 116091 2549
rect 104157 2544 116091 2546
rect 104157 2488 104162 2544
rect 104218 2488 116030 2544
rect 116086 2488 116091 2544
rect 104157 2486 116091 2488
rect 96429 2483 96495 2486
rect 99833 2483 99899 2486
rect 101489 2483 101555 2486
rect 104157 2483 104223 2486
rect 116025 2483 116091 2486
rect 29545 2410 29611 2413
rect 100845 2410 100911 2413
rect 29545 2408 100911 2410
rect 29545 2352 29550 2408
rect 29606 2352 100850 2408
rect 100906 2352 100911 2408
rect 29545 2350 100911 2352
rect 29545 2347 29611 2350
rect 100845 2347 100911 2350
rect 101397 2410 101463 2413
rect 116117 2410 116183 2413
rect 101397 2408 116183 2410
rect 101397 2352 101402 2408
rect 101458 2352 116122 2408
rect 116178 2352 116183 2408
rect 101397 2350 116183 2352
rect 101397 2347 101463 2350
rect 116117 2347 116183 2350
rect 26049 2274 26115 2277
rect 115933 2274 115999 2277
rect 26049 2272 115999 2274
rect 26049 2216 26054 2272
rect 26110 2216 115938 2272
rect 115994 2216 115999 2272
rect 26049 2214 115999 2216
rect 26049 2211 26115 2214
rect 115933 2211 115999 2214
rect 521009 2274 521075 2277
rect 523200 2274 524400 2304
rect 521009 2272 524400 2274
rect 521009 2216 521014 2272
rect 521070 2216 524400 2272
rect 521009 2214 524400 2216
rect 521009 2211 521075 2214
rect 523200 2184 524400 2214
rect 22921 2138 22987 2141
rect 94129 2138 94195 2141
rect 22921 2136 94195 2138
rect 22921 2080 22926 2136
rect 22982 2080 94134 2136
rect 94190 2080 94195 2136
rect 22921 2078 94195 2080
rect 22921 2075 22987 2078
rect 94129 2075 94195 2078
rect 94313 2138 94379 2141
rect 96429 2138 96495 2141
rect 94313 2136 96495 2138
rect 94313 2080 94318 2136
rect 94374 2080 96434 2136
rect 96490 2080 96495 2136
rect 94313 2078 96495 2080
rect 94313 2075 94379 2078
rect 96429 2075 96495 2078
rect 96613 2138 96679 2141
rect 99649 2138 99715 2141
rect 96613 2136 99715 2138
rect 96613 2080 96618 2136
rect 96674 2080 99654 2136
rect 99710 2080 99715 2136
rect 96613 2078 99715 2080
rect 96613 2075 96679 2078
rect 99649 2075 99715 2078
rect 99833 2138 99899 2141
rect 104157 2138 104223 2141
rect 99833 2136 104223 2138
rect 99833 2080 99838 2136
rect 99894 2080 104162 2136
rect 104218 2080 104223 2136
rect 99833 2078 104223 2080
rect 99833 2075 99899 2078
rect 104157 2075 104223 2078
rect 104341 2138 104407 2141
rect 116526 2138 116532 2140
rect 104341 2136 116532 2138
rect 104341 2080 104346 2136
rect 104402 2080 116532 2136
rect 104341 2078 116532 2080
rect 104341 2075 104407 2078
rect 116526 2076 116532 2078
rect 116596 2076 116602 2140
rect 19609 2002 19675 2005
rect 100753 2002 100819 2005
rect 19609 2000 100819 2002
rect 19609 1944 19614 2000
rect 19670 1944 100758 2000
rect 100814 1944 100819 2000
rect 19609 1942 100819 1944
rect 19609 1939 19675 1942
rect 100753 1939 100819 1942
rect 101213 2002 101279 2005
rect 116710 2002 116716 2004
rect 101213 2000 116716 2002
rect 101213 1944 101218 2000
rect 101274 1944 116716 2000
rect 101213 1942 116716 1944
rect 101213 1939 101279 1942
rect 116710 1940 116716 1942
rect 116780 1940 116786 2004
rect 15929 1866 15995 1869
rect 116894 1866 116900 1868
rect 15929 1864 116900 1866
rect 15929 1808 15934 1864
rect 15990 1808 116900 1864
rect 15929 1806 116900 1808
rect 15929 1803 15995 1806
rect 116894 1804 116900 1806
rect 116964 1804 116970 1868
rect 5993 1730 6059 1733
rect 109493 1730 109559 1733
rect 5993 1728 109559 1730
rect 5993 1672 5998 1728
rect 6054 1672 109498 1728
rect 109554 1672 109559 1728
rect 5993 1670 109559 1672
rect 5993 1667 6059 1670
rect 109493 1667 109559 1670
rect 12617 1594 12683 1597
rect 117262 1594 117268 1596
rect 12617 1592 117268 1594
rect 12617 1536 12622 1592
rect 12678 1536 117268 1592
rect 12617 1534 117268 1536
rect 12617 1531 12683 1534
rect 117262 1532 117268 1534
rect 117332 1532 117338 1596
rect 229277 1594 229343 1597
rect 293585 1594 293651 1597
rect 229277 1592 293651 1594
rect 229277 1536 229282 1592
rect 229338 1536 293590 1592
rect 293646 1536 293651 1592
rect 229277 1534 293651 1536
rect 229277 1531 229343 1534
rect 293585 1531 293651 1534
rect 9305 1458 9371 1461
rect 117129 1458 117195 1461
rect 9305 1456 117195 1458
rect 9305 1400 9310 1456
rect 9366 1400 117134 1456
rect 117190 1400 117195 1456
rect 9305 1398 117195 1400
rect 9305 1395 9371 1398
rect 117129 1395 117195 1398
rect 163773 1458 163839 1461
rect 243629 1458 243695 1461
rect 163773 1456 243695 1458
rect 163773 1400 163778 1456
rect 163834 1400 243634 1456
rect 243690 1400 243695 1456
rect 163773 1398 243695 1400
rect 163773 1395 163839 1398
rect 243629 1395 243695 1398
rect 360285 1458 360351 1461
rect 393589 1458 393655 1461
rect 360285 1456 393655 1458
rect 360285 1400 360290 1456
rect 360346 1400 393594 1456
rect 393650 1400 393655 1456
rect 360285 1398 393655 1400
rect 360285 1395 360351 1398
rect 393589 1395 393655 1398
rect 85941 1322 86007 1325
rect 98269 1322 98335 1325
rect 103329 1322 103395 1325
rect 85941 1320 98194 1322
rect 85941 1264 85946 1320
rect 86002 1264 98194 1320
rect 85941 1262 98194 1264
rect 85941 1259 86007 1262
rect 98134 1186 98194 1262
rect 98269 1320 103395 1322
rect 98269 1264 98274 1320
rect 98330 1264 103334 1320
rect 103390 1264 103395 1320
rect 98269 1262 103395 1264
rect 98269 1259 98335 1262
rect 103329 1259 103395 1262
rect 108205 1322 108271 1325
rect 110413 1322 110479 1325
rect 108205 1320 110479 1322
rect 108205 1264 108210 1320
rect 108266 1264 110418 1320
rect 110474 1264 110479 1320
rect 108205 1262 110479 1264
rect 108205 1259 108271 1262
rect 110413 1259 110479 1262
rect 103421 1186 103487 1189
rect 98134 1184 103487 1186
rect 98134 1128 103426 1184
rect 103482 1128 103487 1184
rect 98134 1126 103487 1128
rect 103421 1123 103487 1126
rect 103881 1186 103947 1189
rect 108297 1186 108363 1189
rect 103881 1184 108363 1186
rect 103881 1128 103886 1184
rect 103942 1128 108302 1184
rect 108358 1128 108363 1184
rect 103881 1126 108363 1128
rect 103881 1123 103947 1126
rect 108297 1123 108363 1126
rect 95969 1050 96035 1053
rect 110045 1050 110111 1053
rect 95969 1048 110111 1050
rect 95969 992 95974 1048
rect 96030 992 110050 1048
rect 110106 992 110111 1048
rect 95969 990 110111 992
rect 95969 987 96035 990
rect 110045 987 110111 990
rect 89253 914 89319 917
rect 101489 914 101555 917
rect 89253 912 101555 914
rect 89253 856 89258 912
rect 89314 856 101494 912
rect 101550 856 101555 912
rect 89253 854 101555 856
rect 89253 851 89319 854
rect 101489 851 101555 854
rect 521101 778 521167 781
rect 523200 778 524400 808
rect 521101 776 524400 778
rect 521101 720 521106 776
rect 521162 720 524400 776
rect 521101 718 524400 720
rect 521101 715 521167 718
rect 523200 688 524400 718
<< via3 >>
rect 116532 14452 116596 14516
rect 116716 12548 116780 12612
rect 116900 10644 116964 10708
rect 117268 8740 117332 8804
rect 116532 2076 116596 2140
rect 116716 1940 116780 2004
rect 116900 1804 116964 1868
rect 117268 1532 117332 1596
<< metal4 >>
rect 1664 144454 1984 144496
rect 1664 144218 1706 144454
rect 1942 144218 1984 144454
rect 1664 144134 1984 144218
rect 1664 143898 1706 144134
rect 1942 143898 1984 144134
rect 1664 143856 1984 143898
rect 109956 144454 110276 144496
rect 109956 144218 109998 144454
rect 110234 144218 110276 144454
rect 109956 144134 110276 144218
rect 109956 143898 109998 144134
rect 110234 143898 110276 144134
rect 109956 143856 110276 143898
rect 119664 144454 119984 144496
rect 119664 144218 119706 144454
rect 119942 144218 119984 144454
rect 119664 144134 119984 144218
rect 119664 143898 119706 144134
rect 119942 143898 119984 144134
rect 119664 143856 119984 143898
rect 517940 144454 518260 144496
rect 517940 144218 517982 144454
rect 518218 144218 518260 144454
rect 517940 144134 518260 144218
rect 517940 143898 517982 144134
rect 518218 143898 518260 144134
rect 517940 143856 518260 143898
rect 1096 131454 1332 131496
rect 1096 131134 1332 131218
rect 1096 130856 1332 130898
rect 110616 131454 110936 131496
rect 110616 131218 110658 131454
rect 110894 131218 110936 131454
rect 110616 131134 110936 131218
rect 110616 130898 110658 131134
rect 110894 130898 110936 131134
rect 110616 130856 110936 130898
rect 119004 131454 119324 131496
rect 119004 131218 119046 131454
rect 119282 131218 119324 131454
rect 119004 131134 119324 131218
rect 119004 130898 119046 131134
rect 119282 130898 119324 131134
rect 119004 130856 119324 130898
rect 518600 131454 518920 131496
rect 518600 131218 518642 131454
rect 518878 131218 518920 131454
rect 518600 131134 518920 131218
rect 518600 130898 518642 131134
rect 518878 130898 518920 131134
rect 518600 130856 518920 130898
rect 1664 118454 1984 118496
rect 1664 118218 1706 118454
rect 1942 118218 1984 118454
rect 1664 118134 1984 118218
rect 1664 117898 1706 118134
rect 1942 117898 1984 118134
rect 1664 117856 1984 117898
rect 109956 118454 110276 118496
rect 109956 118218 109998 118454
rect 110234 118218 110276 118454
rect 109956 118134 110276 118218
rect 109956 117898 109998 118134
rect 110234 117898 110276 118134
rect 109956 117856 110276 117898
rect 119664 118454 119984 118496
rect 119664 118218 119706 118454
rect 119942 118218 119984 118454
rect 119664 118134 119984 118218
rect 119664 117898 119706 118134
rect 119942 117898 119984 118134
rect 119664 117856 119984 117898
rect 517940 118454 518260 118496
rect 517940 118218 517982 118454
rect 518218 118218 518260 118454
rect 517940 118134 518260 118218
rect 517940 117898 517982 118134
rect 518218 117898 518260 118134
rect 517940 117856 518260 117898
rect 1096 105454 1332 105496
rect 1096 105134 1332 105218
rect 1096 104856 1332 104898
rect 110616 105454 110936 105496
rect 110616 105218 110658 105454
rect 110894 105218 110936 105454
rect 110616 105134 110936 105218
rect 110616 104898 110658 105134
rect 110894 104898 110936 105134
rect 110616 104856 110936 104898
rect 119004 105454 119324 105496
rect 119004 105218 119046 105454
rect 119282 105218 119324 105454
rect 119004 105134 119324 105218
rect 119004 104898 119046 105134
rect 119282 104898 119324 105134
rect 119004 104856 119324 104898
rect 518600 105454 518920 105496
rect 518600 105218 518642 105454
rect 518878 105218 518920 105454
rect 518600 105134 518920 105218
rect 518600 104898 518642 105134
rect 518878 104898 518920 105134
rect 518600 104856 518920 104898
rect 1664 92454 1984 92496
rect 1664 92218 1706 92454
rect 1942 92218 1984 92454
rect 1664 92134 1984 92218
rect 1664 91898 1706 92134
rect 1942 91898 1984 92134
rect 1664 91856 1984 91898
rect 109956 92454 110276 92496
rect 109956 92218 109998 92454
rect 110234 92218 110276 92454
rect 109956 92134 110276 92218
rect 109956 91898 109998 92134
rect 110234 91898 110276 92134
rect 109956 91856 110276 91898
rect 119664 92454 119984 92496
rect 119664 92218 119706 92454
rect 119942 92218 119984 92454
rect 119664 92134 119984 92218
rect 119664 91898 119706 92134
rect 119942 91898 119984 92134
rect 119664 91856 119984 91898
rect 517940 92454 518260 92496
rect 517940 92218 517982 92454
rect 518218 92218 518260 92454
rect 517940 92134 518260 92218
rect 517940 91898 517982 92134
rect 518218 91898 518260 92134
rect 517940 91856 518260 91898
rect 1096 79454 1332 79496
rect 1096 79134 1332 79218
rect 1096 78856 1332 78898
rect 110616 79454 110936 79496
rect 110616 79218 110658 79454
rect 110894 79218 110936 79454
rect 110616 79134 110936 79218
rect 110616 78898 110658 79134
rect 110894 78898 110936 79134
rect 110616 78856 110936 78898
rect 119004 79454 119324 79496
rect 119004 79218 119046 79454
rect 119282 79218 119324 79454
rect 119004 79134 119324 79218
rect 119004 78898 119046 79134
rect 119282 78898 119324 79134
rect 119004 78856 119324 78898
rect 518600 79454 518920 79496
rect 518600 79218 518642 79454
rect 518878 79218 518920 79454
rect 518600 79134 518920 79218
rect 518600 78898 518642 79134
rect 518878 78898 518920 79134
rect 518600 78856 518920 78898
rect 1664 66454 1984 66496
rect 1664 66218 1706 66454
rect 1942 66218 1984 66454
rect 1664 66134 1984 66218
rect 1664 65898 1706 66134
rect 1942 65898 1984 66134
rect 1664 65856 1984 65898
rect 109956 66454 110276 66496
rect 109956 66218 109998 66454
rect 110234 66218 110276 66454
rect 109956 66134 110276 66218
rect 109956 65898 109998 66134
rect 110234 65898 110276 66134
rect 109956 65856 110276 65898
rect 119664 66454 119984 66496
rect 119664 66218 119706 66454
rect 119942 66218 119984 66454
rect 119664 66134 119984 66218
rect 119664 65898 119706 66134
rect 119942 65898 119984 66134
rect 119664 65856 119984 65898
rect 517940 66454 518260 66496
rect 517940 66218 517982 66454
rect 518218 66218 518260 66454
rect 517940 66134 518260 66218
rect 517940 65898 517982 66134
rect 518218 65898 518260 66134
rect 517940 65856 518260 65898
rect 1096 53454 1332 53496
rect 1096 53134 1332 53218
rect 1096 52856 1332 52898
rect 110616 53454 110936 53496
rect 110616 53218 110658 53454
rect 110894 53218 110936 53454
rect 110616 53134 110936 53218
rect 110616 52898 110658 53134
rect 110894 52898 110936 53134
rect 110616 52856 110936 52898
rect 119004 53454 119324 53496
rect 119004 53218 119046 53454
rect 119282 53218 119324 53454
rect 119004 53134 119324 53218
rect 119004 52898 119046 53134
rect 119282 52898 119324 53134
rect 119004 52856 119324 52898
rect 518600 53454 518920 53496
rect 518600 53218 518642 53454
rect 518878 53218 518920 53454
rect 518600 53134 518920 53218
rect 518600 52898 518642 53134
rect 518878 52898 518920 53134
rect 518600 52856 518920 52898
rect 1664 40454 1984 40496
rect 1664 40218 1706 40454
rect 1942 40218 1984 40454
rect 1664 40134 1984 40218
rect 1664 39898 1706 40134
rect 1942 39898 1984 40134
rect 1664 39856 1984 39898
rect 109956 40454 110276 40496
rect 109956 40218 109998 40454
rect 110234 40218 110276 40454
rect 109956 40134 110276 40218
rect 109956 39898 109998 40134
rect 110234 39898 110276 40134
rect 109956 39856 110276 39898
rect 119664 40454 119984 40496
rect 119664 40218 119706 40454
rect 119942 40218 119984 40454
rect 119664 40134 119984 40218
rect 119664 39898 119706 40134
rect 119942 39898 119984 40134
rect 119664 39856 119984 39898
rect 517940 40454 518260 40496
rect 517940 40218 517982 40454
rect 518218 40218 518260 40454
rect 517940 40134 518260 40218
rect 517940 39898 517982 40134
rect 518218 39898 518260 40134
rect 517940 39856 518260 39898
rect 1096 27454 1332 27496
rect 1096 27134 1332 27218
rect 1096 26856 1332 26898
rect 110616 27454 110936 27496
rect 110616 27218 110658 27454
rect 110894 27218 110936 27454
rect 110616 27134 110936 27218
rect 110616 26898 110658 27134
rect 110894 26898 110936 27134
rect 110616 26856 110936 26898
rect 119004 27454 119324 27496
rect 119004 27218 119046 27454
rect 119282 27218 119324 27454
rect 119004 27134 119324 27218
rect 119004 26898 119046 27134
rect 119282 26898 119324 27134
rect 119004 26856 119324 26898
rect 518600 27454 518920 27496
rect 518600 27218 518642 27454
rect 518878 27218 518920 27454
rect 518600 27134 518920 27218
rect 518600 26898 518642 27134
rect 518878 26898 518920 27134
rect 518600 26856 518920 26898
rect 116531 14516 116597 14517
rect 1664 14454 1984 14496
rect 1664 14218 1706 14454
rect 1942 14218 1984 14454
rect 1664 14134 1984 14218
rect 1664 13898 1706 14134
rect 1942 13898 1984 14134
rect 1664 13856 1984 13898
rect 109956 14454 110276 14496
rect 109956 14218 109998 14454
rect 110234 14218 110276 14454
rect 116531 14452 116532 14516
rect 116596 14452 116597 14516
rect 116531 14451 116597 14452
rect 119664 14454 119984 14496
rect 109956 14134 110276 14218
rect 109956 13898 109998 14134
rect 110234 13898 110276 14134
rect 109956 13856 110276 13898
rect 116534 2141 116594 14451
rect 119664 14218 119706 14454
rect 119942 14218 119984 14454
rect 119664 14134 119984 14218
rect 119664 13898 119706 14134
rect 119942 13898 119984 14134
rect 119664 13856 119984 13898
rect 517940 14454 518260 14496
rect 517940 14218 517982 14454
rect 518218 14218 518260 14454
rect 517940 14134 518260 14218
rect 517940 13898 517982 14134
rect 518218 13898 518260 14134
rect 517940 13856 518260 13898
rect 116715 12612 116781 12613
rect 116715 12548 116716 12612
rect 116780 12548 116781 12612
rect 116715 12547 116781 12548
rect 116531 2140 116597 2141
rect 116531 2076 116532 2140
rect 116596 2076 116597 2140
rect 116531 2075 116597 2076
rect 116718 2005 116778 12547
rect 116899 10708 116965 10709
rect 116899 10644 116900 10708
rect 116964 10644 116965 10708
rect 116899 10643 116965 10644
rect 116715 2004 116781 2005
rect 116715 1940 116716 2004
rect 116780 1940 116781 2004
rect 116715 1939 116781 1940
rect 116902 1869 116962 10643
rect 117267 8804 117333 8805
rect 117267 8740 117268 8804
rect 117332 8740 117333 8804
rect 117267 8739 117333 8740
rect 116899 1868 116965 1869
rect 116899 1804 116900 1868
rect 116964 1804 116965 1868
rect 116899 1803 116965 1804
rect 117270 1597 117330 8739
rect 117267 1596 117333 1597
rect 117267 1532 117268 1596
rect 117332 1532 117333 1596
rect 117267 1531 117333 1532
<< via4 >>
rect 1706 144218 1942 144454
rect 1706 143898 1942 144134
rect 109998 144218 110234 144454
rect 109998 143898 110234 144134
rect 119706 144218 119942 144454
rect 119706 143898 119942 144134
rect 517982 144218 518218 144454
rect 517982 143898 518218 144134
rect 1096 131218 1332 131454
rect 1096 130898 1332 131134
rect 110658 131218 110894 131454
rect 110658 130898 110894 131134
rect 119046 131218 119282 131454
rect 119046 130898 119282 131134
rect 518642 131218 518878 131454
rect 518642 130898 518878 131134
rect 1706 118218 1942 118454
rect 1706 117898 1942 118134
rect 109998 118218 110234 118454
rect 109998 117898 110234 118134
rect 119706 118218 119942 118454
rect 119706 117898 119942 118134
rect 517982 118218 518218 118454
rect 517982 117898 518218 118134
rect 1096 105218 1332 105454
rect 1096 104898 1332 105134
rect 110658 105218 110894 105454
rect 110658 104898 110894 105134
rect 119046 105218 119282 105454
rect 119046 104898 119282 105134
rect 518642 105218 518878 105454
rect 518642 104898 518878 105134
rect 1706 92218 1942 92454
rect 1706 91898 1942 92134
rect 109998 92218 110234 92454
rect 109998 91898 110234 92134
rect 119706 92218 119942 92454
rect 119706 91898 119942 92134
rect 517982 92218 518218 92454
rect 517982 91898 518218 92134
rect 1096 79218 1332 79454
rect 1096 78898 1332 79134
rect 110658 79218 110894 79454
rect 110658 78898 110894 79134
rect 119046 79218 119282 79454
rect 119046 78898 119282 79134
rect 518642 79218 518878 79454
rect 518642 78898 518878 79134
rect 1706 66218 1942 66454
rect 1706 65898 1942 66134
rect 109998 66218 110234 66454
rect 109998 65898 110234 66134
rect 119706 66218 119942 66454
rect 119706 65898 119942 66134
rect 517982 66218 518218 66454
rect 517982 65898 518218 66134
rect 1096 53218 1332 53454
rect 1096 52898 1332 53134
rect 110658 53218 110894 53454
rect 110658 52898 110894 53134
rect 119046 53218 119282 53454
rect 119046 52898 119282 53134
rect 518642 53218 518878 53454
rect 518642 52898 518878 53134
rect 1706 40218 1942 40454
rect 1706 39898 1942 40134
rect 109998 40218 110234 40454
rect 109998 39898 110234 40134
rect 119706 40218 119942 40454
rect 119706 39898 119942 40134
rect 517982 40218 518218 40454
rect 517982 39898 518218 40134
rect 1096 27218 1332 27454
rect 1096 26898 1332 27134
rect 110658 27218 110894 27454
rect 110658 26898 110894 27134
rect 119046 27218 119282 27454
rect 119046 26898 119282 27134
rect 518642 27218 518878 27454
rect 518642 26898 518878 27134
rect 1706 14218 1942 14454
rect 1706 13898 1942 14134
rect 109998 14218 110234 14454
rect 109998 13898 110234 14134
rect 119706 14218 119942 14454
rect 119706 13898 119942 14134
rect 517982 14218 518218 14454
rect 517982 13898 518218 14134
<< metal5 >>
rect 1104 156856 522836 157496
rect 1104 144454 2200 144496
rect 1104 144218 1706 144454
rect 1942 144218 2200 144454
rect 1104 144134 2200 144218
rect 1104 143898 1706 144134
rect 1942 143898 2200 144134
rect 1104 143856 2200 143898
rect 109800 144454 120200 144496
rect 109800 144218 109998 144454
rect 110234 144218 119706 144454
rect 119942 144218 120200 144454
rect 109800 144134 120200 144218
rect 109800 143898 109998 144134
rect 110234 143898 119706 144134
rect 119942 143898 120200 144134
rect 109800 143856 120200 143898
rect 517800 144454 522836 144496
rect 517800 144218 517982 144454
rect 518218 144218 522836 144454
rect 517800 144134 522836 144218
rect 517800 143898 517982 144134
rect 518218 143898 522836 144134
rect 517800 143856 522836 143898
rect 1072 131454 2200 131496
rect 1072 131218 1096 131454
rect 1332 131218 2200 131454
rect 1072 131134 2200 131218
rect 1072 130898 1096 131134
rect 1332 130898 2200 131134
rect 1072 130856 2200 130898
rect 109800 131454 120200 131496
rect 109800 131218 110658 131454
rect 110894 131218 119046 131454
rect 119282 131218 120200 131454
rect 109800 131134 120200 131218
rect 109800 130898 110658 131134
rect 110894 130898 119046 131134
rect 119282 130898 120200 131134
rect 109800 130856 120200 130898
rect 517800 131454 522836 131496
rect 517800 131218 518642 131454
rect 518878 131218 522836 131454
rect 517800 131134 522836 131218
rect 517800 130898 518642 131134
rect 518878 130898 522836 131134
rect 517800 130856 522836 130898
rect 1104 118454 2200 118496
rect 1104 118218 1706 118454
rect 1942 118218 2200 118454
rect 1104 118134 2200 118218
rect 1104 117898 1706 118134
rect 1942 117898 2200 118134
rect 1104 117856 2200 117898
rect 109800 118454 120200 118496
rect 109800 118218 109998 118454
rect 110234 118218 119706 118454
rect 119942 118218 120200 118454
rect 109800 118134 120200 118218
rect 109800 117898 109998 118134
rect 110234 117898 119706 118134
rect 119942 117898 120200 118134
rect 109800 117856 120200 117898
rect 517800 118454 522836 118496
rect 517800 118218 517982 118454
rect 518218 118218 522836 118454
rect 517800 118134 522836 118218
rect 517800 117898 517982 118134
rect 518218 117898 522836 118134
rect 517800 117856 522836 117898
rect 1072 105454 2200 105496
rect 1072 105218 1096 105454
rect 1332 105218 2200 105454
rect 1072 105134 2200 105218
rect 1072 104898 1096 105134
rect 1332 104898 2200 105134
rect 1072 104856 2200 104898
rect 109800 105454 120200 105496
rect 109800 105218 110658 105454
rect 110894 105218 119046 105454
rect 119282 105218 120200 105454
rect 109800 105134 120200 105218
rect 109800 104898 110658 105134
rect 110894 104898 119046 105134
rect 119282 104898 120200 105134
rect 109800 104856 120200 104898
rect 517800 105454 522836 105496
rect 517800 105218 518642 105454
rect 518878 105218 522836 105454
rect 517800 105134 522836 105218
rect 517800 104898 518642 105134
rect 518878 104898 522836 105134
rect 517800 104856 522836 104898
rect 1104 92454 2200 92496
rect 1104 92218 1706 92454
rect 1942 92218 2200 92454
rect 1104 92134 2200 92218
rect 1104 91898 1706 92134
rect 1942 91898 2200 92134
rect 1104 91856 2200 91898
rect 109800 92454 120200 92496
rect 109800 92218 109998 92454
rect 110234 92218 119706 92454
rect 119942 92218 120200 92454
rect 109800 92134 120200 92218
rect 109800 91898 109998 92134
rect 110234 91898 119706 92134
rect 119942 91898 120200 92134
rect 109800 91856 120200 91898
rect 517800 92454 522836 92496
rect 517800 92218 517982 92454
rect 518218 92218 522836 92454
rect 517800 92134 522836 92218
rect 517800 91898 517982 92134
rect 518218 91898 522836 92134
rect 517800 91856 522836 91898
rect 1072 79454 2200 79496
rect 1072 79218 1096 79454
rect 1332 79218 2200 79454
rect 1072 79134 2200 79218
rect 1072 78898 1096 79134
rect 1332 78898 2200 79134
rect 1072 78856 2200 78898
rect 109800 79454 120200 79496
rect 109800 79218 110658 79454
rect 110894 79218 119046 79454
rect 119282 79218 120200 79454
rect 109800 79134 120200 79218
rect 109800 78898 110658 79134
rect 110894 78898 119046 79134
rect 119282 78898 120200 79134
rect 109800 78856 120200 78898
rect 517800 79454 522836 79496
rect 517800 79218 518642 79454
rect 518878 79218 522836 79454
rect 517800 79134 522836 79218
rect 517800 78898 518642 79134
rect 518878 78898 522836 79134
rect 517800 78856 522836 78898
rect 1104 66454 2200 66496
rect 1104 66218 1706 66454
rect 1942 66218 2200 66454
rect 1104 66134 2200 66218
rect 1104 65898 1706 66134
rect 1942 65898 2200 66134
rect 1104 65856 2200 65898
rect 109800 66454 120200 66496
rect 109800 66218 109998 66454
rect 110234 66218 119706 66454
rect 119942 66218 120200 66454
rect 109800 66134 120200 66218
rect 109800 65898 109998 66134
rect 110234 65898 119706 66134
rect 119942 65898 120200 66134
rect 109800 65856 120200 65898
rect 517800 66454 522836 66496
rect 517800 66218 517982 66454
rect 518218 66218 522836 66454
rect 517800 66134 522836 66218
rect 517800 65898 517982 66134
rect 518218 65898 522836 66134
rect 517800 65856 522836 65898
rect 1072 53454 2200 53496
rect 1072 53218 1096 53454
rect 1332 53218 2200 53454
rect 1072 53134 2200 53218
rect 1072 52898 1096 53134
rect 1332 52898 2200 53134
rect 1072 52856 2200 52898
rect 109800 53454 120200 53496
rect 109800 53218 110658 53454
rect 110894 53218 119046 53454
rect 119282 53218 120200 53454
rect 109800 53134 120200 53218
rect 109800 52898 110658 53134
rect 110894 52898 119046 53134
rect 119282 52898 120200 53134
rect 109800 52856 120200 52898
rect 517800 53454 522836 53496
rect 517800 53218 518642 53454
rect 518878 53218 522836 53454
rect 517800 53134 522836 53218
rect 517800 52898 518642 53134
rect 518878 52898 522836 53134
rect 517800 52856 522836 52898
rect 1104 40454 2200 40496
rect 1104 40218 1706 40454
rect 1942 40218 2200 40454
rect 1104 40134 2200 40218
rect 1104 39898 1706 40134
rect 1942 39898 2200 40134
rect 1104 39856 2200 39898
rect 109800 40454 120200 40496
rect 109800 40218 109998 40454
rect 110234 40218 119706 40454
rect 119942 40218 120200 40454
rect 109800 40134 120200 40218
rect 109800 39898 109998 40134
rect 110234 39898 119706 40134
rect 119942 39898 120200 40134
rect 109800 39856 120200 39898
rect 517800 40454 522836 40496
rect 517800 40218 517982 40454
rect 518218 40218 522836 40454
rect 517800 40134 522836 40218
rect 517800 39898 517982 40134
rect 518218 39898 522836 40134
rect 517800 39856 522836 39898
rect 1072 27454 2200 27496
rect 1072 27218 1096 27454
rect 1332 27218 2200 27454
rect 1072 27134 2200 27218
rect 1072 26898 1096 27134
rect 1332 26898 2200 27134
rect 1072 26856 2200 26898
rect 109800 27454 120200 27496
rect 109800 27218 110658 27454
rect 110894 27218 119046 27454
rect 119282 27218 120200 27454
rect 109800 27134 120200 27218
rect 109800 26898 110658 27134
rect 110894 26898 119046 27134
rect 119282 26898 120200 27134
rect 109800 26856 120200 26898
rect 517800 27454 522836 27496
rect 517800 27218 518642 27454
rect 518878 27218 522836 27454
rect 517800 27134 522836 27218
rect 517800 26898 518642 27134
rect 518878 26898 522836 27134
rect 517800 26856 522836 26898
rect 1104 14454 2200 14496
rect 1104 14218 1706 14454
rect 1942 14218 2200 14454
rect 1104 14134 2200 14218
rect 1104 13898 1706 14134
rect 1942 13898 2200 14134
rect 1104 13856 2200 13898
rect 109800 14454 120200 14496
rect 109800 14218 109998 14454
rect 110234 14218 119706 14454
rect 119942 14218 120200 14454
rect 109800 14134 120200 14218
rect 109800 13898 109998 14134
rect 110234 13898 119706 14134
rect 119942 13898 120200 14134
rect 109800 13856 120200 13898
rect 517800 14454 522836 14496
rect 517800 14218 517982 14454
rect 518218 14218 522836 14454
rect 517800 14134 522836 14218
rect 517800 13898 517982 14134
rect 518218 13898 522836 14134
rect 517800 13856 522836 13898
use mgmt_core  core
timestamp 1638474025
transform 1 0 119000 0 1 2000
box 0 0 400000 148000
use DFFRAM  DFFRAM
timestamp 1638474025
transform 1 0 1000 0 1 2000
box 4 0 110000 148000
<< labels >>
rlabel metal5 s 1104 26856 2200 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 26856 120200 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 26856 522836 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 52856 2200 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 52856 120200 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 52856 522836 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 78856 2200 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 78856 120200 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 78856 522836 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 104856 2200 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 104856 120200 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 104856 522836 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 130856 2200 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 130856 120200 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 130856 522836 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 156856 522836 157496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 13856 2200 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 13856 120200 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 13856 522836 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 39856 2200 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 39856 120200 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 39856 522836 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 65856 2200 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 65856 120200 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 65856 522836 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 91856 2200 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 91856 120200 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 91856 522836 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 117856 2200 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 117856 120200 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 117856 522836 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 143856 2200 144496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 143856 120200 144496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 143856 522836 144496 6 VPWR
port 1 nsew power input
rlabel metal2 s 294786 -400 294842 800 6 core_clk
port 2 nsew signal input
rlabel metal2 s 98274 -400 98330 800 6 core_rstn
port 3 nsew signal input
rlabel metal3 s 523200 63792 524400 63912 6 debug_in
port 4 nsew signal input
rlabel metal3 s 523200 65288 524400 65408 6 debug_mode
port 5 nsew signal tristate
rlabel metal3 s 523200 66784 524400 66904 6 debug_oeb
port 6 nsew signal tristate
rlabel metal3 s 523200 68280 524400 68400 6 debug_out
port 7 nsew signal tristate
rlabel metal3 s 523200 145120 524400 145240 6 flash_clk
port 8 nsew signal tristate
rlabel metal3 s 523200 143624 524400 143744 6 flash_csb
port 9 nsew signal tristate
rlabel metal3 s 523200 146616 524400 146736 6 flash_io0_di
port 10 nsew signal input
rlabel metal3 s 523200 148112 524400 148232 6 flash_io0_do
port 11 nsew signal tristate
rlabel metal3 s 523200 149608 524400 149728 6 flash_io0_oeb
port 12 nsew signal tristate
rlabel metal3 s 523200 151104 524400 151224 6 flash_io1_di
port 13 nsew signal input
rlabel metal3 s 523200 152600 524400 152720 6 flash_io1_do
port 14 nsew signal tristate
rlabel metal3 s 523200 154096 524400 154216 6 flash_io1_oeb
port 15 nsew signal tristate
rlabel metal3 s 523200 155592 524400 155712 6 flash_io2_di
port 16 nsew signal input
rlabel metal3 s 523200 157088 524400 157208 6 flash_io2_do
port 17 nsew signal tristate
rlabel metal3 s 523200 158584 524400 158704 6 flash_io2_oeb
port 18 nsew signal tristate
rlabel metal3 s 523200 160080 524400 160200 6 flash_io3_di
port 19 nsew signal input
rlabel metal3 s 523200 161576 524400 161696 6 flash_io3_do
port 20 nsew signal tristate
rlabel metal3 s 523200 163072 524400 163192 6 flash_io3_oeb
port 21 nsew signal tristate
rlabel metal2 s 32770 -400 32826 800 6 gpio_in_pad
port 22 nsew signal input
rlabel metal2 s 163778 -400 163834 800 6 gpio_inenb_pad
port 23 nsew signal tristate
rlabel metal2 s 229282 -400 229338 800 6 gpio_mode0_pad
port 24 nsew signal tristate
rlabel metal2 s 360290 -400 360346 800 6 gpio_mode1_pad
port 25 nsew signal tristate
rlabel metal2 s 425794 -400 425850 800 6 gpio_out_pad
port 26 nsew signal tristate
rlabel metal2 s 491298 -400 491354 800 6 gpio_outenb_pad
port 27 nsew signal tristate
rlabel metal3 s 523200 90856 524400 90976 6 hk_ack_i
port 28 nsew signal input
rlabel metal3 s 523200 93848 524400 93968 6 hk_cyc_o
port 29 nsew signal tristate
rlabel metal3 s 523200 95480 524400 95600 6 hk_dat_i[0]
port 30 nsew signal input
rlabel metal3 s 523200 110440 524400 110560 6 hk_dat_i[10]
port 31 nsew signal input
rlabel metal3 s 523200 111936 524400 112056 6 hk_dat_i[11]
port 32 nsew signal input
rlabel metal3 s 523200 113432 524400 113552 6 hk_dat_i[12]
port 33 nsew signal input
rlabel metal3 s 523200 114928 524400 115048 6 hk_dat_i[13]
port 34 nsew signal input
rlabel metal3 s 523200 116424 524400 116544 6 hk_dat_i[14]
port 35 nsew signal input
rlabel metal3 s 523200 118056 524400 118176 6 hk_dat_i[15]
port 36 nsew signal input
rlabel metal3 s 523200 119552 524400 119672 6 hk_dat_i[16]
port 37 nsew signal input
rlabel metal3 s 523200 121048 524400 121168 6 hk_dat_i[17]
port 38 nsew signal input
rlabel metal3 s 523200 122544 524400 122664 6 hk_dat_i[18]
port 39 nsew signal input
rlabel metal3 s 523200 124040 524400 124160 6 hk_dat_i[19]
port 40 nsew signal input
rlabel metal3 s 523200 96976 524400 97096 6 hk_dat_i[1]
port 41 nsew signal input
rlabel metal3 s 523200 125536 524400 125656 6 hk_dat_i[20]
port 42 nsew signal input
rlabel metal3 s 523200 127032 524400 127152 6 hk_dat_i[21]
port 43 nsew signal input
rlabel metal3 s 523200 128528 524400 128648 6 hk_dat_i[22]
port 44 nsew signal input
rlabel metal3 s 523200 130024 524400 130144 6 hk_dat_i[23]
port 45 nsew signal input
rlabel metal3 s 523200 131520 524400 131640 6 hk_dat_i[24]
port 46 nsew signal input
rlabel metal3 s 523200 133016 524400 133136 6 hk_dat_i[25]
port 47 nsew signal input
rlabel metal3 s 523200 134512 524400 134632 6 hk_dat_i[26]
port 48 nsew signal input
rlabel metal3 s 523200 136008 524400 136128 6 hk_dat_i[27]
port 49 nsew signal input
rlabel metal3 s 523200 137504 524400 137624 6 hk_dat_i[28]
port 50 nsew signal input
rlabel metal3 s 523200 139000 524400 139120 6 hk_dat_i[29]
port 51 nsew signal input
rlabel metal3 s 523200 98472 524400 98592 6 hk_dat_i[2]
port 52 nsew signal input
rlabel metal3 s 523200 140496 524400 140616 6 hk_dat_i[30]
port 53 nsew signal input
rlabel metal3 s 523200 142128 524400 142248 6 hk_dat_i[31]
port 54 nsew signal input
rlabel metal3 s 523200 99968 524400 100088 6 hk_dat_i[3]
port 55 nsew signal input
rlabel metal3 s 523200 101464 524400 101584 6 hk_dat_i[4]
port 56 nsew signal input
rlabel metal3 s 523200 102960 524400 103080 6 hk_dat_i[5]
port 57 nsew signal input
rlabel metal3 s 523200 104456 524400 104576 6 hk_dat_i[6]
port 58 nsew signal input
rlabel metal3 s 523200 105952 524400 106072 6 hk_dat_i[7]
port 59 nsew signal input
rlabel metal3 s 523200 107448 524400 107568 6 hk_dat_i[8]
port 60 nsew signal input
rlabel metal3 s 523200 108944 524400 109064 6 hk_dat_i[9]
port 61 nsew signal input
rlabel metal3 s 523200 92352 524400 92472 6 hk_stb_o
port 62 nsew signal tristate
rlabel metal2 s 521842 163200 521898 164400 6 irq[0]
port 63 nsew signal input
rlabel metal2 s 522670 163200 522726 164400 6 irq[1]
port 64 nsew signal input
rlabel metal2 s 523498 163200 523554 164400 6 irq[2]
port 65 nsew signal input
rlabel metal3 s 523200 74400 524400 74520 6 irq[3]
port 66 nsew signal input
rlabel metal3 s 523200 72904 524400 73024 6 irq[4]
port 67 nsew signal input
rlabel metal3 s 523200 71408 524400 71528 6 irq[5]
port 68 nsew signal input
rlabel metal2 s 386 163200 442 164400 6 la_iena[0]
port 69 nsew signal tristate
rlabel metal2 s 336830 163200 336886 164400 6 la_iena[100]
port 70 nsew signal tristate
rlabel metal2 s 340142 163200 340198 164400 6 la_iena[101]
port 71 nsew signal tristate
rlabel metal2 s 343546 163200 343602 164400 6 la_iena[102]
port 72 nsew signal tristate
rlabel metal2 s 346858 163200 346914 164400 6 la_iena[103]
port 73 nsew signal tristate
rlabel metal2 s 350262 163200 350318 164400 6 la_iena[104]
port 74 nsew signal tristate
rlabel metal2 s 353666 163200 353722 164400 6 la_iena[105]
port 75 nsew signal tristate
rlabel metal2 s 356978 163200 357034 164400 6 la_iena[106]
port 76 nsew signal tristate
rlabel metal2 s 360382 163200 360438 164400 6 la_iena[107]
port 77 nsew signal tristate
rlabel metal2 s 363694 163200 363750 164400 6 la_iena[108]
port 78 nsew signal tristate
rlabel metal2 s 367098 163200 367154 164400 6 la_iena[109]
port 79 nsew signal tristate
rlabel metal2 s 33966 163200 34022 164400 6 la_iena[10]
port 80 nsew signal tristate
rlabel metal2 s 370410 163200 370466 164400 6 la_iena[110]
port 81 nsew signal tristate
rlabel metal2 s 373814 163200 373870 164400 6 la_iena[111]
port 82 nsew signal tristate
rlabel metal2 s 377218 163200 377274 164400 6 la_iena[112]
port 83 nsew signal tristate
rlabel metal2 s 380530 163200 380586 164400 6 la_iena[113]
port 84 nsew signal tristate
rlabel metal2 s 383934 163200 383990 164400 6 la_iena[114]
port 85 nsew signal tristate
rlabel metal2 s 387246 163200 387302 164400 6 la_iena[115]
port 86 nsew signal tristate
rlabel metal2 s 390650 163200 390706 164400 6 la_iena[116]
port 87 nsew signal tristate
rlabel metal2 s 393962 163200 394018 164400 6 la_iena[117]
port 88 nsew signal tristate
rlabel metal2 s 397366 163200 397422 164400 6 la_iena[118]
port 89 nsew signal tristate
rlabel metal2 s 400770 163200 400826 164400 6 la_iena[119]
port 90 nsew signal tristate
rlabel metal2 s 37370 163200 37426 164400 6 la_iena[11]
port 91 nsew signal tristate
rlabel metal2 s 404082 163200 404138 164400 6 la_iena[120]
port 92 nsew signal tristate
rlabel metal2 s 407486 163200 407542 164400 6 la_iena[121]
port 93 nsew signal tristate
rlabel metal2 s 410798 163200 410854 164400 6 la_iena[122]
port 94 nsew signal tristate
rlabel metal2 s 414202 163200 414258 164400 6 la_iena[123]
port 95 nsew signal tristate
rlabel metal2 s 417514 163200 417570 164400 6 la_iena[124]
port 96 nsew signal tristate
rlabel metal2 s 420918 163200 420974 164400 6 la_iena[125]
port 97 nsew signal tristate
rlabel metal2 s 424322 163200 424378 164400 6 la_iena[126]
port 98 nsew signal tristate
rlabel metal2 s 427634 163200 427690 164400 6 la_iena[127]
port 99 nsew signal tristate
rlabel metal2 s 40682 163200 40738 164400 6 la_iena[12]
port 100 nsew signal tristate
rlabel metal2 s 44086 163200 44142 164400 6 la_iena[13]
port 101 nsew signal tristate
rlabel metal2 s 47490 163200 47546 164400 6 la_iena[14]
port 102 nsew signal tristate
rlabel metal2 s 50802 163200 50858 164400 6 la_iena[15]
port 103 nsew signal tristate
rlabel metal2 s 54206 163200 54262 164400 6 la_iena[16]
port 104 nsew signal tristate
rlabel metal2 s 57518 163200 57574 164400 6 la_iena[17]
port 105 nsew signal tristate
rlabel metal2 s 60922 163200 60978 164400 6 la_iena[18]
port 106 nsew signal tristate
rlabel metal2 s 64234 163200 64290 164400 6 la_iena[19]
port 107 nsew signal tristate
rlabel metal2 s 3698 163200 3754 164400 6 la_iena[1]
port 108 nsew signal tristate
rlabel metal2 s 67638 163200 67694 164400 6 la_iena[20]
port 109 nsew signal tristate
rlabel metal2 s 71042 163200 71098 164400 6 la_iena[21]
port 110 nsew signal tristate
rlabel metal2 s 74354 163200 74410 164400 6 la_iena[22]
port 111 nsew signal tristate
rlabel metal2 s 77758 163200 77814 164400 6 la_iena[23]
port 112 nsew signal tristate
rlabel metal2 s 81070 163200 81126 164400 6 la_iena[24]
port 113 nsew signal tristate
rlabel metal2 s 84474 163200 84530 164400 6 la_iena[25]
port 114 nsew signal tristate
rlabel metal2 s 87786 163200 87842 164400 6 la_iena[26]
port 115 nsew signal tristate
rlabel metal2 s 91190 163200 91246 164400 6 la_iena[27]
port 116 nsew signal tristate
rlabel metal2 s 94594 163200 94650 164400 6 la_iena[28]
port 117 nsew signal tristate
rlabel metal2 s 97906 163200 97962 164400 6 la_iena[29]
port 118 nsew signal tristate
rlabel metal2 s 7102 163200 7158 164400 6 la_iena[2]
port 119 nsew signal tristate
rlabel metal2 s 101310 163200 101366 164400 6 la_iena[30]
port 120 nsew signal tristate
rlabel metal2 s 104622 163200 104678 164400 6 la_iena[31]
port 121 nsew signal tristate
rlabel metal2 s 108026 163200 108082 164400 6 la_iena[32]
port 122 nsew signal tristate
rlabel metal2 s 111338 163200 111394 164400 6 la_iena[33]
port 123 nsew signal tristate
rlabel metal2 s 114742 163200 114798 164400 6 la_iena[34]
port 124 nsew signal tristate
rlabel metal2 s 118146 163200 118202 164400 6 la_iena[35]
port 125 nsew signal tristate
rlabel metal2 s 121458 163200 121514 164400 6 la_iena[36]
port 126 nsew signal tristate
rlabel metal2 s 124862 163200 124918 164400 6 la_iena[37]
port 127 nsew signal tristate
rlabel metal2 s 128174 163200 128230 164400 6 la_iena[38]
port 128 nsew signal tristate
rlabel metal2 s 131578 163200 131634 164400 6 la_iena[39]
port 129 nsew signal tristate
rlabel metal2 s 10414 163200 10470 164400 6 la_iena[3]
port 130 nsew signal tristate
rlabel metal2 s 134890 163200 134946 164400 6 la_iena[40]
port 131 nsew signal tristate
rlabel metal2 s 138294 163200 138350 164400 6 la_iena[41]
port 132 nsew signal tristate
rlabel metal2 s 141698 163200 141754 164400 6 la_iena[42]
port 133 nsew signal tristate
rlabel metal2 s 145010 163200 145066 164400 6 la_iena[43]
port 134 nsew signal tristate
rlabel metal2 s 148414 163200 148470 164400 6 la_iena[44]
port 135 nsew signal tristate
rlabel metal2 s 151726 163200 151782 164400 6 la_iena[45]
port 136 nsew signal tristate
rlabel metal2 s 155130 163200 155186 164400 6 la_iena[46]
port 137 nsew signal tristate
rlabel metal2 s 158442 163200 158498 164400 6 la_iena[47]
port 138 nsew signal tristate
rlabel metal2 s 161846 163200 161902 164400 6 la_iena[48]
port 139 nsew signal tristate
rlabel metal2 s 165250 163200 165306 164400 6 la_iena[49]
port 140 nsew signal tristate
rlabel metal2 s 13818 163200 13874 164400 6 la_iena[4]
port 141 nsew signal tristate
rlabel metal2 s 168562 163200 168618 164400 6 la_iena[50]
port 142 nsew signal tristate
rlabel metal2 s 171966 163200 172022 164400 6 la_iena[51]
port 143 nsew signal tristate
rlabel metal2 s 175278 163200 175334 164400 6 la_iena[52]
port 144 nsew signal tristate
rlabel metal2 s 178682 163200 178738 164400 6 la_iena[53]
port 145 nsew signal tristate
rlabel metal2 s 181994 163200 182050 164400 6 la_iena[54]
port 146 nsew signal tristate
rlabel metal2 s 185398 163200 185454 164400 6 la_iena[55]
port 147 nsew signal tristate
rlabel metal2 s 188802 163200 188858 164400 6 la_iena[56]
port 148 nsew signal tristate
rlabel metal2 s 192114 163200 192170 164400 6 la_iena[57]
port 149 nsew signal tristate
rlabel metal2 s 195518 163200 195574 164400 6 la_iena[58]
port 150 nsew signal tristate
rlabel metal2 s 198830 163200 198886 164400 6 la_iena[59]
port 151 nsew signal tristate
rlabel metal2 s 17130 163200 17186 164400 6 la_iena[5]
port 152 nsew signal tristate
rlabel metal2 s 202234 163200 202290 164400 6 la_iena[60]
port 153 nsew signal tristate
rlabel metal2 s 205546 163200 205602 164400 6 la_iena[61]
port 154 nsew signal tristate
rlabel metal2 s 208950 163200 209006 164400 6 la_iena[62]
port 155 nsew signal tristate
rlabel metal2 s 212354 163200 212410 164400 6 la_iena[63]
port 156 nsew signal tristate
rlabel metal2 s 215666 163200 215722 164400 6 la_iena[64]
port 157 nsew signal tristate
rlabel metal2 s 219070 163200 219126 164400 6 la_iena[65]
port 158 nsew signal tristate
rlabel metal2 s 222382 163200 222438 164400 6 la_iena[66]
port 159 nsew signal tristate
rlabel metal2 s 225786 163200 225842 164400 6 la_iena[67]
port 160 nsew signal tristate
rlabel metal2 s 229098 163200 229154 164400 6 la_iena[68]
port 161 nsew signal tristate
rlabel metal2 s 232502 163200 232558 164400 6 la_iena[69]
port 162 nsew signal tristate
rlabel metal2 s 20534 163200 20590 164400 6 la_iena[6]
port 163 nsew signal tristate
rlabel metal2 s 235906 163200 235962 164400 6 la_iena[70]
port 164 nsew signal tristate
rlabel metal2 s 239218 163200 239274 164400 6 la_iena[71]
port 165 nsew signal tristate
rlabel metal2 s 242622 163200 242678 164400 6 la_iena[72]
port 166 nsew signal tristate
rlabel metal2 s 245934 163200 245990 164400 6 la_iena[73]
port 167 nsew signal tristate
rlabel metal2 s 249338 163200 249394 164400 6 la_iena[74]
port 168 nsew signal tristate
rlabel metal2 s 252650 163200 252706 164400 6 la_iena[75]
port 169 nsew signal tristate
rlabel metal2 s 256054 163200 256110 164400 6 la_iena[76]
port 170 nsew signal tristate
rlabel metal2 s 259458 163200 259514 164400 6 la_iena[77]
port 171 nsew signal tristate
rlabel metal2 s 262770 163200 262826 164400 6 la_iena[78]
port 172 nsew signal tristate
rlabel metal2 s 266174 163200 266230 164400 6 la_iena[79]
port 173 nsew signal tristate
rlabel metal2 s 23938 163200 23994 164400 6 la_iena[7]
port 174 nsew signal tristate
rlabel metal2 s 269486 163200 269542 164400 6 la_iena[80]
port 175 nsew signal tristate
rlabel metal2 s 272890 163200 272946 164400 6 la_iena[81]
port 176 nsew signal tristate
rlabel metal2 s 276202 163200 276258 164400 6 la_iena[82]
port 177 nsew signal tristate
rlabel metal2 s 279606 163200 279662 164400 6 la_iena[83]
port 178 nsew signal tristate
rlabel metal2 s 283010 163200 283066 164400 6 la_iena[84]
port 179 nsew signal tristate
rlabel metal2 s 286322 163200 286378 164400 6 la_iena[85]
port 180 nsew signal tristate
rlabel metal2 s 289726 163200 289782 164400 6 la_iena[86]
port 181 nsew signal tristate
rlabel metal2 s 293038 163200 293094 164400 6 la_iena[87]
port 182 nsew signal tristate
rlabel metal2 s 296442 163200 296498 164400 6 la_iena[88]
port 183 nsew signal tristate
rlabel metal2 s 299754 163200 299810 164400 6 la_iena[89]
port 184 nsew signal tristate
rlabel metal2 s 27250 163200 27306 164400 6 la_iena[8]
port 185 nsew signal tristate
rlabel metal2 s 303158 163200 303214 164400 6 la_iena[90]
port 186 nsew signal tristate
rlabel metal2 s 306562 163200 306618 164400 6 la_iena[91]
port 187 nsew signal tristate
rlabel metal2 s 309874 163200 309930 164400 6 la_iena[92]
port 188 nsew signal tristate
rlabel metal2 s 313278 163200 313334 164400 6 la_iena[93]
port 189 nsew signal tristate
rlabel metal2 s 316590 163200 316646 164400 6 la_iena[94]
port 190 nsew signal tristate
rlabel metal2 s 319994 163200 320050 164400 6 la_iena[95]
port 191 nsew signal tristate
rlabel metal2 s 323306 163200 323362 164400 6 la_iena[96]
port 192 nsew signal tristate
rlabel metal2 s 326710 163200 326766 164400 6 la_iena[97]
port 193 nsew signal tristate
rlabel metal2 s 330114 163200 330170 164400 6 la_iena[98]
port 194 nsew signal tristate
rlabel metal2 s 333426 163200 333482 164400 6 la_iena[99]
port 195 nsew signal tristate
rlabel metal2 s 30654 163200 30710 164400 6 la_iena[9]
port 196 nsew signal tristate
rlabel metal2 s 1214 163200 1270 164400 6 la_input[0]
port 197 nsew signal input
rlabel metal2 s 337658 163200 337714 164400 6 la_input[100]
port 198 nsew signal input
rlabel metal2 s 340970 163200 341026 164400 6 la_input[101]
port 199 nsew signal input
rlabel metal2 s 344374 163200 344430 164400 6 la_input[102]
port 200 nsew signal input
rlabel metal2 s 347778 163200 347834 164400 6 la_input[103]
port 201 nsew signal input
rlabel metal2 s 351090 163200 351146 164400 6 la_input[104]
port 202 nsew signal input
rlabel metal2 s 354494 163200 354550 164400 6 la_input[105]
port 203 nsew signal input
rlabel metal2 s 357806 163200 357862 164400 6 la_input[106]
port 204 nsew signal input
rlabel metal2 s 361210 163200 361266 164400 6 la_input[107]
port 205 nsew signal input
rlabel metal2 s 364522 163200 364578 164400 6 la_input[108]
port 206 nsew signal input
rlabel metal2 s 367926 163200 367982 164400 6 la_input[109]
port 207 nsew signal input
rlabel metal2 s 34794 163200 34850 164400 6 la_input[10]
port 208 nsew signal input
rlabel metal2 s 371330 163200 371386 164400 6 la_input[110]
port 209 nsew signal input
rlabel metal2 s 374642 163200 374698 164400 6 la_input[111]
port 210 nsew signal input
rlabel metal2 s 378046 163200 378102 164400 6 la_input[112]
port 211 nsew signal input
rlabel metal2 s 381358 163200 381414 164400 6 la_input[113]
port 212 nsew signal input
rlabel metal2 s 384762 163200 384818 164400 6 la_input[114]
port 213 nsew signal input
rlabel metal2 s 388074 163200 388130 164400 6 la_input[115]
port 214 nsew signal input
rlabel metal2 s 391478 163200 391534 164400 6 la_input[116]
port 215 nsew signal input
rlabel metal2 s 394882 163200 394938 164400 6 la_input[117]
port 216 nsew signal input
rlabel metal2 s 398194 163200 398250 164400 6 la_input[118]
port 217 nsew signal input
rlabel metal2 s 401598 163200 401654 164400 6 la_input[119]
port 218 nsew signal input
rlabel metal2 s 38198 163200 38254 164400 6 la_input[11]
port 219 nsew signal input
rlabel metal2 s 404910 163200 404966 164400 6 la_input[120]
port 220 nsew signal input
rlabel metal2 s 408314 163200 408370 164400 6 la_input[121]
port 221 nsew signal input
rlabel metal2 s 411626 163200 411682 164400 6 la_input[122]
port 222 nsew signal input
rlabel metal2 s 415030 163200 415086 164400 6 la_input[123]
port 223 nsew signal input
rlabel metal2 s 418434 163200 418490 164400 6 la_input[124]
port 224 nsew signal input
rlabel metal2 s 421746 163200 421802 164400 6 la_input[125]
port 225 nsew signal input
rlabel metal2 s 425150 163200 425206 164400 6 la_input[126]
port 226 nsew signal input
rlabel metal2 s 428462 163200 428518 164400 6 la_input[127]
port 227 nsew signal input
rlabel metal2 s 41602 163200 41658 164400 6 la_input[12]
port 228 nsew signal input
rlabel metal2 s 44914 163200 44970 164400 6 la_input[13]
port 229 nsew signal input
rlabel metal2 s 48318 163200 48374 164400 6 la_input[14]
port 230 nsew signal input
rlabel metal2 s 51630 163200 51686 164400 6 la_input[15]
port 231 nsew signal input
rlabel metal2 s 55034 163200 55090 164400 6 la_input[16]
port 232 nsew signal input
rlabel metal2 s 58346 163200 58402 164400 6 la_input[17]
port 233 nsew signal input
rlabel metal2 s 61750 163200 61806 164400 6 la_input[18]
port 234 nsew signal input
rlabel metal2 s 65154 163200 65210 164400 6 la_input[19]
port 235 nsew signal input
rlabel metal2 s 4526 163200 4582 164400 6 la_input[1]
port 236 nsew signal input
rlabel metal2 s 68466 163200 68522 164400 6 la_input[20]
port 237 nsew signal input
rlabel metal2 s 71870 163200 71926 164400 6 la_input[21]
port 238 nsew signal input
rlabel metal2 s 75182 163200 75238 164400 6 la_input[22]
port 239 nsew signal input
rlabel metal2 s 78586 163200 78642 164400 6 la_input[23]
port 240 nsew signal input
rlabel metal2 s 81898 163200 81954 164400 6 la_input[24]
port 241 nsew signal input
rlabel metal2 s 85302 163200 85358 164400 6 la_input[25]
port 242 nsew signal input
rlabel metal2 s 88706 163200 88762 164400 6 la_input[26]
port 243 nsew signal input
rlabel metal2 s 92018 163200 92074 164400 6 la_input[27]
port 244 nsew signal input
rlabel metal2 s 95422 163200 95478 164400 6 la_input[28]
port 245 nsew signal input
rlabel metal2 s 98734 163200 98790 164400 6 la_input[29]
port 246 nsew signal input
rlabel metal2 s 7930 163200 7986 164400 6 la_input[2]
port 247 nsew signal input
rlabel metal2 s 102138 163200 102194 164400 6 la_input[30]
port 248 nsew signal input
rlabel metal2 s 105450 163200 105506 164400 6 la_input[31]
port 249 nsew signal input
rlabel metal2 s 108854 163200 108910 164400 6 la_input[32]
port 250 nsew signal input
rlabel metal2 s 112258 163200 112314 164400 6 la_input[33]
port 251 nsew signal input
rlabel metal2 s 115570 163200 115626 164400 6 la_input[34]
port 252 nsew signal input
rlabel metal2 s 118974 163200 119030 164400 6 la_input[35]
port 253 nsew signal input
rlabel metal2 s 122286 163200 122342 164400 6 la_input[36]
port 254 nsew signal input
rlabel metal2 s 125690 163200 125746 164400 6 la_input[37]
port 255 nsew signal input
rlabel metal2 s 129002 163200 129058 164400 6 la_input[38]
port 256 nsew signal input
rlabel metal2 s 132406 163200 132462 164400 6 la_input[39]
port 257 nsew signal input
rlabel metal2 s 11242 163200 11298 164400 6 la_input[3]
port 258 nsew signal input
rlabel metal2 s 135810 163200 135866 164400 6 la_input[40]
port 259 nsew signal input
rlabel metal2 s 139122 163200 139178 164400 6 la_input[41]
port 260 nsew signal input
rlabel metal2 s 142526 163200 142582 164400 6 la_input[42]
port 261 nsew signal input
rlabel metal2 s 145838 163200 145894 164400 6 la_input[43]
port 262 nsew signal input
rlabel metal2 s 149242 163200 149298 164400 6 la_input[44]
port 263 nsew signal input
rlabel metal2 s 152554 163200 152610 164400 6 la_input[45]
port 264 nsew signal input
rlabel metal2 s 155958 163200 156014 164400 6 la_input[46]
port 265 nsew signal input
rlabel metal2 s 159362 163200 159418 164400 6 la_input[47]
port 266 nsew signal input
rlabel metal2 s 162674 163200 162730 164400 6 la_input[48]
port 267 nsew signal input
rlabel metal2 s 166078 163200 166134 164400 6 la_input[49]
port 268 nsew signal input
rlabel metal2 s 14646 163200 14702 164400 6 la_input[4]
port 269 nsew signal input
rlabel metal2 s 169390 163200 169446 164400 6 la_input[50]
port 270 nsew signal input
rlabel metal2 s 172794 163200 172850 164400 6 la_input[51]
port 271 nsew signal input
rlabel metal2 s 176106 163200 176162 164400 6 la_input[52]
port 272 nsew signal input
rlabel metal2 s 179510 163200 179566 164400 6 la_input[53]
port 273 nsew signal input
rlabel metal2 s 182914 163200 182970 164400 6 la_input[54]
port 274 nsew signal input
rlabel metal2 s 186226 163200 186282 164400 6 la_input[55]
port 275 nsew signal input
rlabel metal2 s 189630 163200 189686 164400 6 la_input[56]
port 276 nsew signal input
rlabel metal2 s 192942 163200 192998 164400 6 la_input[57]
port 277 nsew signal input
rlabel metal2 s 196346 163200 196402 164400 6 la_input[58]
port 278 nsew signal input
rlabel metal2 s 199658 163200 199714 164400 6 la_input[59]
port 279 nsew signal input
rlabel metal2 s 18050 163200 18106 164400 6 la_input[5]
port 280 nsew signal input
rlabel metal2 s 203062 163200 203118 164400 6 la_input[60]
port 281 nsew signal input
rlabel metal2 s 206466 163200 206522 164400 6 la_input[61]
port 282 nsew signal input
rlabel metal2 s 209778 163200 209834 164400 6 la_input[62]
port 283 nsew signal input
rlabel metal2 s 213182 163200 213238 164400 6 la_input[63]
port 284 nsew signal input
rlabel metal2 s 216494 163200 216550 164400 6 la_input[64]
port 285 nsew signal input
rlabel metal2 s 219898 163200 219954 164400 6 la_input[65]
port 286 nsew signal input
rlabel metal2 s 223210 163200 223266 164400 6 la_input[66]
port 287 nsew signal input
rlabel metal2 s 226614 163200 226670 164400 6 la_input[67]
port 288 nsew signal input
rlabel metal2 s 230018 163200 230074 164400 6 la_input[68]
port 289 nsew signal input
rlabel metal2 s 233330 163200 233386 164400 6 la_input[69]
port 290 nsew signal input
rlabel metal2 s 21362 163200 21418 164400 6 la_input[6]
port 291 nsew signal input
rlabel metal2 s 236734 163200 236790 164400 6 la_input[70]
port 292 nsew signal input
rlabel metal2 s 240046 163200 240102 164400 6 la_input[71]
port 293 nsew signal input
rlabel metal2 s 243450 163200 243506 164400 6 la_input[72]
port 294 nsew signal input
rlabel metal2 s 246762 163200 246818 164400 6 la_input[73]
port 295 nsew signal input
rlabel metal2 s 250166 163200 250222 164400 6 la_input[74]
port 296 nsew signal input
rlabel metal2 s 253570 163200 253626 164400 6 la_input[75]
port 297 nsew signal input
rlabel metal2 s 256882 163200 256938 164400 6 la_input[76]
port 298 nsew signal input
rlabel metal2 s 260286 163200 260342 164400 6 la_input[77]
port 299 nsew signal input
rlabel metal2 s 263598 163200 263654 164400 6 la_input[78]
port 300 nsew signal input
rlabel metal2 s 267002 163200 267058 164400 6 la_input[79]
port 301 nsew signal input
rlabel metal2 s 24766 163200 24822 164400 6 la_input[7]
port 302 nsew signal input
rlabel metal2 s 270314 163200 270370 164400 6 la_input[80]
port 303 nsew signal input
rlabel metal2 s 273718 163200 273774 164400 6 la_input[81]
port 304 nsew signal input
rlabel metal2 s 277122 163200 277178 164400 6 la_input[82]
port 305 nsew signal input
rlabel metal2 s 280434 163200 280490 164400 6 la_input[83]
port 306 nsew signal input
rlabel metal2 s 283838 163200 283894 164400 6 la_input[84]
port 307 nsew signal input
rlabel metal2 s 287150 163200 287206 164400 6 la_input[85]
port 308 nsew signal input
rlabel metal2 s 290554 163200 290610 164400 6 la_input[86]
port 309 nsew signal input
rlabel metal2 s 293866 163200 293922 164400 6 la_input[87]
port 310 nsew signal input
rlabel metal2 s 297270 163200 297326 164400 6 la_input[88]
port 311 nsew signal input
rlabel metal2 s 300674 163200 300730 164400 6 la_input[89]
port 312 nsew signal input
rlabel metal2 s 28078 163200 28134 164400 6 la_input[8]
port 313 nsew signal input
rlabel metal2 s 303986 163200 304042 164400 6 la_input[90]
port 314 nsew signal input
rlabel metal2 s 307390 163200 307446 164400 6 la_input[91]
port 315 nsew signal input
rlabel metal2 s 310702 163200 310758 164400 6 la_input[92]
port 316 nsew signal input
rlabel metal2 s 314106 163200 314162 164400 6 la_input[93]
port 317 nsew signal input
rlabel metal2 s 317418 163200 317474 164400 6 la_input[94]
port 318 nsew signal input
rlabel metal2 s 320822 163200 320878 164400 6 la_input[95]
port 319 nsew signal input
rlabel metal2 s 324226 163200 324282 164400 6 la_input[96]
port 320 nsew signal input
rlabel metal2 s 327538 163200 327594 164400 6 la_input[97]
port 321 nsew signal input
rlabel metal2 s 330942 163200 330998 164400 6 la_input[98]
port 322 nsew signal input
rlabel metal2 s 334254 163200 334310 164400 6 la_input[99]
port 323 nsew signal input
rlabel metal2 s 31482 163200 31538 164400 6 la_input[9]
port 324 nsew signal input
rlabel metal2 s 2042 163200 2098 164400 6 la_oenb[0]
port 325 nsew signal tristate
rlabel metal2 s 338486 163200 338542 164400 6 la_oenb[100]
port 326 nsew signal tristate
rlabel metal2 s 341890 163200 341946 164400 6 la_oenb[101]
port 327 nsew signal tristate
rlabel metal2 s 345202 163200 345258 164400 6 la_oenb[102]
port 328 nsew signal tristate
rlabel metal2 s 348606 163200 348662 164400 6 la_oenb[103]
port 329 nsew signal tristate
rlabel metal2 s 351918 163200 351974 164400 6 la_oenb[104]
port 330 nsew signal tristate
rlabel metal2 s 355322 163200 355378 164400 6 la_oenb[105]
port 331 nsew signal tristate
rlabel metal2 s 358634 163200 358690 164400 6 la_oenb[106]
port 332 nsew signal tristate
rlabel metal2 s 362038 163200 362094 164400 6 la_oenb[107]
port 333 nsew signal tristate
rlabel metal2 s 365442 163200 365498 164400 6 la_oenb[108]
port 334 nsew signal tristate
rlabel metal2 s 368754 163200 368810 164400 6 la_oenb[109]
port 335 nsew signal tristate
rlabel metal2 s 35714 163200 35770 164400 6 la_oenb[10]
port 336 nsew signal tristate
rlabel metal2 s 372158 163200 372214 164400 6 la_oenb[110]
port 337 nsew signal tristate
rlabel metal2 s 375470 163200 375526 164400 6 la_oenb[111]
port 338 nsew signal tristate
rlabel metal2 s 378874 163200 378930 164400 6 la_oenb[112]
port 339 nsew signal tristate
rlabel metal2 s 382186 163200 382242 164400 6 la_oenb[113]
port 340 nsew signal tristate
rlabel metal2 s 385590 163200 385646 164400 6 la_oenb[114]
port 341 nsew signal tristate
rlabel metal2 s 388994 163200 389050 164400 6 la_oenb[115]
port 342 nsew signal tristate
rlabel metal2 s 392306 163200 392362 164400 6 la_oenb[116]
port 343 nsew signal tristate
rlabel metal2 s 395710 163200 395766 164400 6 la_oenb[117]
port 344 nsew signal tristate
rlabel metal2 s 399022 163200 399078 164400 6 la_oenb[118]
port 345 nsew signal tristate
rlabel metal2 s 402426 163200 402482 164400 6 la_oenb[119]
port 346 nsew signal tristate
rlabel metal2 s 39026 163200 39082 164400 6 la_oenb[11]
port 347 nsew signal tristate
rlabel metal2 s 405738 163200 405794 164400 6 la_oenb[120]
port 348 nsew signal tristate
rlabel metal2 s 409142 163200 409198 164400 6 la_oenb[121]
port 349 nsew signal tristate
rlabel metal2 s 412546 163200 412602 164400 6 la_oenb[122]
port 350 nsew signal tristate
rlabel metal2 s 415858 163200 415914 164400 6 la_oenb[123]
port 351 nsew signal tristate
rlabel metal2 s 419262 163200 419318 164400 6 la_oenb[124]
port 352 nsew signal tristate
rlabel metal2 s 422574 163200 422630 164400 6 la_oenb[125]
port 353 nsew signal tristate
rlabel metal2 s 425978 163200 426034 164400 6 la_oenb[126]
port 354 nsew signal tristate
rlabel metal2 s 429290 163200 429346 164400 6 la_oenb[127]
port 355 nsew signal tristate
rlabel metal2 s 42430 163200 42486 164400 6 la_oenb[12]
port 356 nsew signal tristate
rlabel metal2 s 45742 163200 45798 164400 6 la_oenb[13]
port 357 nsew signal tristate
rlabel metal2 s 49146 163200 49202 164400 6 la_oenb[14]
port 358 nsew signal tristate
rlabel metal2 s 52458 163200 52514 164400 6 la_oenb[15]
port 359 nsew signal tristate
rlabel metal2 s 55862 163200 55918 164400 6 la_oenb[16]
port 360 nsew signal tristate
rlabel metal2 s 59266 163200 59322 164400 6 la_oenb[17]
port 361 nsew signal tristate
rlabel metal2 s 62578 163200 62634 164400 6 la_oenb[18]
port 362 nsew signal tristate
rlabel metal2 s 65982 163200 66038 164400 6 la_oenb[19]
port 363 nsew signal tristate
rlabel metal2 s 5354 163200 5410 164400 6 la_oenb[1]
port 364 nsew signal tristate
rlabel metal2 s 69294 163200 69350 164400 6 la_oenb[20]
port 365 nsew signal tristate
rlabel metal2 s 72698 163200 72754 164400 6 la_oenb[21]
port 366 nsew signal tristate
rlabel metal2 s 76010 163200 76066 164400 6 la_oenb[22]
port 367 nsew signal tristate
rlabel metal2 s 79414 163200 79470 164400 6 la_oenb[23]
port 368 nsew signal tristate
rlabel metal2 s 82818 163200 82874 164400 6 la_oenb[24]
port 369 nsew signal tristate
rlabel metal2 s 86130 163200 86186 164400 6 la_oenb[25]
port 370 nsew signal tristate
rlabel metal2 s 89534 163200 89590 164400 6 la_oenb[26]
port 371 nsew signal tristate
rlabel metal2 s 92846 163200 92902 164400 6 la_oenb[27]
port 372 nsew signal tristate
rlabel metal2 s 96250 163200 96306 164400 6 la_oenb[28]
port 373 nsew signal tristate
rlabel metal2 s 99562 163200 99618 164400 6 la_oenb[29]
port 374 nsew signal tristate
rlabel metal2 s 8758 163200 8814 164400 6 la_oenb[2]
port 375 nsew signal tristate
rlabel metal2 s 102966 163200 103022 164400 6 la_oenb[30]
port 376 nsew signal tristate
rlabel metal2 s 106370 163200 106426 164400 6 la_oenb[31]
port 377 nsew signal tristate
rlabel metal2 s 109682 163200 109738 164400 6 la_oenb[32]
port 378 nsew signal tristate
rlabel metal2 s 113086 163200 113142 164400 6 la_oenb[33]
port 379 nsew signal tristate
rlabel metal2 s 116398 163200 116454 164400 6 la_oenb[34]
port 380 nsew signal tristate
rlabel metal2 s 119802 163200 119858 164400 6 la_oenb[35]
port 381 nsew signal tristate
rlabel metal2 s 123114 163200 123170 164400 6 la_oenb[36]
port 382 nsew signal tristate
rlabel metal2 s 126518 163200 126574 164400 6 la_oenb[37]
port 383 nsew signal tristate
rlabel metal2 s 129922 163200 129978 164400 6 la_oenb[38]
port 384 nsew signal tristate
rlabel metal2 s 133234 163200 133290 164400 6 la_oenb[39]
port 385 nsew signal tristate
rlabel metal2 s 12162 163200 12218 164400 6 la_oenb[3]
port 386 nsew signal tristate
rlabel metal2 s 136638 163200 136694 164400 6 la_oenb[40]
port 387 nsew signal tristate
rlabel metal2 s 139950 163200 140006 164400 6 la_oenb[41]
port 388 nsew signal tristate
rlabel metal2 s 143354 163200 143410 164400 6 la_oenb[42]
port 389 nsew signal tristate
rlabel metal2 s 146666 163200 146722 164400 6 la_oenb[43]
port 390 nsew signal tristate
rlabel metal2 s 150070 163200 150126 164400 6 la_oenb[44]
port 391 nsew signal tristate
rlabel metal2 s 153474 163200 153530 164400 6 la_oenb[45]
port 392 nsew signal tristate
rlabel metal2 s 156786 163200 156842 164400 6 la_oenb[46]
port 393 nsew signal tristate
rlabel metal2 s 160190 163200 160246 164400 6 la_oenb[47]
port 394 nsew signal tristate
rlabel metal2 s 163502 163200 163558 164400 6 la_oenb[48]
port 395 nsew signal tristate
rlabel metal2 s 166906 163200 166962 164400 6 la_oenb[49]
port 396 nsew signal tristate
rlabel metal2 s 15474 163200 15530 164400 6 la_oenb[4]
port 397 nsew signal tristate
rlabel metal2 s 170218 163200 170274 164400 6 la_oenb[50]
port 398 nsew signal tristate
rlabel metal2 s 173622 163200 173678 164400 6 la_oenb[51]
port 399 nsew signal tristate
rlabel metal2 s 177026 163200 177082 164400 6 la_oenb[52]
port 400 nsew signal tristate
rlabel metal2 s 180338 163200 180394 164400 6 la_oenb[53]
port 401 nsew signal tristate
rlabel metal2 s 183742 163200 183798 164400 6 la_oenb[54]
port 402 nsew signal tristate
rlabel metal2 s 187054 163200 187110 164400 6 la_oenb[55]
port 403 nsew signal tristate
rlabel metal2 s 190458 163200 190514 164400 6 la_oenb[56]
port 404 nsew signal tristate
rlabel metal2 s 193770 163200 193826 164400 6 la_oenb[57]
port 405 nsew signal tristate
rlabel metal2 s 197174 163200 197230 164400 6 la_oenb[58]
port 406 nsew signal tristate
rlabel metal2 s 200578 163200 200634 164400 6 la_oenb[59]
port 407 nsew signal tristate
rlabel metal2 s 18878 163200 18934 164400 6 la_oenb[5]
port 408 nsew signal tristate
rlabel metal2 s 203890 163200 203946 164400 6 la_oenb[60]
port 409 nsew signal tristate
rlabel metal2 s 207294 163200 207350 164400 6 la_oenb[61]
port 410 nsew signal tristate
rlabel metal2 s 210606 163200 210662 164400 6 la_oenb[62]
port 411 nsew signal tristate
rlabel metal2 s 214010 163200 214066 164400 6 la_oenb[63]
port 412 nsew signal tristate
rlabel metal2 s 217322 163200 217378 164400 6 la_oenb[64]
port 413 nsew signal tristate
rlabel metal2 s 220726 163200 220782 164400 6 la_oenb[65]
port 414 nsew signal tristate
rlabel metal2 s 224130 163200 224186 164400 6 la_oenb[66]
port 415 nsew signal tristate
rlabel metal2 s 227442 163200 227498 164400 6 la_oenb[67]
port 416 nsew signal tristate
rlabel metal2 s 230846 163200 230902 164400 6 la_oenb[68]
port 417 nsew signal tristate
rlabel metal2 s 234158 163200 234214 164400 6 la_oenb[69]
port 418 nsew signal tristate
rlabel metal2 s 22190 163200 22246 164400 6 la_oenb[6]
port 419 nsew signal tristate
rlabel metal2 s 237562 163200 237618 164400 6 la_oenb[70]
port 420 nsew signal tristate
rlabel metal2 s 240874 163200 240930 164400 6 la_oenb[71]
port 421 nsew signal tristate
rlabel metal2 s 244278 163200 244334 164400 6 la_oenb[72]
port 422 nsew signal tristate
rlabel metal2 s 247682 163200 247738 164400 6 la_oenb[73]
port 423 nsew signal tristate
rlabel metal2 s 250994 163200 251050 164400 6 la_oenb[74]
port 424 nsew signal tristate
rlabel metal2 s 254398 163200 254454 164400 6 la_oenb[75]
port 425 nsew signal tristate
rlabel metal2 s 257710 163200 257766 164400 6 la_oenb[76]
port 426 nsew signal tristate
rlabel metal2 s 261114 163200 261170 164400 6 la_oenb[77]
port 427 nsew signal tristate
rlabel metal2 s 264426 163200 264482 164400 6 la_oenb[78]
port 428 nsew signal tristate
rlabel metal2 s 267830 163200 267886 164400 6 la_oenb[79]
port 429 nsew signal tristate
rlabel metal2 s 25594 163200 25650 164400 6 la_oenb[7]
port 430 nsew signal tristate
rlabel metal2 s 271234 163200 271290 164400 6 la_oenb[80]
port 431 nsew signal tristate
rlabel metal2 s 274546 163200 274602 164400 6 la_oenb[81]
port 432 nsew signal tristate
rlabel metal2 s 277950 163200 278006 164400 6 la_oenb[82]
port 433 nsew signal tristate
rlabel metal2 s 281262 163200 281318 164400 6 la_oenb[83]
port 434 nsew signal tristate
rlabel metal2 s 284666 163200 284722 164400 6 la_oenb[84]
port 435 nsew signal tristate
rlabel metal2 s 287978 163200 288034 164400 6 la_oenb[85]
port 436 nsew signal tristate
rlabel metal2 s 291382 163200 291438 164400 6 la_oenb[86]
port 437 nsew signal tristate
rlabel metal2 s 294786 163200 294842 164400 6 la_oenb[87]
port 438 nsew signal tristate
rlabel metal2 s 298098 163200 298154 164400 6 la_oenb[88]
port 439 nsew signal tristate
rlabel metal2 s 301502 163200 301558 164400 6 la_oenb[89]
port 440 nsew signal tristate
rlabel metal2 s 28906 163200 28962 164400 6 la_oenb[8]
port 441 nsew signal tristate
rlabel metal2 s 304814 163200 304870 164400 6 la_oenb[90]
port 442 nsew signal tristate
rlabel metal2 s 308218 163200 308274 164400 6 la_oenb[91]
port 443 nsew signal tristate
rlabel metal2 s 311530 163200 311586 164400 6 la_oenb[92]
port 444 nsew signal tristate
rlabel metal2 s 314934 163200 314990 164400 6 la_oenb[93]
port 445 nsew signal tristate
rlabel metal2 s 318338 163200 318394 164400 6 la_oenb[94]
port 446 nsew signal tristate
rlabel metal2 s 321650 163200 321706 164400 6 la_oenb[95]
port 447 nsew signal tristate
rlabel metal2 s 325054 163200 325110 164400 6 la_oenb[96]
port 448 nsew signal tristate
rlabel metal2 s 328366 163200 328422 164400 6 la_oenb[97]
port 449 nsew signal tristate
rlabel metal2 s 331770 163200 331826 164400 6 la_oenb[98]
port 450 nsew signal tristate
rlabel metal2 s 335082 163200 335138 164400 6 la_oenb[99]
port 451 nsew signal tristate
rlabel metal2 s 32310 163200 32366 164400 6 la_oenb[9]
port 452 nsew signal tristate
rlabel metal2 s 2870 163200 2926 164400 6 la_output[0]
port 453 nsew signal tristate
rlabel metal2 s 339314 163200 339370 164400 6 la_output[100]
port 454 nsew signal tristate
rlabel metal2 s 342718 163200 342774 164400 6 la_output[101]
port 455 nsew signal tristate
rlabel metal2 s 346030 163200 346086 164400 6 la_output[102]
port 456 nsew signal tristate
rlabel metal2 s 349434 163200 349490 164400 6 la_output[103]
port 457 nsew signal tristate
rlabel metal2 s 352746 163200 352802 164400 6 la_output[104]
port 458 nsew signal tristate
rlabel metal2 s 356150 163200 356206 164400 6 la_output[105]
port 459 nsew signal tristate
rlabel metal2 s 359554 163200 359610 164400 6 la_output[106]
port 460 nsew signal tristate
rlabel metal2 s 362866 163200 362922 164400 6 la_output[107]
port 461 nsew signal tristate
rlabel metal2 s 366270 163200 366326 164400 6 la_output[108]
port 462 nsew signal tristate
rlabel metal2 s 369582 163200 369638 164400 6 la_output[109]
port 463 nsew signal tristate
rlabel metal2 s 36542 163200 36598 164400 6 la_output[10]
port 464 nsew signal tristate
rlabel metal2 s 372986 163200 373042 164400 6 la_output[110]
port 465 nsew signal tristate
rlabel metal2 s 376298 163200 376354 164400 6 la_output[111]
port 466 nsew signal tristate
rlabel metal2 s 379702 163200 379758 164400 6 la_output[112]
port 467 nsew signal tristate
rlabel metal2 s 383106 163200 383162 164400 6 la_output[113]
port 468 nsew signal tristate
rlabel metal2 s 386418 163200 386474 164400 6 la_output[114]
port 469 nsew signal tristate
rlabel metal2 s 389822 163200 389878 164400 6 la_output[115]
port 470 nsew signal tristate
rlabel metal2 s 393134 163200 393190 164400 6 la_output[116]
port 471 nsew signal tristate
rlabel metal2 s 396538 163200 396594 164400 6 la_output[117]
port 472 nsew signal tristate
rlabel metal2 s 399850 163200 399906 164400 6 la_output[118]
port 473 nsew signal tristate
rlabel metal2 s 403254 163200 403310 164400 6 la_output[119]
port 474 nsew signal tristate
rlabel metal2 s 39854 163200 39910 164400 6 la_output[11]
port 475 nsew signal tristate
rlabel metal2 s 406658 163200 406714 164400 6 la_output[120]
port 476 nsew signal tristate
rlabel metal2 s 409970 163200 410026 164400 6 la_output[121]
port 477 nsew signal tristate
rlabel metal2 s 413374 163200 413430 164400 6 la_output[122]
port 478 nsew signal tristate
rlabel metal2 s 416686 163200 416742 164400 6 la_output[123]
port 479 nsew signal tristate
rlabel metal2 s 420090 163200 420146 164400 6 la_output[124]
port 480 nsew signal tristate
rlabel metal2 s 423402 163200 423458 164400 6 la_output[125]
port 481 nsew signal tristate
rlabel metal2 s 426806 163200 426862 164400 6 la_output[126]
port 482 nsew signal tristate
rlabel metal2 s 430210 163200 430266 164400 6 la_output[127]
port 483 nsew signal tristate
rlabel metal2 s 43258 163200 43314 164400 6 la_output[12]
port 484 nsew signal tristate
rlabel metal2 s 46570 163200 46626 164400 6 la_output[13]
port 485 nsew signal tristate
rlabel metal2 s 49974 163200 50030 164400 6 la_output[14]
port 486 nsew signal tristate
rlabel metal2 s 53378 163200 53434 164400 6 la_output[15]
port 487 nsew signal tristate
rlabel metal2 s 56690 163200 56746 164400 6 la_output[16]
port 488 nsew signal tristate
rlabel metal2 s 60094 163200 60150 164400 6 la_output[17]
port 489 nsew signal tristate
rlabel metal2 s 63406 163200 63462 164400 6 la_output[18]
port 490 nsew signal tristate
rlabel metal2 s 66810 163200 66866 164400 6 la_output[19]
port 491 nsew signal tristate
rlabel metal2 s 6274 163200 6330 164400 6 la_output[1]
port 492 nsew signal tristate
rlabel metal2 s 70122 163200 70178 164400 6 la_output[20]
port 493 nsew signal tristate
rlabel metal2 s 73526 163200 73582 164400 6 la_output[21]
port 494 nsew signal tristate
rlabel metal2 s 76930 163200 76986 164400 6 la_output[22]
port 495 nsew signal tristate
rlabel metal2 s 80242 163200 80298 164400 6 la_output[23]
port 496 nsew signal tristate
rlabel metal2 s 83646 163200 83702 164400 6 la_output[24]
port 497 nsew signal tristate
rlabel metal2 s 86958 163200 87014 164400 6 la_output[25]
port 498 nsew signal tristate
rlabel metal2 s 90362 163200 90418 164400 6 la_output[26]
port 499 nsew signal tristate
rlabel metal2 s 93674 163200 93730 164400 6 la_output[27]
port 500 nsew signal tristate
rlabel metal2 s 97078 163200 97134 164400 6 la_output[28]
port 501 nsew signal tristate
rlabel metal2 s 100482 163200 100538 164400 6 la_output[29]
port 502 nsew signal tristate
rlabel metal2 s 9586 163200 9642 164400 6 la_output[2]
port 503 nsew signal tristate
rlabel metal2 s 103794 163200 103850 164400 6 la_output[30]
port 504 nsew signal tristate
rlabel metal2 s 107198 163200 107254 164400 6 la_output[31]
port 505 nsew signal tristate
rlabel metal2 s 110510 163200 110566 164400 6 la_output[32]
port 506 nsew signal tristate
rlabel metal2 s 113914 163200 113970 164400 6 la_output[33]
port 507 nsew signal tristate
rlabel metal2 s 117226 163200 117282 164400 6 la_output[34]
port 508 nsew signal tristate
rlabel metal2 s 120630 163200 120686 164400 6 la_output[35]
port 509 nsew signal tristate
rlabel metal2 s 124034 163200 124090 164400 6 la_output[36]
port 510 nsew signal tristate
rlabel metal2 s 127346 163200 127402 164400 6 la_output[37]
port 511 nsew signal tristate
rlabel metal2 s 130750 163200 130806 164400 6 la_output[38]
port 512 nsew signal tristate
rlabel metal2 s 134062 163200 134118 164400 6 la_output[39]
port 513 nsew signal tristate
rlabel metal2 s 12990 163200 13046 164400 6 la_output[3]
port 514 nsew signal tristate
rlabel metal2 s 137466 163200 137522 164400 6 la_output[40]
port 515 nsew signal tristate
rlabel metal2 s 140778 163200 140834 164400 6 la_output[41]
port 516 nsew signal tristate
rlabel metal2 s 144182 163200 144238 164400 6 la_output[42]
port 517 nsew signal tristate
rlabel metal2 s 147586 163200 147642 164400 6 la_output[43]
port 518 nsew signal tristate
rlabel metal2 s 150898 163200 150954 164400 6 la_output[44]
port 519 nsew signal tristate
rlabel metal2 s 154302 163200 154358 164400 6 la_output[45]
port 520 nsew signal tristate
rlabel metal2 s 157614 163200 157670 164400 6 la_output[46]
port 521 nsew signal tristate
rlabel metal2 s 161018 163200 161074 164400 6 la_output[47]
port 522 nsew signal tristate
rlabel metal2 s 164330 163200 164386 164400 6 la_output[48]
port 523 nsew signal tristate
rlabel metal2 s 167734 163200 167790 164400 6 la_output[49]
port 524 nsew signal tristate
rlabel metal2 s 16302 163200 16358 164400 6 la_output[4]
port 525 nsew signal tristate
rlabel metal2 s 171138 163200 171194 164400 6 la_output[50]
port 526 nsew signal tristate
rlabel metal2 s 174450 163200 174506 164400 6 la_output[51]
port 527 nsew signal tristate
rlabel metal2 s 177854 163200 177910 164400 6 la_output[52]
port 528 nsew signal tristate
rlabel metal2 s 181166 163200 181222 164400 6 la_output[53]
port 529 nsew signal tristate
rlabel metal2 s 184570 163200 184626 164400 6 la_output[54]
port 530 nsew signal tristate
rlabel metal2 s 187882 163200 187938 164400 6 la_output[55]
port 531 nsew signal tristate
rlabel metal2 s 191286 163200 191342 164400 6 la_output[56]
port 532 nsew signal tristate
rlabel metal2 s 194690 163200 194746 164400 6 la_output[57]
port 533 nsew signal tristate
rlabel metal2 s 198002 163200 198058 164400 6 la_output[58]
port 534 nsew signal tristate
rlabel metal2 s 201406 163200 201462 164400 6 la_output[59]
port 535 nsew signal tristate
rlabel metal2 s 19706 163200 19762 164400 6 la_output[5]
port 536 nsew signal tristate
rlabel metal2 s 204718 163200 204774 164400 6 la_output[60]
port 537 nsew signal tristate
rlabel metal2 s 208122 163200 208178 164400 6 la_output[61]
port 538 nsew signal tristate
rlabel metal2 s 211434 163200 211490 164400 6 la_output[62]
port 539 nsew signal tristate
rlabel metal2 s 214838 163200 214894 164400 6 la_output[63]
port 540 nsew signal tristate
rlabel metal2 s 218242 163200 218298 164400 6 la_output[64]
port 541 nsew signal tristate
rlabel metal2 s 221554 163200 221610 164400 6 la_output[65]
port 542 nsew signal tristate
rlabel metal2 s 224958 163200 225014 164400 6 la_output[66]
port 543 nsew signal tristate
rlabel metal2 s 228270 163200 228326 164400 6 la_output[67]
port 544 nsew signal tristate
rlabel metal2 s 231674 163200 231730 164400 6 la_output[68]
port 545 nsew signal tristate
rlabel metal2 s 234986 163200 235042 164400 6 la_output[69]
port 546 nsew signal tristate
rlabel metal2 s 23018 163200 23074 164400 6 la_output[6]
port 547 nsew signal tristate
rlabel metal2 s 238390 163200 238446 164400 6 la_output[70]
port 548 nsew signal tristate
rlabel metal2 s 241794 163200 241850 164400 6 la_output[71]
port 549 nsew signal tristate
rlabel metal2 s 245106 163200 245162 164400 6 la_output[72]
port 550 nsew signal tristate
rlabel metal2 s 248510 163200 248566 164400 6 la_output[73]
port 551 nsew signal tristate
rlabel metal2 s 251822 163200 251878 164400 6 la_output[74]
port 552 nsew signal tristate
rlabel metal2 s 255226 163200 255282 164400 6 la_output[75]
port 553 nsew signal tristate
rlabel metal2 s 258538 163200 258594 164400 6 la_output[76]
port 554 nsew signal tristate
rlabel metal2 s 261942 163200 261998 164400 6 la_output[77]
port 555 nsew signal tristate
rlabel metal2 s 265346 163200 265402 164400 6 la_output[78]
port 556 nsew signal tristate
rlabel metal2 s 268658 163200 268714 164400 6 la_output[79]
port 557 nsew signal tristate
rlabel metal2 s 26422 163200 26478 164400 6 la_output[7]
port 558 nsew signal tristate
rlabel metal2 s 272062 163200 272118 164400 6 la_output[80]
port 559 nsew signal tristate
rlabel metal2 s 275374 163200 275430 164400 6 la_output[81]
port 560 nsew signal tristate
rlabel metal2 s 278778 163200 278834 164400 6 la_output[82]
port 561 nsew signal tristate
rlabel metal2 s 282090 163200 282146 164400 6 la_output[83]
port 562 nsew signal tristate
rlabel metal2 s 285494 163200 285550 164400 6 la_output[84]
port 563 nsew signal tristate
rlabel metal2 s 288898 163200 288954 164400 6 la_output[85]
port 564 nsew signal tristate
rlabel metal2 s 292210 163200 292266 164400 6 la_output[86]
port 565 nsew signal tristate
rlabel metal2 s 295614 163200 295670 164400 6 la_output[87]
port 566 nsew signal tristate
rlabel metal2 s 298926 163200 298982 164400 6 la_output[88]
port 567 nsew signal tristate
rlabel metal2 s 302330 163200 302386 164400 6 la_output[89]
port 568 nsew signal tristate
rlabel metal2 s 29826 163200 29882 164400 6 la_output[8]
port 569 nsew signal tristate
rlabel metal2 s 305642 163200 305698 164400 6 la_output[90]
port 570 nsew signal tristate
rlabel metal2 s 309046 163200 309102 164400 6 la_output[91]
port 571 nsew signal tristate
rlabel metal2 s 312450 163200 312506 164400 6 la_output[92]
port 572 nsew signal tristate
rlabel metal2 s 315762 163200 315818 164400 6 la_output[93]
port 573 nsew signal tristate
rlabel metal2 s 319166 163200 319222 164400 6 la_output[94]
port 574 nsew signal tristate
rlabel metal2 s 322478 163200 322534 164400 6 la_output[95]
port 575 nsew signal tristate
rlabel metal2 s 325882 163200 325938 164400 6 la_output[96]
port 576 nsew signal tristate
rlabel metal2 s 329194 163200 329250 164400 6 la_output[97]
port 577 nsew signal tristate
rlabel metal2 s 332598 163200 332654 164400 6 la_output[98]
port 578 nsew signal tristate
rlabel metal2 s 336002 163200 336058 164400 6 la_output[99]
port 579 nsew signal tristate
rlabel metal2 s 33138 163200 33194 164400 6 la_output[9]
port 580 nsew signal tristate
rlabel metal2 s 431038 163200 431094 164400 6 mprj_ack_i
port 581 nsew signal input
rlabel metal2 s 435178 163200 435234 164400 6 mprj_adr_o[0]
port 582 nsew signal tristate
rlabel metal2 s 463790 163200 463846 164400 6 mprj_adr_o[10]
port 583 nsew signal tristate
rlabel metal2 s 466366 163200 466422 164400 6 mprj_adr_o[11]
port 584 nsew signal tristate
rlabel metal2 s 468850 163200 468906 164400 6 mprj_adr_o[12]
port 585 nsew signal tristate
rlabel metal2 s 471426 163200 471482 164400 6 mprj_adr_o[13]
port 586 nsew signal tristate
rlabel metal2 s 473910 163200 473966 164400 6 mprj_adr_o[14]
port 587 nsew signal tristate
rlabel metal2 s 476394 163200 476450 164400 6 mprj_adr_o[15]
port 588 nsew signal tristate
rlabel metal2 s 478970 163200 479026 164400 6 mprj_adr_o[16]
port 589 nsew signal tristate
rlabel metal2 s 481454 163200 481510 164400 6 mprj_adr_o[17]
port 590 nsew signal tristate
rlabel metal2 s 484030 163200 484086 164400 6 mprj_adr_o[18]
port 591 nsew signal tristate
rlabel metal2 s 486514 163200 486570 164400 6 mprj_adr_o[19]
port 592 nsew signal tristate
rlabel metal2 s 438582 163200 438638 164400 6 mprj_adr_o[1]
port 593 nsew signal tristate
rlabel metal2 s 489090 163200 489146 164400 6 mprj_adr_o[20]
port 594 nsew signal tristate
rlabel metal2 s 491574 163200 491630 164400 6 mprj_adr_o[21]
port 595 nsew signal tristate
rlabel metal2 s 494058 163200 494114 164400 6 mprj_adr_o[22]
port 596 nsew signal tristate
rlabel metal2 s 496634 163200 496690 164400 6 mprj_adr_o[23]
port 597 nsew signal tristate
rlabel metal2 s 499118 163200 499174 164400 6 mprj_adr_o[24]
port 598 nsew signal tristate
rlabel metal2 s 501694 163200 501750 164400 6 mprj_adr_o[25]
port 599 nsew signal tristate
rlabel metal2 s 504178 163200 504234 164400 6 mprj_adr_o[26]
port 600 nsew signal tristate
rlabel metal2 s 506754 163200 506810 164400 6 mprj_adr_o[27]
port 601 nsew signal tristate
rlabel metal2 s 509238 163200 509294 164400 6 mprj_adr_o[28]
port 602 nsew signal tristate
rlabel metal2 s 511722 163200 511778 164400 6 mprj_adr_o[29]
port 603 nsew signal tristate
rlabel metal2 s 441986 163200 442042 164400 6 mprj_adr_o[2]
port 604 nsew signal tristate
rlabel metal2 s 514298 163200 514354 164400 6 mprj_adr_o[30]
port 605 nsew signal tristate
rlabel metal2 s 516782 163200 516838 164400 6 mprj_adr_o[31]
port 606 nsew signal tristate
rlabel metal2 s 445298 163200 445354 164400 6 mprj_adr_o[3]
port 607 nsew signal tristate
rlabel metal2 s 448702 163200 448758 164400 6 mprj_adr_o[4]
port 608 nsew signal tristate
rlabel metal2 s 451186 163200 451242 164400 6 mprj_adr_o[5]
port 609 nsew signal tristate
rlabel metal2 s 453762 163200 453818 164400 6 mprj_adr_o[6]
port 610 nsew signal tristate
rlabel metal2 s 456246 163200 456302 164400 6 mprj_adr_o[7]
port 611 nsew signal tristate
rlabel metal2 s 458730 163200 458786 164400 6 mprj_adr_o[8]
port 612 nsew signal tristate
rlabel metal2 s 461306 163200 461362 164400 6 mprj_adr_o[9]
port 613 nsew signal tristate
rlabel metal2 s 431866 163200 431922 164400 6 mprj_cyc_o
port 614 nsew signal tristate
rlabel metal2 s 436098 163200 436154 164400 6 mprj_dat_i[0]
port 615 nsew signal input
rlabel metal2 s 464618 163200 464674 164400 6 mprj_dat_i[10]
port 616 nsew signal input
rlabel metal2 s 467194 163200 467250 164400 6 mprj_dat_i[11]
port 617 nsew signal input
rlabel metal2 s 469678 163200 469734 164400 6 mprj_dat_i[12]
port 618 nsew signal input
rlabel metal2 s 472254 163200 472310 164400 6 mprj_dat_i[13]
port 619 nsew signal input
rlabel metal2 s 474738 163200 474794 164400 6 mprj_dat_i[14]
port 620 nsew signal input
rlabel metal2 s 477314 163200 477370 164400 6 mprj_dat_i[15]
port 621 nsew signal input
rlabel metal2 s 479798 163200 479854 164400 6 mprj_dat_i[16]
port 622 nsew signal input
rlabel metal2 s 482282 163200 482338 164400 6 mprj_dat_i[17]
port 623 nsew signal input
rlabel metal2 s 484858 163200 484914 164400 6 mprj_dat_i[18]
port 624 nsew signal input
rlabel metal2 s 487342 163200 487398 164400 6 mprj_dat_i[19]
port 625 nsew signal input
rlabel metal2 s 439410 163200 439466 164400 6 mprj_dat_i[1]
port 626 nsew signal input
rlabel metal2 s 489918 163200 489974 164400 6 mprj_dat_i[20]
port 627 nsew signal input
rlabel metal2 s 492402 163200 492458 164400 6 mprj_dat_i[21]
port 628 nsew signal input
rlabel metal2 s 494978 163200 495034 164400 6 mprj_dat_i[22]
port 629 nsew signal input
rlabel metal2 s 497462 163200 497518 164400 6 mprj_dat_i[23]
port 630 nsew signal input
rlabel metal2 s 499946 163200 500002 164400 6 mprj_dat_i[24]
port 631 nsew signal input
rlabel metal2 s 502522 163200 502578 164400 6 mprj_dat_i[25]
port 632 nsew signal input
rlabel metal2 s 505006 163200 505062 164400 6 mprj_dat_i[26]
port 633 nsew signal input
rlabel metal2 s 507582 163200 507638 164400 6 mprj_dat_i[27]
port 634 nsew signal input
rlabel metal2 s 510066 163200 510122 164400 6 mprj_dat_i[28]
port 635 nsew signal input
rlabel metal2 s 512642 163200 512698 164400 6 mprj_dat_i[29]
port 636 nsew signal input
rlabel metal2 s 442814 163200 442870 164400 6 mprj_dat_i[2]
port 637 nsew signal input
rlabel metal2 s 515126 163200 515182 164400 6 mprj_dat_i[30]
port 638 nsew signal input
rlabel metal2 s 517610 163200 517666 164400 6 mprj_dat_i[31]
port 639 nsew signal input
rlabel metal2 s 446126 163200 446182 164400 6 mprj_dat_i[3]
port 640 nsew signal input
rlabel metal2 s 449530 163200 449586 164400 6 mprj_dat_i[4]
port 641 nsew signal input
rlabel metal2 s 452014 163200 452070 164400 6 mprj_dat_i[5]
port 642 nsew signal input
rlabel metal2 s 454590 163200 454646 164400 6 mprj_dat_i[6]
port 643 nsew signal input
rlabel metal2 s 457074 163200 457130 164400 6 mprj_dat_i[7]
port 644 nsew signal input
rlabel metal2 s 459650 163200 459706 164400 6 mprj_dat_i[8]
port 645 nsew signal input
rlabel metal2 s 462134 163200 462190 164400 6 mprj_dat_i[9]
port 646 nsew signal input
rlabel metal2 s 436926 163200 436982 164400 6 mprj_dat_o[0]
port 647 nsew signal tristate
rlabel metal2 s 465538 163200 465594 164400 6 mprj_dat_o[10]
port 648 nsew signal tristate
rlabel metal2 s 468022 163200 468078 164400 6 mprj_dat_o[11]
port 649 nsew signal tristate
rlabel metal2 s 470506 163200 470562 164400 6 mprj_dat_o[12]
port 650 nsew signal tristate
rlabel metal2 s 473082 163200 473138 164400 6 mprj_dat_o[13]
port 651 nsew signal tristate
rlabel metal2 s 475566 163200 475622 164400 6 mprj_dat_o[14]
port 652 nsew signal tristate
rlabel metal2 s 478142 163200 478198 164400 6 mprj_dat_o[15]
port 653 nsew signal tristate
rlabel metal2 s 480626 163200 480682 164400 6 mprj_dat_o[16]
port 654 nsew signal tristate
rlabel metal2 s 483202 163200 483258 164400 6 mprj_dat_o[17]
port 655 nsew signal tristate
rlabel metal2 s 485686 163200 485742 164400 6 mprj_dat_o[18]
port 656 nsew signal tristate
rlabel metal2 s 488170 163200 488226 164400 6 mprj_dat_o[19]
port 657 nsew signal tristate
rlabel metal2 s 440238 163200 440294 164400 6 mprj_dat_o[1]
port 658 nsew signal tristate
rlabel metal2 s 490746 163200 490802 164400 6 mprj_dat_o[20]
port 659 nsew signal tristate
rlabel metal2 s 493230 163200 493286 164400 6 mprj_dat_o[21]
port 660 nsew signal tristate
rlabel metal2 s 495806 163200 495862 164400 6 mprj_dat_o[22]
port 661 nsew signal tristate
rlabel metal2 s 498290 163200 498346 164400 6 mprj_dat_o[23]
port 662 nsew signal tristate
rlabel metal2 s 500866 163200 500922 164400 6 mprj_dat_o[24]
port 663 nsew signal tristate
rlabel metal2 s 503350 163200 503406 164400 6 mprj_dat_o[25]
port 664 nsew signal tristate
rlabel metal2 s 505834 163200 505890 164400 6 mprj_dat_o[26]
port 665 nsew signal tristate
rlabel metal2 s 508410 163200 508466 164400 6 mprj_dat_o[27]
port 666 nsew signal tristate
rlabel metal2 s 510894 163200 510950 164400 6 mprj_dat_o[28]
port 667 nsew signal tristate
rlabel metal2 s 513470 163200 513526 164400 6 mprj_dat_o[29]
port 668 nsew signal tristate
rlabel metal2 s 443642 163200 443698 164400 6 mprj_dat_o[2]
port 669 nsew signal tristate
rlabel metal2 s 515954 163200 516010 164400 6 mprj_dat_o[30]
port 670 nsew signal tristate
rlabel metal2 s 518530 163200 518586 164400 6 mprj_dat_o[31]
port 671 nsew signal tristate
rlabel metal2 s 446954 163200 447010 164400 6 mprj_dat_o[3]
port 672 nsew signal tristate
rlabel metal2 s 450358 163200 450414 164400 6 mprj_dat_o[4]
port 673 nsew signal tristate
rlabel metal2 s 452842 163200 452898 164400 6 mprj_dat_o[5]
port 674 nsew signal tristate
rlabel metal2 s 455418 163200 455474 164400 6 mprj_dat_o[6]
port 675 nsew signal tristate
rlabel metal2 s 457902 163200 457958 164400 6 mprj_dat_o[7]
port 676 nsew signal tristate
rlabel metal2 s 460478 163200 460534 164400 6 mprj_dat_o[8]
port 677 nsew signal tristate
rlabel metal2 s 462962 163200 463018 164400 6 mprj_dat_o[9]
port 678 nsew signal tristate
rlabel metal2 s 437754 163200 437810 164400 6 mprj_sel_o[0]
port 679 nsew signal tristate
rlabel metal2 s 441066 163200 441122 164400 6 mprj_sel_o[1]
port 680 nsew signal tristate
rlabel metal2 s 444470 163200 444526 164400 6 mprj_sel_o[2]
port 681 nsew signal tristate
rlabel metal2 s 447874 163200 447930 164400 6 mprj_sel_o[3]
port 682 nsew signal tristate
rlabel metal2 s 432694 163200 432750 164400 6 mprj_stb_o
port 683 nsew signal tristate
rlabel metal2 s 433522 163200 433578 164400 6 mprj_wb_iena
port 684 nsew signal tristate
rlabel metal2 s 434350 163200 434406 164400 6 mprj_we_o
port 685 nsew signal tristate
rlabel metal3 s 523200 89360 524400 89480 6 qspi_enabled
port 686 nsew signal tristate
rlabel metal3 s 523200 83376 524400 83496 6 ser_rx
port 687 nsew signal input
rlabel metal3 s 523200 84872 524400 84992 6 ser_tx
port 688 nsew signal tristate
rlabel metal3 s 523200 80384 524400 80504 6 spi_csb
port 689 nsew signal tristate
rlabel metal3 s 523200 86368 524400 86488 6 spi_enabled
port 690 nsew signal tristate
rlabel metal3 s 523200 78888 524400 79008 6 spi_sck
port 691 nsew signal tristate
rlabel metal3 s 523200 81880 524400 82000 6 spi_sdi
port 692 nsew signal input
rlabel metal3 s 523200 77392 524400 77512 6 spi_sdo
port 693 nsew signal tristate
rlabel metal3 s 523200 75896 524400 76016 6 spi_sdoenb
port 694 nsew signal tristate
rlabel metal3 s 523200 2184 524400 2304 6 sram_ro_addr[0]
port 695 nsew signal input
rlabel metal3 s 523200 3680 524400 3800 6 sram_ro_addr[1]
port 696 nsew signal input
rlabel metal3 s 523200 5176 524400 5296 6 sram_ro_addr[2]
port 697 nsew signal input
rlabel metal3 s 523200 6672 524400 6792 6 sram_ro_addr[3]
port 698 nsew signal input
rlabel metal3 s 523200 8168 524400 8288 6 sram_ro_addr[4]
port 699 nsew signal input
rlabel metal3 s 523200 9664 524400 9784 6 sram_ro_addr[5]
port 700 nsew signal input
rlabel metal3 s 523200 11160 524400 11280 6 sram_ro_addr[6]
port 701 nsew signal input
rlabel metal3 s 523200 12656 524400 12776 6 sram_ro_addr[7]
port 702 nsew signal input
rlabel metal3 s 523200 14152 524400 14272 6 sram_ro_clk
port 703 nsew signal input
rlabel metal3 s 523200 688 524400 808 6 sram_ro_csb
port 704 nsew signal input
rlabel metal3 s 523200 15648 524400 15768 6 sram_ro_data[0]
port 705 nsew signal tristate
rlabel metal3 s 523200 30744 524400 30864 6 sram_ro_data[10]
port 706 nsew signal tristate
rlabel metal3 s 523200 32240 524400 32360 6 sram_ro_data[11]
port 707 nsew signal tristate
rlabel metal3 s 523200 33736 524400 33856 6 sram_ro_data[12]
port 708 nsew signal tristate
rlabel metal3 s 523200 35232 524400 35352 6 sram_ro_data[13]
port 709 nsew signal tristate
rlabel metal3 s 523200 36728 524400 36848 6 sram_ro_data[14]
port 710 nsew signal tristate
rlabel metal3 s 523200 38224 524400 38344 6 sram_ro_data[15]
port 711 nsew signal tristate
rlabel metal3 s 523200 39720 524400 39840 6 sram_ro_data[16]
port 712 nsew signal tristate
rlabel metal3 s 523200 41216 524400 41336 6 sram_ro_data[17]
port 713 nsew signal tristate
rlabel metal3 s 523200 42712 524400 42832 6 sram_ro_data[18]
port 714 nsew signal tristate
rlabel metal3 s 523200 44208 524400 44328 6 sram_ro_data[19]
port 715 nsew signal tristate
rlabel metal3 s 523200 17144 524400 17264 6 sram_ro_data[1]
port 716 nsew signal tristate
rlabel metal3 s 523200 45704 524400 45824 6 sram_ro_data[20]
port 717 nsew signal tristate
rlabel metal3 s 523200 47200 524400 47320 6 sram_ro_data[21]
port 718 nsew signal tristate
rlabel metal3 s 523200 48832 524400 48952 6 sram_ro_data[22]
port 719 nsew signal tristate
rlabel metal3 s 523200 50328 524400 50448 6 sram_ro_data[23]
port 720 nsew signal tristate
rlabel metal3 s 523200 51824 524400 51944 6 sram_ro_data[24]
port 721 nsew signal tristate
rlabel metal3 s 523200 53320 524400 53440 6 sram_ro_data[25]
port 722 nsew signal tristate
rlabel metal3 s 523200 54816 524400 54936 6 sram_ro_data[26]
port 723 nsew signal tristate
rlabel metal3 s 523200 56312 524400 56432 6 sram_ro_data[27]
port 724 nsew signal tristate
rlabel metal3 s 523200 57808 524400 57928 6 sram_ro_data[28]
port 725 nsew signal tristate
rlabel metal3 s 523200 59304 524400 59424 6 sram_ro_data[29]
port 726 nsew signal tristate
rlabel metal3 s 523200 18640 524400 18760 6 sram_ro_data[2]
port 727 nsew signal tristate
rlabel metal3 s 523200 60800 524400 60920 6 sram_ro_data[30]
port 728 nsew signal tristate
rlabel metal3 s 523200 62296 524400 62416 6 sram_ro_data[31]
port 729 nsew signal tristate
rlabel metal3 s 523200 20136 524400 20256 6 sram_ro_data[3]
port 730 nsew signal tristate
rlabel metal3 s 523200 21632 524400 21752 6 sram_ro_data[4]
port 731 nsew signal tristate
rlabel metal3 s 523200 23128 524400 23248 6 sram_ro_data[5]
port 732 nsew signal tristate
rlabel metal3 s 523200 24760 524400 24880 6 sram_ro_data[6]
port 733 nsew signal tristate
rlabel metal3 s 523200 26256 524400 26376 6 sram_ro_data[7]
port 734 nsew signal tristate
rlabel metal3 s 523200 27752 524400 27872 6 sram_ro_data[8]
port 735 nsew signal tristate
rlabel metal3 s 523200 29248 524400 29368 6 sram_ro_data[9]
port 736 nsew signal tristate
rlabel metal3 s 523200 69776 524400 69896 6 trap
port 737 nsew signal tristate
rlabel metal3 s 523200 87864 524400 87984 6 uart_enabled
port 738 nsew signal tristate
rlabel metal2 s 519358 163200 519414 164400 6 user_irq_ena[0]
port 739 nsew signal tristate
rlabel metal2 s 520186 163200 520242 164400 6 user_irq_ena[1]
port 740 nsew signal tristate
rlabel metal2 s 521014 163200 521070 164400 6 user_irq_ena[2]
port 741 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 524000 164000
<< end >>
