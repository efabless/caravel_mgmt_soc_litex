magic
tech sky130A
magscale 1 2
timestamp 1638311469
<< obsli1 >>
rect 2869 4159 516900 147809
<< obsm1 >>
rect 382 348 523558 158568
<< metal2 >>
rect 386 159200 442 160400
rect 1214 159200 1270 160400
rect 2042 159200 2098 160400
rect 2870 159200 2926 160400
rect 3698 159200 3754 160400
rect 4526 159200 4582 160400
rect 5354 159200 5410 160400
rect 6182 159200 6238 160400
rect 7102 159200 7158 160400
rect 7930 159200 7986 160400
rect 8758 159200 8814 160400
rect 9586 159200 9642 160400
rect 10414 159200 10470 160400
rect 11242 159200 11298 160400
rect 12070 159200 12126 160400
rect 12898 159200 12954 160400
rect 13818 159200 13874 160400
rect 14646 159200 14702 160400
rect 15474 159200 15530 160400
rect 16302 159200 16358 160400
rect 17130 159200 17186 160400
rect 17958 159200 18014 160400
rect 18786 159200 18842 160400
rect 19614 159200 19670 160400
rect 20534 159200 20590 160400
rect 21362 159200 21418 160400
rect 22190 159200 22246 160400
rect 23018 159200 23074 160400
rect 23846 159200 23902 160400
rect 24674 159200 24730 160400
rect 25502 159200 25558 160400
rect 26330 159200 26386 160400
rect 27250 159200 27306 160400
rect 28078 159200 28134 160400
rect 28906 159200 28962 160400
rect 29734 159200 29790 160400
rect 30562 159200 30618 160400
rect 31390 159200 31446 160400
rect 32218 159200 32274 160400
rect 33138 159200 33194 160400
rect 33966 159200 34022 160400
rect 34794 159200 34850 160400
rect 35622 159200 35678 160400
rect 36450 159200 36506 160400
rect 37278 159200 37334 160400
rect 38106 159200 38162 160400
rect 38934 159200 38990 160400
rect 39854 159200 39910 160400
rect 40682 159200 40738 160400
rect 41510 159200 41566 160400
rect 42338 159200 42394 160400
rect 43166 159200 43222 160400
rect 43994 159200 44050 160400
rect 44822 159200 44878 160400
rect 45650 159200 45706 160400
rect 46570 159200 46626 160400
rect 47398 159200 47454 160400
rect 48226 159200 48282 160400
rect 49054 159200 49110 160400
rect 49882 159200 49938 160400
rect 50710 159200 50766 160400
rect 51538 159200 51594 160400
rect 52366 159200 52422 160400
rect 53286 159200 53342 160400
rect 54114 159200 54170 160400
rect 54942 159200 54998 160400
rect 55770 159200 55826 160400
rect 56598 159200 56654 160400
rect 57426 159200 57482 160400
rect 58254 159200 58310 160400
rect 59082 159200 59138 160400
rect 60002 159200 60058 160400
rect 60830 159200 60886 160400
rect 61658 159200 61714 160400
rect 62486 159200 62542 160400
rect 63314 159200 63370 160400
rect 64142 159200 64198 160400
rect 64970 159200 65026 160400
rect 65890 159200 65946 160400
rect 66718 159200 66774 160400
rect 67546 159200 67602 160400
rect 68374 159200 68430 160400
rect 69202 159200 69258 160400
rect 70030 159200 70086 160400
rect 70858 159200 70914 160400
rect 71686 159200 71742 160400
rect 72606 159200 72662 160400
rect 73434 159200 73490 160400
rect 74262 159200 74318 160400
rect 75090 159200 75146 160400
rect 75918 159200 75974 160400
rect 76746 159200 76802 160400
rect 77574 159200 77630 160400
rect 78402 159200 78458 160400
rect 79322 159200 79378 160400
rect 80150 159200 80206 160400
rect 80978 159200 81034 160400
rect 81806 159200 81862 160400
rect 82634 159200 82690 160400
rect 83462 159200 83518 160400
rect 84290 159200 84346 160400
rect 85118 159200 85174 160400
rect 86038 159200 86094 160400
rect 86866 159200 86922 160400
rect 87694 159200 87750 160400
rect 88522 159200 88578 160400
rect 89350 159200 89406 160400
rect 90178 159200 90234 160400
rect 91006 159200 91062 160400
rect 91834 159200 91890 160400
rect 92754 159200 92810 160400
rect 93582 159200 93638 160400
rect 94410 159200 94466 160400
rect 95238 159200 95294 160400
rect 96066 159200 96122 160400
rect 96894 159200 96950 160400
rect 97722 159200 97778 160400
rect 98642 159200 98698 160400
rect 99470 159200 99526 160400
rect 100298 159200 100354 160400
rect 101126 159200 101182 160400
rect 101954 159200 102010 160400
rect 102782 159200 102838 160400
rect 103610 159200 103666 160400
rect 104438 159200 104494 160400
rect 105358 159200 105414 160400
rect 106186 159200 106242 160400
rect 107014 159200 107070 160400
rect 107842 159200 107898 160400
rect 108670 159200 108726 160400
rect 109498 159200 109554 160400
rect 110326 159200 110382 160400
rect 111154 159200 111210 160400
rect 112074 159200 112130 160400
rect 112902 159200 112958 160400
rect 113730 159200 113786 160400
rect 114558 159200 114614 160400
rect 115386 159200 115442 160400
rect 116214 159200 116270 160400
rect 117042 159200 117098 160400
rect 117870 159200 117926 160400
rect 118790 159200 118846 160400
rect 119618 159200 119674 160400
rect 120446 159200 120502 160400
rect 121274 159200 121330 160400
rect 122102 159200 122158 160400
rect 122930 159200 122986 160400
rect 123758 159200 123814 160400
rect 124586 159200 124642 160400
rect 125506 159200 125562 160400
rect 126334 159200 126390 160400
rect 127162 159200 127218 160400
rect 127990 159200 128046 160400
rect 128818 159200 128874 160400
rect 129646 159200 129702 160400
rect 130474 159200 130530 160400
rect 131394 159200 131450 160400
rect 132222 159200 132278 160400
rect 133050 159200 133106 160400
rect 133878 159200 133934 160400
rect 134706 159200 134762 160400
rect 135534 159200 135590 160400
rect 136362 159200 136418 160400
rect 137190 159200 137246 160400
rect 138110 159200 138166 160400
rect 138938 159200 138994 160400
rect 139766 159200 139822 160400
rect 140594 159200 140650 160400
rect 141422 159200 141478 160400
rect 142250 159200 142306 160400
rect 143078 159200 143134 160400
rect 143906 159200 143962 160400
rect 144826 159200 144882 160400
rect 145654 159200 145710 160400
rect 146482 159200 146538 160400
rect 147310 159200 147366 160400
rect 148138 159200 148194 160400
rect 148966 159200 149022 160400
rect 149794 159200 149850 160400
rect 150622 159200 150678 160400
rect 151542 159200 151598 160400
rect 152370 159200 152426 160400
rect 153198 159200 153254 160400
rect 154026 159200 154082 160400
rect 154854 159200 154910 160400
rect 155682 159200 155738 160400
rect 156510 159200 156566 160400
rect 157338 159200 157394 160400
rect 158258 159200 158314 160400
rect 159086 159200 159142 160400
rect 159914 159200 159970 160400
rect 160742 159200 160798 160400
rect 161570 159200 161626 160400
rect 162398 159200 162454 160400
rect 163226 159200 163282 160400
rect 164146 159200 164202 160400
rect 164974 159200 165030 160400
rect 165802 159200 165858 160400
rect 166630 159200 166686 160400
rect 167458 159200 167514 160400
rect 168286 159200 168342 160400
rect 169114 159200 169170 160400
rect 169942 159200 169998 160400
rect 170862 159200 170918 160400
rect 171690 159200 171746 160400
rect 172518 159200 172574 160400
rect 173346 159200 173402 160400
rect 174174 159200 174230 160400
rect 175002 159200 175058 160400
rect 175830 159200 175886 160400
rect 176658 159200 176714 160400
rect 177578 159200 177634 160400
rect 178406 159200 178462 160400
rect 179234 159200 179290 160400
rect 180062 159200 180118 160400
rect 180890 159200 180946 160400
rect 181718 159200 181774 160400
rect 182546 159200 182602 160400
rect 183374 159200 183430 160400
rect 184294 159200 184350 160400
rect 185122 159200 185178 160400
rect 185950 159200 186006 160400
rect 186778 159200 186834 160400
rect 187606 159200 187662 160400
rect 188434 159200 188490 160400
rect 189262 159200 189318 160400
rect 190090 159200 190146 160400
rect 191010 159200 191066 160400
rect 191838 159200 191894 160400
rect 192666 159200 192722 160400
rect 193494 159200 193550 160400
rect 194322 159200 194378 160400
rect 195150 159200 195206 160400
rect 195978 159200 196034 160400
rect 196898 159200 196954 160400
rect 197726 159200 197782 160400
rect 198554 159200 198610 160400
rect 199382 159200 199438 160400
rect 200210 159200 200266 160400
rect 201038 159200 201094 160400
rect 201866 159200 201922 160400
rect 202694 159200 202750 160400
rect 203614 159200 203670 160400
rect 204442 159200 204498 160400
rect 205270 159200 205326 160400
rect 206098 159200 206154 160400
rect 206926 159200 206982 160400
rect 207754 159200 207810 160400
rect 208582 159200 208638 160400
rect 209410 159200 209466 160400
rect 210330 159200 210386 160400
rect 211158 159200 211214 160400
rect 211986 159200 212042 160400
rect 212814 159200 212870 160400
rect 213642 159200 213698 160400
rect 214470 159200 214526 160400
rect 215298 159200 215354 160400
rect 216126 159200 216182 160400
rect 217046 159200 217102 160400
rect 217874 159200 217930 160400
rect 218702 159200 218758 160400
rect 219530 159200 219586 160400
rect 220358 159200 220414 160400
rect 221186 159200 221242 160400
rect 222014 159200 222070 160400
rect 222842 159200 222898 160400
rect 223762 159200 223818 160400
rect 224590 159200 224646 160400
rect 225418 159200 225474 160400
rect 226246 159200 226302 160400
rect 227074 159200 227130 160400
rect 227902 159200 227958 160400
rect 228730 159200 228786 160400
rect 229650 159200 229706 160400
rect 230478 159200 230534 160400
rect 231306 159200 231362 160400
rect 232134 159200 232190 160400
rect 232962 159200 233018 160400
rect 233790 159200 233846 160400
rect 234618 159200 234674 160400
rect 235446 159200 235502 160400
rect 236366 159200 236422 160400
rect 237194 159200 237250 160400
rect 238022 159200 238078 160400
rect 238850 159200 238906 160400
rect 239678 159200 239734 160400
rect 240506 159200 240562 160400
rect 241334 159200 241390 160400
rect 242162 159200 242218 160400
rect 243082 159200 243138 160400
rect 243910 159200 243966 160400
rect 244738 159200 244794 160400
rect 245566 159200 245622 160400
rect 246394 159200 246450 160400
rect 247222 159200 247278 160400
rect 248050 159200 248106 160400
rect 248878 159200 248934 160400
rect 249798 159200 249854 160400
rect 250626 159200 250682 160400
rect 251454 159200 251510 160400
rect 252282 159200 252338 160400
rect 253110 159200 253166 160400
rect 253938 159200 253994 160400
rect 254766 159200 254822 160400
rect 255594 159200 255650 160400
rect 256514 159200 256570 160400
rect 257342 159200 257398 160400
rect 258170 159200 258226 160400
rect 258998 159200 259054 160400
rect 259826 159200 259882 160400
rect 260654 159200 260710 160400
rect 261482 159200 261538 160400
rect 262402 159200 262458 160400
rect 263230 159200 263286 160400
rect 264058 159200 264114 160400
rect 264886 159200 264942 160400
rect 265714 159200 265770 160400
rect 266542 159200 266598 160400
rect 267370 159200 267426 160400
rect 268198 159200 268254 160400
rect 269118 159200 269174 160400
rect 269946 159200 270002 160400
rect 270774 159200 270830 160400
rect 271602 159200 271658 160400
rect 272430 159200 272486 160400
rect 273258 159200 273314 160400
rect 274086 159200 274142 160400
rect 274914 159200 274970 160400
rect 275834 159200 275890 160400
rect 276662 159200 276718 160400
rect 277490 159200 277546 160400
rect 278318 159200 278374 160400
rect 279146 159200 279202 160400
rect 279974 159200 280030 160400
rect 280802 159200 280858 160400
rect 281630 159200 281686 160400
rect 282550 159200 282606 160400
rect 283378 159200 283434 160400
rect 284206 159200 284262 160400
rect 285034 159200 285090 160400
rect 285862 159200 285918 160400
rect 286690 159200 286746 160400
rect 287518 159200 287574 160400
rect 288346 159200 288402 160400
rect 289266 159200 289322 160400
rect 290094 159200 290150 160400
rect 290922 159200 290978 160400
rect 291750 159200 291806 160400
rect 292578 159200 292634 160400
rect 293406 159200 293462 160400
rect 294234 159200 294290 160400
rect 295154 159200 295210 160400
rect 295982 159200 296038 160400
rect 296810 159200 296866 160400
rect 297638 159200 297694 160400
rect 298466 159200 298522 160400
rect 299294 159200 299350 160400
rect 300122 159200 300178 160400
rect 300950 159200 301006 160400
rect 301870 159200 301926 160400
rect 302698 159200 302754 160400
rect 303526 159200 303582 160400
rect 304354 159200 304410 160400
rect 305182 159200 305238 160400
rect 306010 159200 306066 160400
rect 306838 159200 306894 160400
rect 307666 159200 307722 160400
rect 308586 159200 308642 160400
rect 309414 159200 309470 160400
rect 310242 159200 310298 160400
rect 311070 159200 311126 160400
rect 311898 159200 311954 160400
rect 312726 159200 312782 160400
rect 313554 159200 313610 160400
rect 314382 159200 314438 160400
rect 315302 159200 315358 160400
rect 316130 159200 316186 160400
rect 316958 159200 317014 160400
rect 317786 159200 317842 160400
rect 318614 159200 318670 160400
rect 319442 159200 319498 160400
rect 320270 159200 320326 160400
rect 321098 159200 321154 160400
rect 322018 159200 322074 160400
rect 322846 159200 322902 160400
rect 323674 159200 323730 160400
rect 324502 159200 324558 160400
rect 325330 159200 325386 160400
rect 326158 159200 326214 160400
rect 326986 159200 327042 160400
rect 327906 159200 327962 160400
rect 328734 159200 328790 160400
rect 329562 159200 329618 160400
rect 330390 159200 330446 160400
rect 331218 159200 331274 160400
rect 332046 159200 332102 160400
rect 332874 159200 332930 160400
rect 333702 159200 333758 160400
rect 334622 159200 334678 160400
rect 335450 159200 335506 160400
rect 336278 159200 336334 160400
rect 337106 159200 337162 160400
rect 337934 159200 337990 160400
rect 338762 159200 338818 160400
rect 339590 159200 339646 160400
rect 340418 159200 340474 160400
rect 341338 159200 341394 160400
rect 342166 159200 342222 160400
rect 342994 159200 343050 160400
rect 343822 159200 343878 160400
rect 344650 159200 344706 160400
rect 345478 159200 345534 160400
rect 346306 159200 346362 160400
rect 347134 159200 347190 160400
rect 348054 159200 348110 160400
rect 348882 159200 348938 160400
rect 349710 159200 349766 160400
rect 350538 159200 350594 160400
rect 351366 159200 351422 160400
rect 352194 159200 352250 160400
rect 353022 159200 353078 160400
rect 353850 159200 353906 160400
rect 354770 159200 354826 160400
rect 355598 159200 355654 160400
rect 356426 159200 356482 160400
rect 357254 159200 357310 160400
rect 358082 159200 358138 160400
rect 358910 159200 358966 160400
rect 359738 159200 359794 160400
rect 360658 159200 360714 160400
rect 361486 159200 361542 160400
rect 362314 159200 362370 160400
rect 363142 159200 363198 160400
rect 363970 159200 364026 160400
rect 364798 159200 364854 160400
rect 365626 159200 365682 160400
rect 366454 159200 366510 160400
rect 367374 159200 367430 160400
rect 368202 159200 368258 160400
rect 369030 159200 369086 160400
rect 369858 159200 369914 160400
rect 370686 159200 370742 160400
rect 371514 159200 371570 160400
rect 372342 159200 372398 160400
rect 373170 159200 373226 160400
rect 374090 159200 374146 160400
rect 374918 159200 374974 160400
rect 375746 159200 375802 160400
rect 376574 159200 376630 160400
rect 377402 159200 377458 160400
rect 378230 159200 378286 160400
rect 379058 159200 379114 160400
rect 379886 159200 379942 160400
rect 380806 159200 380862 160400
rect 381634 159200 381690 160400
rect 382462 159200 382518 160400
rect 383290 159200 383346 160400
rect 384118 159200 384174 160400
rect 384946 159200 385002 160400
rect 385774 159200 385830 160400
rect 386602 159200 386658 160400
rect 387522 159200 387578 160400
rect 388350 159200 388406 160400
rect 389178 159200 389234 160400
rect 390006 159200 390062 160400
rect 390834 159200 390890 160400
rect 391662 159200 391718 160400
rect 392490 159200 392546 160400
rect 393410 159200 393466 160400
rect 394238 159200 394294 160400
rect 395066 159200 395122 160400
rect 395894 159200 395950 160400
rect 396722 159200 396778 160400
rect 397550 159200 397606 160400
rect 398378 159200 398434 160400
rect 399206 159200 399262 160400
rect 400126 159200 400182 160400
rect 400954 159200 401010 160400
rect 401782 159200 401838 160400
rect 402610 159200 402666 160400
rect 403438 159200 403494 160400
rect 404266 159200 404322 160400
rect 405094 159200 405150 160400
rect 405922 159200 405978 160400
rect 406842 159200 406898 160400
rect 407670 159200 407726 160400
rect 408498 159200 408554 160400
rect 409326 159200 409382 160400
rect 410154 159200 410210 160400
rect 410982 159200 411038 160400
rect 411810 159200 411866 160400
rect 412638 159200 412694 160400
rect 413558 159200 413614 160400
rect 414386 159200 414442 160400
rect 415214 159200 415270 160400
rect 416042 159200 416098 160400
rect 416870 159200 416926 160400
rect 417698 159200 417754 160400
rect 418526 159200 418582 160400
rect 419354 159200 419410 160400
rect 420274 159200 420330 160400
rect 421102 159200 421158 160400
rect 421930 159200 421986 160400
rect 422758 159200 422814 160400
rect 423586 159200 423642 160400
rect 424414 159200 424470 160400
rect 425242 159200 425298 160400
rect 426162 159200 426218 160400
rect 426990 159200 427046 160400
rect 427818 159200 427874 160400
rect 428646 159200 428702 160400
rect 429474 159200 429530 160400
rect 430302 159200 430358 160400
rect 431130 159200 431186 160400
rect 431958 159200 432014 160400
rect 432878 159200 432934 160400
rect 433706 159200 433762 160400
rect 434534 159200 434590 160400
rect 435362 159200 435418 160400
rect 436190 159200 436246 160400
rect 437018 159200 437074 160400
rect 437846 159200 437902 160400
rect 438674 159200 438730 160400
rect 439594 159200 439650 160400
rect 440422 159200 440478 160400
rect 441250 159200 441306 160400
rect 442078 159200 442134 160400
rect 442906 159200 442962 160400
rect 443734 159200 443790 160400
rect 444562 159200 444618 160400
rect 445390 159200 445446 160400
rect 446310 159200 446366 160400
rect 447138 159200 447194 160400
rect 447966 159200 448022 160400
rect 448794 159200 448850 160400
rect 449622 159200 449678 160400
rect 450450 159200 450506 160400
rect 451278 159200 451334 160400
rect 452106 159200 452162 160400
rect 453026 159200 453082 160400
rect 453854 159200 453910 160400
rect 454682 159200 454738 160400
rect 455510 159200 455566 160400
rect 456338 159200 456394 160400
rect 457166 159200 457222 160400
rect 457994 159200 458050 160400
rect 458914 159200 458970 160400
rect 459742 159200 459798 160400
rect 460570 159200 460626 160400
rect 461398 159200 461454 160400
rect 462226 159200 462282 160400
rect 463054 159200 463110 160400
rect 463882 159200 463938 160400
rect 464710 159200 464766 160400
rect 465630 159200 465686 160400
rect 466458 159200 466514 160400
rect 467286 159200 467342 160400
rect 468114 159200 468170 160400
rect 468942 159200 468998 160400
rect 469770 159200 469826 160400
rect 470598 159200 470654 160400
rect 471426 159200 471482 160400
rect 472346 159200 472402 160400
rect 473174 159200 473230 160400
rect 474002 159200 474058 160400
rect 474830 159200 474886 160400
rect 475658 159200 475714 160400
rect 476486 159200 476542 160400
rect 477314 159200 477370 160400
rect 478142 159200 478198 160400
rect 479062 159200 479118 160400
rect 479890 159200 479946 160400
rect 480718 159200 480774 160400
rect 481546 159200 481602 160400
rect 482374 159200 482430 160400
rect 483202 159200 483258 160400
rect 484030 159200 484086 160400
rect 484858 159200 484914 160400
rect 485778 159200 485834 160400
rect 486606 159200 486662 160400
rect 487434 159200 487490 160400
rect 488262 159200 488318 160400
rect 489090 159200 489146 160400
rect 489918 159200 489974 160400
rect 490746 159200 490802 160400
rect 491666 159200 491722 160400
rect 492494 159200 492550 160400
rect 493322 159200 493378 160400
rect 494150 159200 494206 160400
rect 494978 159200 495034 160400
rect 495806 159200 495862 160400
rect 496634 159200 496690 160400
rect 497462 159200 497518 160400
rect 498382 159200 498438 160400
rect 499210 159200 499266 160400
rect 500038 159200 500094 160400
rect 500866 159200 500922 160400
rect 501694 159200 501750 160400
rect 502522 159200 502578 160400
rect 503350 159200 503406 160400
rect 504178 159200 504234 160400
rect 505098 159200 505154 160400
rect 505926 159200 505982 160400
rect 506754 159200 506810 160400
rect 507582 159200 507638 160400
rect 508410 159200 508466 160400
rect 509238 159200 509294 160400
rect 510066 159200 510122 160400
rect 510894 159200 510950 160400
rect 511814 159200 511870 160400
rect 512642 159200 512698 160400
rect 513470 159200 513526 160400
rect 514298 159200 514354 160400
rect 515126 159200 515182 160400
rect 515954 159200 516010 160400
rect 516782 159200 516838 160400
rect 517610 159200 517666 160400
rect 518530 159200 518586 160400
rect 519358 159200 519414 160400
rect 520186 159200 520242 160400
rect 521014 159200 521070 160400
rect 521842 159200 521898 160400
rect 522670 159200 522726 160400
rect 523498 159200 523554 160400
rect 32770 -400 32826 800
rect 98274 -400 98330 800
rect 163778 -400 163834 800
rect 229282 -400 229338 800
rect 294786 -400 294842 800
rect 360290 -400 360346 800
rect 425794 -400 425850 800
rect 491298 -400 491354 800
<< obsm2 >>
rect 498 159144 1158 159338
rect 1326 159144 1986 159338
rect 2154 159144 2814 159338
rect 2982 159144 3642 159338
rect 3810 159144 4470 159338
rect 4638 159144 5298 159338
rect 5466 159144 6126 159338
rect 6294 159144 7046 159338
rect 7214 159144 7874 159338
rect 8042 159144 8702 159338
rect 8870 159144 9530 159338
rect 9698 159144 10358 159338
rect 10526 159144 11186 159338
rect 11354 159144 12014 159338
rect 12182 159144 12842 159338
rect 13010 159144 13762 159338
rect 13930 159144 14590 159338
rect 14758 159144 15418 159338
rect 15586 159144 16246 159338
rect 16414 159144 17074 159338
rect 17242 159144 17902 159338
rect 18070 159144 18730 159338
rect 18898 159144 19558 159338
rect 19726 159144 20478 159338
rect 20646 159144 21306 159338
rect 21474 159144 22134 159338
rect 22302 159144 22962 159338
rect 23130 159144 23790 159338
rect 23958 159144 24618 159338
rect 24786 159144 25446 159338
rect 25614 159144 26274 159338
rect 26442 159144 27194 159338
rect 27362 159144 28022 159338
rect 28190 159144 28850 159338
rect 29018 159144 29678 159338
rect 29846 159144 30506 159338
rect 30674 159144 31334 159338
rect 31502 159144 32162 159338
rect 32330 159144 33082 159338
rect 33250 159144 33910 159338
rect 34078 159144 34738 159338
rect 34906 159144 35566 159338
rect 35734 159144 36394 159338
rect 36562 159144 37222 159338
rect 37390 159144 38050 159338
rect 38218 159144 38878 159338
rect 39046 159144 39798 159338
rect 39966 159144 40626 159338
rect 40794 159144 41454 159338
rect 41622 159144 42282 159338
rect 42450 159144 43110 159338
rect 43278 159144 43938 159338
rect 44106 159144 44766 159338
rect 44934 159144 45594 159338
rect 45762 159144 46514 159338
rect 46682 159144 47342 159338
rect 47510 159144 48170 159338
rect 48338 159144 48998 159338
rect 49166 159144 49826 159338
rect 49994 159144 50654 159338
rect 50822 159144 51482 159338
rect 51650 159144 52310 159338
rect 52478 159144 53230 159338
rect 53398 159144 54058 159338
rect 54226 159144 54886 159338
rect 55054 159144 55714 159338
rect 55882 159144 56542 159338
rect 56710 159144 57370 159338
rect 57538 159144 58198 159338
rect 58366 159144 59026 159338
rect 59194 159144 59946 159338
rect 60114 159144 60774 159338
rect 60942 159144 61602 159338
rect 61770 159144 62430 159338
rect 62598 159144 63258 159338
rect 63426 159144 64086 159338
rect 64254 159144 64914 159338
rect 65082 159144 65834 159338
rect 66002 159144 66662 159338
rect 66830 159144 67490 159338
rect 67658 159144 68318 159338
rect 68486 159144 69146 159338
rect 69314 159144 69974 159338
rect 70142 159144 70802 159338
rect 70970 159144 71630 159338
rect 71798 159144 72550 159338
rect 72718 159144 73378 159338
rect 73546 159144 74206 159338
rect 74374 159144 75034 159338
rect 75202 159144 75862 159338
rect 76030 159144 76690 159338
rect 76858 159144 77518 159338
rect 77686 159144 78346 159338
rect 78514 159144 79266 159338
rect 79434 159144 80094 159338
rect 80262 159144 80922 159338
rect 81090 159144 81750 159338
rect 81918 159144 82578 159338
rect 82746 159144 83406 159338
rect 83574 159144 84234 159338
rect 84402 159144 85062 159338
rect 85230 159144 85982 159338
rect 86150 159144 86810 159338
rect 86978 159144 87638 159338
rect 87806 159144 88466 159338
rect 88634 159144 89294 159338
rect 89462 159144 90122 159338
rect 90290 159144 90950 159338
rect 91118 159144 91778 159338
rect 91946 159144 92698 159338
rect 92866 159144 93526 159338
rect 93694 159144 94354 159338
rect 94522 159144 95182 159338
rect 95350 159144 96010 159338
rect 96178 159144 96838 159338
rect 97006 159144 97666 159338
rect 97834 159144 98586 159338
rect 98754 159144 99414 159338
rect 99582 159144 100242 159338
rect 100410 159144 101070 159338
rect 101238 159144 101898 159338
rect 102066 159144 102726 159338
rect 102894 159144 103554 159338
rect 103722 159144 104382 159338
rect 104550 159144 105302 159338
rect 105470 159144 106130 159338
rect 106298 159144 106958 159338
rect 107126 159144 107786 159338
rect 107954 159144 108614 159338
rect 108782 159144 109442 159338
rect 109610 159144 110270 159338
rect 110438 159144 111098 159338
rect 111266 159144 112018 159338
rect 112186 159144 112846 159338
rect 113014 159144 113674 159338
rect 113842 159144 114502 159338
rect 114670 159144 115330 159338
rect 115498 159144 116158 159338
rect 116326 159144 116986 159338
rect 117154 159144 117814 159338
rect 117982 159144 118734 159338
rect 118902 159144 119562 159338
rect 119730 159144 120390 159338
rect 120558 159144 121218 159338
rect 121386 159144 122046 159338
rect 122214 159144 122874 159338
rect 123042 159144 123702 159338
rect 123870 159144 124530 159338
rect 124698 159144 125450 159338
rect 125618 159144 126278 159338
rect 126446 159144 127106 159338
rect 127274 159144 127934 159338
rect 128102 159144 128762 159338
rect 128930 159144 129590 159338
rect 129758 159144 130418 159338
rect 130586 159144 131338 159338
rect 131506 159144 132166 159338
rect 132334 159144 132994 159338
rect 133162 159144 133822 159338
rect 133990 159144 134650 159338
rect 134818 159144 135478 159338
rect 135646 159144 136306 159338
rect 136474 159144 137134 159338
rect 137302 159144 138054 159338
rect 138222 159144 138882 159338
rect 139050 159144 139710 159338
rect 139878 159144 140538 159338
rect 140706 159144 141366 159338
rect 141534 159144 142194 159338
rect 142362 159144 143022 159338
rect 143190 159144 143850 159338
rect 144018 159144 144770 159338
rect 144938 159144 145598 159338
rect 145766 159144 146426 159338
rect 146594 159144 147254 159338
rect 147422 159144 148082 159338
rect 148250 159144 148910 159338
rect 149078 159144 149738 159338
rect 149906 159144 150566 159338
rect 150734 159144 151486 159338
rect 151654 159144 152314 159338
rect 152482 159144 153142 159338
rect 153310 159144 153970 159338
rect 154138 159144 154798 159338
rect 154966 159144 155626 159338
rect 155794 159144 156454 159338
rect 156622 159144 157282 159338
rect 157450 159144 158202 159338
rect 158370 159144 159030 159338
rect 159198 159144 159858 159338
rect 160026 159144 160686 159338
rect 160854 159144 161514 159338
rect 161682 159144 162342 159338
rect 162510 159144 163170 159338
rect 163338 159144 164090 159338
rect 164258 159144 164918 159338
rect 165086 159144 165746 159338
rect 165914 159144 166574 159338
rect 166742 159144 167402 159338
rect 167570 159144 168230 159338
rect 168398 159144 169058 159338
rect 169226 159144 169886 159338
rect 170054 159144 170806 159338
rect 170974 159144 171634 159338
rect 171802 159144 172462 159338
rect 172630 159144 173290 159338
rect 173458 159144 174118 159338
rect 174286 159144 174946 159338
rect 175114 159144 175774 159338
rect 175942 159144 176602 159338
rect 176770 159144 177522 159338
rect 177690 159144 178350 159338
rect 178518 159144 179178 159338
rect 179346 159144 180006 159338
rect 180174 159144 180834 159338
rect 181002 159144 181662 159338
rect 181830 159144 182490 159338
rect 182658 159144 183318 159338
rect 183486 159144 184238 159338
rect 184406 159144 185066 159338
rect 185234 159144 185894 159338
rect 186062 159144 186722 159338
rect 186890 159144 187550 159338
rect 187718 159144 188378 159338
rect 188546 159144 189206 159338
rect 189374 159144 190034 159338
rect 190202 159144 190954 159338
rect 191122 159144 191782 159338
rect 191950 159144 192610 159338
rect 192778 159144 193438 159338
rect 193606 159144 194266 159338
rect 194434 159144 195094 159338
rect 195262 159144 195922 159338
rect 196090 159144 196842 159338
rect 197010 159144 197670 159338
rect 197838 159144 198498 159338
rect 198666 159144 199326 159338
rect 199494 159144 200154 159338
rect 200322 159144 200982 159338
rect 201150 159144 201810 159338
rect 201978 159144 202638 159338
rect 202806 159144 203558 159338
rect 203726 159144 204386 159338
rect 204554 159144 205214 159338
rect 205382 159144 206042 159338
rect 206210 159144 206870 159338
rect 207038 159144 207698 159338
rect 207866 159144 208526 159338
rect 208694 159144 209354 159338
rect 209522 159144 210274 159338
rect 210442 159144 211102 159338
rect 211270 159144 211930 159338
rect 212098 159144 212758 159338
rect 212926 159144 213586 159338
rect 213754 159144 214414 159338
rect 214582 159144 215242 159338
rect 215410 159144 216070 159338
rect 216238 159144 216990 159338
rect 217158 159144 217818 159338
rect 217986 159144 218646 159338
rect 218814 159144 219474 159338
rect 219642 159144 220302 159338
rect 220470 159144 221130 159338
rect 221298 159144 221958 159338
rect 222126 159144 222786 159338
rect 222954 159144 223706 159338
rect 223874 159144 224534 159338
rect 224702 159144 225362 159338
rect 225530 159144 226190 159338
rect 226358 159144 227018 159338
rect 227186 159144 227846 159338
rect 228014 159144 228674 159338
rect 228842 159144 229594 159338
rect 229762 159144 230422 159338
rect 230590 159144 231250 159338
rect 231418 159144 232078 159338
rect 232246 159144 232906 159338
rect 233074 159144 233734 159338
rect 233902 159144 234562 159338
rect 234730 159144 235390 159338
rect 235558 159144 236310 159338
rect 236478 159144 237138 159338
rect 237306 159144 237966 159338
rect 238134 159144 238794 159338
rect 238962 159144 239622 159338
rect 239790 159144 240450 159338
rect 240618 159144 241278 159338
rect 241446 159144 242106 159338
rect 242274 159144 243026 159338
rect 243194 159144 243854 159338
rect 244022 159144 244682 159338
rect 244850 159144 245510 159338
rect 245678 159144 246338 159338
rect 246506 159144 247166 159338
rect 247334 159144 247994 159338
rect 248162 159144 248822 159338
rect 248990 159144 249742 159338
rect 249910 159144 250570 159338
rect 250738 159144 251398 159338
rect 251566 159144 252226 159338
rect 252394 159144 253054 159338
rect 253222 159144 253882 159338
rect 254050 159144 254710 159338
rect 254878 159144 255538 159338
rect 255706 159144 256458 159338
rect 256626 159144 257286 159338
rect 257454 159144 258114 159338
rect 258282 159144 258942 159338
rect 259110 159144 259770 159338
rect 259938 159144 260598 159338
rect 260766 159144 261426 159338
rect 261594 159144 262346 159338
rect 262514 159144 263174 159338
rect 263342 159144 264002 159338
rect 264170 159144 264830 159338
rect 264998 159144 265658 159338
rect 265826 159144 266486 159338
rect 266654 159144 267314 159338
rect 267482 159144 268142 159338
rect 268310 159144 269062 159338
rect 269230 159144 269890 159338
rect 270058 159144 270718 159338
rect 270886 159144 271546 159338
rect 271714 159144 272374 159338
rect 272542 159144 273202 159338
rect 273370 159144 274030 159338
rect 274198 159144 274858 159338
rect 275026 159144 275778 159338
rect 275946 159144 276606 159338
rect 276774 159144 277434 159338
rect 277602 159144 278262 159338
rect 278430 159144 279090 159338
rect 279258 159144 279918 159338
rect 280086 159144 280746 159338
rect 280914 159144 281574 159338
rect 281742 159144 282494 159338
rect 282662 159144 283322 159338
rect 283490 159144 284150 159338
rect 284318 159144 284978 159338
rect 285146 159144 285806 159338
rect 285974 159144 286634 159338
rect 286802 159144 287462 159338
rect 287630 159144 288290 159338
rect 288458 159144 289210 159338
rect 289378 159144 290038 159338
rect 290206 159144 290866 159338
rect 291034 159144 291694 159338
rect 291862 159144 292522 159338
rect 292690 159144 293350 159338
rect 293518 159144 294178 159338
rect 294346 159144 295098 159338
rect 295266 159144 295926 159338
rect 296094 159144 296754 159338
rect 296922 159144 297582 159338
rect 297750 159144 298410 159338
rect 298578 159144 299238 159338
rect 299406 159144 300066 159338
rect 300234 159144 300894 159338
rect 301062 159144 301814 159338
rect 301982 159144 302642 159338
rect 302810 159144 303470 159338
rect 303638 159144 304298 159338
rect 304466 159144 305126 159338
rect 305294 159144 305954 159338
rect 306122 159144 306782 159338
rect 306950 159144 307610 159338
rect 307778 159144 308530 159338
rect 308698 159144 309358 159338
rect 309526 159144 310186 159338
rect 310354 159144 311014 159338
rect 311182 159144 311842 159338
rect 312010 159144 312670 159338
rect 312838 159144 313498 159338
rect 313666 159144 314326 159338
rect 314494 159144 315246 159338
rect 315414 159144 316074 159338
rect 316242 159144 316902 159338
rect 317070 159144 317730 159338
rect 317898 159144 318558 159338
rect 318726 159144 319386 159338
rect 319554 159144 320214 159338
rect 320382 159144 321042 159338
rect 321210 159144 321962 159338
rect 322130 159144 322790 159338
rect 322958 159144 323618 159338
rect 323786 159144 324446 159338
rect 324614 159144 325274 159338
rect 325442 159144 326102 159338
rect 326270 159144 326930 159338
rect 327098 159144 327850 159338
rect 328018 159144 328678 159338
rect 328846 159144 329506 159338
rect 329674 159144 330334 159338
rect 330502 159144 331162 159338
rect 331330 159144 331990 159338
rect 332158 159144 332818 159338
rect 332986 159144 333646 159338
rect 333814 159144 334566 159338
rect 334734 159144 335394 159338
rect 335562 159144 336222 159338
rect 336390 159144 337050 159338
rect 337218 159144 337878 159338
rect 338046 159144 338706 159338
rect 338874 159144 339534 159338
rect 339702 159144 340362 159338
rect 340530 159144 341282 159338
rect 341450 159144 342110 159338
rect 342278 159144 342938 159338
rect 343106 159144 343766 159338
rect 343934 159144 344594 159338
rect 344762 159144 345422 159338
rect 345590 159144 346250 159338
rect 346418 159144 347078 159338
rect 347246 159144 347998 159338
rect 348166 159144 348826 159338
rect 348994 159144 349654 159338
rect 349822 159144 350482 159338
rect 350650 159144 351310 159338
rect 351478 159144 352138 159338
rect 352306 159144 352966 159338
rect 353134 159144 353794 159338
rect 353962 159144 354714 159338
rect 354882 159144 355542 159338
rect 355710 159144 356370 159338
rect 356538 159144 357198 159338
rect 357366 159144 358026 159338
rect 358194 159144 358854 159338
rect 359022 159144 359682 159338
rect 359850 159144 360602 159338
rect 360770 159144 361430 159338
rect 361598 159144 362258 159338
rect 362426 159144 363086 159338
rect 363254 159144 363914 159338
rect 364082 159144 364742 159338
rect 364910 159144 365570 159338
rect 365738 159144 366398 159338
rect 366566 159144 367318 159338
rect 367486 159144 368146 159338
rect 368314 159144 368974 159338
rect 369142 159144 369802 159338
rect 369970 159144 370630 159338
rect 370798 159144 371458 159338
rect 371626 159144 372286 159338
rect 372454 159144 373114 159338
rect 373282 159144 374034 159338
rect 374202 159144 374862 159338
rect 375030 159144 375690 159338
rect 375858 159144 376518 159338
rect 376686 159144 377346 159338
rect 377514 159144 378174 159338
rect 378342 159144 379002 159338
rect 379170 159144 379830 159338
rect 379998 159144 380750 159338
rect 380918 159144 381578 159338
rect 381746 159144 382406 159338
rect 382574 159144 383234 159338
rect 383402 159144 384062 159338
rect 384230 159144 384890 159338
rect 385058 159144 385718 159338
rect 385886 159144 386546 159338
rect 386714 159144 387466 159338
rect 387634 159144 388294 159338
rect 388462 159144 389122 159338
rect 389290 159144 389950 159338
rect 390118 159144 390778 159338
rect 390946 159144 391606 159338
rect 391774 159144 392434 159338
rect 392602 159144 393354 159338
rect 393522 159144 394182 159338
rect 394350 159144 395010 159338
rect 395178 159144 395838 159338
rect 396006 159144 396666 159338
rect 396834 159144 397494 159338
rect 397662 159144 398322 159338
rect 398490 159144 399150 159338
rect 399318 159144 400070 159338
rect 400238 159144 400898 159338
rect 401066 159144 401726 159338
rect 401894 159144 402554 159338
rect 402722 159144 403382 159338
rect 403550 159144 404210 159338
rect 404378 159144 405038 159338
rect 405206 159144 405866 159338
rect 406034 159144 406786 159338
rect 406954 159144 407614 159338
rect 407782 159144 408442 159338
rect 408610 159144 409270 159338
rect 409438 159144 410098 159338
rect 410266 159144 410926 159338
rect 411094 159144 411754 159338
rect 411922 159144 412582 159338
rect 412750 159144 413502 159338
rect 413670 159144 414330 159338
rect 414498 159144 415158 159338
rect 415326 159144 415986 159338
rect 416154 159144 416814 159338
rect 416982 159144 417642 159338
rect 417810 159144 418470 159338
rect 418638 159144 419298 159338
rect 419466 159144 420218 159338
rect 420386 159144 421046 159338
rect 421214 159144 421874 159338
rect 422042 159144 422702 159338
rect 422870 159144 423530 159338
rect 423698 159144 424358 159338
rect 424526 159144 425186 159338
rect 425354 159144 426106 159338
rect 426274 159144 426934 159338
rect 427102 159144 427762 159338
rect 427930 159144 428590 159338
rect 428758 159144 429418 159338
rect 429586 159144 430246 159338
rect 430414 159144 431074 159338
rect 431242 159144 431902 159338
rect 432070 159144 432822 159338
rect 432990 159144 433650 159338
rect 433818 159144 434478 159338
rect 434646 159144 435306 159338
rect 435474 159144 436134 159338
rect 436302 159144 436962 159338
rect 437130 159144 437790 159338
rect 437958 159144 438618 159338
rect 438786 159144 439538 159338
rect 439706 159144 440366 159338
rect 440534 159144 441194 159338
rect 441362 159144 442022 159338
rect 442190 159144 442850 159338
rect 443018 159144 443678 159338
rect 443846 159144 444506 159338
rect 444674 159144 445334 159338
rect 445502 159144 446254 159338
rect 446422 159144 447082 159338
rect 447250 159144 447910 159338
rect 448078 159144 448738 159338
rect 448906 159144 449566 159338
rect 449734 159144 450394 159338
rect 450562 159144 451222 159338
rect 451390 159144 452050 159338
rect 452218 159144 452970 159338
rect 453138 159144 453798 159338
rect 453966 159144 454626 159338
rect 454794 159144 455454 159338
rect 455622 159144 456282 159338
rect 456450 159144 457110 159338
rect 457278 159144 457938 159338
rect 458106 159144 458858 159338
rect 459026 159144 459686 159338
rect 459854 159144 460514 159338
rect 460682 159144 461342 159338
rect 461510 159144 462170 159338
rect 462338 159144 462998 159338
rect 463166 159144 463826 159338
rect 463994 159144 464654 159338
rect 464822 159144 465574 159338
rect 465742 159144 466402 159338
rect 466570 159144 467230 159338
rect 467398 159144 468058 159338
rect 468226 159144 468886 159338
rect 469054 159144 469714 159338
rect 469882 159144 470542 159338
rect 470710 159144 471370 159338
rect 471538 159144 472290 159338
rect 472458 159144 473118 159338
rect 473286 159144 473946 159338
rect 474114 159144 474774 159338
rect 474942 159144 475602 159338
rect 475770 159144 476430 159338
rect 476598 159144 477258 159338
rect 477426 159144 478086 159338
rect 478254 159144 479006 159338
rect 479174 159144 479834 159338
rect 480002 159144 480662 159338
rect 480830 159144 481490 159338
rect 481658 159144 482318 159338
rect 482486 159144 483146 159338
rect 483314 159144 483974 159338
rect 484142 159144 484802 159338
rect 484970 159144 485722 159338
rect 485890 159144 486550 159338
rect 486718 159144 487378 159338
rect 487546 159144 488206 159338
rect 488374 159144 489034 159338
rect 489202 159144 489862 159338
rect 490030 159144 490690 159338
rect 490858 159144 491610 159338
rect 491778 159144 492438 159338
rect 492606 159144 493266 159338
rect 493434 159144 494094 159338
rect 494262 159144 494922 159338
rect 495090 159144 495750 159338
rect 495918 159144 496578 159338
rect 496746 159144 497406 159338
rect 497574 159144 498326 159338
rect 498494 159144 499154 159338
rect 499322 159144 499982 159338
rect 500150 159144 500810 159338
rect 500978 159144 501638 159338
rect 501806 159144 502466 159338
rect 502634 159144 503294 159338
rect 503462 159144 504122 159338
rect 504290 159144 505042 159338
rect 505210 159144 505870 159338
rect 506038 159144 506698 159338
rect 506866 159144 507526 159338
rect 507694 159144 508354 159338
rect 508522 159144 509182 159338
rect 509350 159144 510010 159338
rect 510178 159144 510838 159338
rect 511006 159144 511758 159338
rect 511926 159144 512586 159338
rect 512754 159144 513414 159338
rect 513582 159144 514242 159338
rect 514410 159144 515070 159338
rect 515238 159144 515898 159338
rect 516066 159144 516726 159338
rect 516894 159144 517554 159338
rect 517722 159144 518474 159338
rect 518642 159144 519302 159338
rect 519470 159144 520130 159338
rect 520298 159144 520958 159338
rect 521126 159144 521786 159338
rect 521954 159144 522614 159338
rect 522782 159144 523442 159338
rect 388 856 523552 159144
rect 388 342 32714 856
rect 32882 342 98218 856
rect 98386 342 163722 856
rect 163890 342 229226 856
rect 229394 342 294730 856
rect 294898 342 360234 856
rect 360402 342 425738 856
rect 425906 342 491242 856
rect 491410 342 523552 856
<< metal3 >>
rect 523200 159128 524400 159248
rect 523200 157632 524400 157752
rect 523200 156136 524400 156256
rect 523200 154640 524400 154760
rect 523200 153144 524400 153264
rect 523200 151648 524400 151768
rect 523200 150152 524400 150272
rect 523200 148656 524400 148776
rect 523200 147296 524400 147416
rect 523200 145800 524400 145920
rect 523200 144304 524400 144424
rect 523200 142808 524400 142928
rect 523200 141312 524400 141432
rect 523200 139816 524400 139936
rect 523200 138320 524400 138440
rect 523200 136824 524400 136944
rect 523200 135328 524400 135448
rect 523200 133968 524400 134088
rect 523200 132472 524400 132592
rect 523200 130976 524400 131096
rect 523200 129480 524400 129600
rect 523200 127984 524400 128104
rect 523200 126488 524400 126608
rect 523200 124992 524400 125112
rect 523200 123496 524400 123616
rect 523200 122000 524400 122120
rect 523200 120640 524400 120760
rect 523200 119144 524400 119264
rect 523200 117648 524400 117768
rect 523200 116152 524400 116272
rect 523200 114656 524400 114776
rect 523200 113160 524400 113280
rect 523200 111664 524400 111784
rect 523200 110168 524400 110288
rect 523200 108672 524400 108792
rect 523200 107312 524400 107432
rect 523200 105816 524400 105936
rect 523200 104320 524400 104440
rect 523200 102824 524400 102944
rect 523200 101328 524400 101448
rect 523200 99832 524400 99952
rect 523200 98336 524400 98456
rect 523200 96840 524400 96960
rect 523200 95344 524400 95464
rect 523200 93984 524400 94104
rect 523200 92488 524400 92608
rect 523200 90992 524400 91112
rect 523200 89496 524400 89616
rect 523200 88000 524400 88120
rect 523200 86504 524400 86624
rect 523200 85008 524400 85128
rect 523200 83512 524400 83632
rect 523200 82016 524400 82136
rect 523200 80656 524400 80776
rect 523200 79160 524400 79280
rect 523200 77664 524400 77784
rect 523200 76168 524400 76288
rect 523200 74672 524400 74792
rect 523200 73176 524400 73296
rect 523200 71680 524400 71800
rect 523200 70184 524400 70304
rect 523200 68688 524400 68808
rect 523200 67328 524400 67448
rect 523200 65832 524400 65952
rect 523200 64336 524400 64456
rect 523200 62840 524400 62960
rect 523200 61344 524400 61464
rect 523200 59848 524400 59968
rect 523200 58352 524400 58472
rect 523200 56856 524400 56976
rect 523200 55360 524400 55480
rect 523200 54000 524400 54120
rect 523200 52504 524400 52624
rect 523200 51008 524400 51128
rect 523200 49512 524400 49632
rect 523200 48016 524400 48136
rect 523200 46520 524400 46640
rect 523200 45024 524400 45144
rect 523200 43528 524400 43648
rect 523200 42032 524400 42152
rect 523200 40672 524400 40792
rect 523200 39176 524400 39296
rect 523200 37680 524400 37800
rect 523200 36184 524400 36304
rect 523200 34688 524400 34808
rect 523200 33192 524400 33312
rect 523200 31696 524400 31816
rect 523200 30200 524400 30320
rect 523200 28704 524400 28824
rect 523200 27344 524400 27464
rect 523200 25848 524400 25968
rect 523200 24352 524400 24472
rect 523200 22856 524400 22976
rect 523200 21360 524400 21480
rect 523200 19864 524400 19984
rect 523200 18368 524400 18488
rect 523200 16872 524400 16992
rect 523200 15376 524400 15496
rect 523200 14016 524400 14136
rect 523200 12520 524400 12640
rect 523200 11024 524400 11144
rect 523200 9528 524400 9648
rect 523200 8032 524400 8152
rect 523200 6536 524400 6656
rect 523200 5040 524400 5160
rect 523200 3544 524400 3664
rect 523200 2048 524400 2168
rect 523200 688 524400 808
<< obsm3 >>
rect 2037 159048 523120 159221
rect 2037 157832 523200 159048
rect 2037 157552 523120 157832
rect 2037 156336 523200 157552
rect 2037 156056 523120 156336
rect 2037 154840 523200 156056
rect 2037 154560 523120 154840
rect 2037 153344 523200 154560
rect 2037 153064 523120 153344
rect 2037 151848 523200 153064
rect 2037 151568 523120 151848
rect 2037 150352 523200 151568
rect 2037 150072 523120 150352
rect 2037 148856 523200 150072
rect 2037 148576 523120 148856
rect 2037 147496 523200 148576
rect 2037 147216 523120 147496
rect 2037 146000 523200 147216
rect 2037 145720 523120 146000
rect 2037 144504 523200 145720
rect 2037 144224 523120 144504
rect 2037 143008 523200 144224
rect 2037 142728 523120 143008
rect 2037 141512 523200 142728
rect 2037 141232 523120 141512
rect 2037 140016 523200 141232
rect 2037 139736 523120 140016
rect 2037 138520 523200 139736
rect 2037 138240 523120 138520
rect 2037 137024 523200 138240
rect 2037 136744 523120 137024
rect 2037 135528 523200 136744
rect 2037 135248 523120 135528
rect 2037 134168 523200 135248
rect 2037 133888 523120 134168
rect 2037 132672 523200 133888
rect 2037 132392 523120 132672
rect 2037 131176 523200 132392
rect 2037 130896 523120 131176
rect 2037 129680 523200 130896
rect 2037 129400 523120 129680
rect 2037 128184 523200 129400
rect 2037 127904 523120 128184
rect 2037 126688 523200 127904
rect 2037 126408 523120 126688
rect 2037 125192 523200 126408
rect 2037 124912 523120 125192
rect 2037 123696 523200 124912
rect 2037 123416 523120 123696
rect 2037 122200 523200 123416
rect 2037 121920 523120 122200
rect 2037 120840 523200 121920
rect 2037 120560 523120 120840
rect 2037 119344 523200 120560
rect 2037 119064 523120 119344
rect 2037 117848 523200 119064
rect 2037 117568 523120 117848
rect 2037 116352 523200 117568
rect 2037 116072 523120 116352
rect 2037 114856 523200 116072
rect 2037 114576 523120 114856
rect 2037 113360 523200 114576
rect 2037 113080 523120 113360
rect 2037 111864 523200 113080
rect 2037 111584 523120 111864
rect 2037 110368 523200 111584
rect 2037 110088 523120 110368
rect 2037 108872 523200 110088
rect 2037 108592 523120 108872
rect 2037 107512 523200 108592
rect 2037 107232 523120 107512
rect 2037 106016 523200 107232
rect 2037 105736 523120 106016
rect 2037 104520 523200 105736
rect 2037 104240 523120 104520
rect 2037 103024 523200 104240
rect 2037 102744 523120 103024
rect 2037 101528 523200 102744
rect 2037 101248 523120 101528
rect 2037 100032 523200 101248
rect 2037 99752 523120 100032
rect 2037 98536 523200 99752
rect 2037 98256 523120 98536
rect 2037 97040 523200 98256
rect 2037 96760 523120 97040
rect 2037 95544 523200 96760
rect 2037 95264 523120 95544
rect 2037 94184 523200 95264
rect 2037 93904 523120 94184
rect 2037 92688 523200 93904
rect 2037 92408 523120 92688
rect 2037 91192 523200 92408
rect 2037 90912 523120 91192
rect 2037 89696 523200 90912
rect 2037 89416 523120 89696
rect 2037 88200 523200 89416
rect 2037 87920 523120 88200
rect 2037 86704 523200 87920
rect 2037 86424 523120 86704
rect 2037 85208 523200 86424
rect 2037 84928 523120 85208
rect 2037 83712 523200 84928
rect 2037 83432 523120 83712
rect 2037 82216 523200 83432
rect 2037 81936 523120 82216
rect 2037 80856 523200 81936
rect 2037 80576 523120 80856
rect 2037 79360 523200 80576
rect 2037 79080 523120 79360
rect 2037 77864 523200 79080
rect 2037 77584 523120 77864
rect 2037 76368 523200 77584
rect 2037 76088 523120 76368
rect 2037 74872 523200 76088
rect 2037 74592 523120 74872
rect 2037 73376 523200 74592
rect 2037 73096 523120 73376
rect 2037 71880 523200 73096
rect 2037 71600 523120 71880
rect 2037 70384 523200 71600
rect 2037 70104 523120 70384
rect 2037 68888 523200 70104
rect 2037 68608 523120 68888
rect 2037 67528 523200 68608
rect 2037 67248 523120 67528
rect 2037 66032 523200 67248
rect 2037 65752 523120 66032
rect 2037 64536 523200 65752
rect 2037 64256 523120 64536
rect 2037 63040 523200 64256
rect 2037 62760 523120 63040
rect 2037 61544 523200 62760
rect 2037 61264 523120 61544
rect 2037 60048 523200 61264
rect 2037 59768 523120 60048
rect 2037 58552 523200 59768
rect 2037 58272 523120 58552
rect 2037 57056 523200 58272
rect 2037 56776 523120 57056
rect 2037 55560 523200 56776
rect 2037 55280 523120 55560
rect 2037 54200 523200 55280
rect 2037 53920 523120 54200
rect 2037 52704 523200 53920
rect 2037 52424 523120 52704
rect 2037 51208 523200 52424
rect 2037 50928 523120 51208
rect 2037 49712 523200 50928
rect 2037 49432 523120 49712
rect 2037 48216 523200 49432
rect 2037 47936 523120 48216
rect 2037 46720 523200 47936
rect 2037 46440 523120 46720
rect 2037 45224 523200 46440
rect 2037 44944 523120 45224
rect 2037 43728 523200 44944
rect 2037 43448 523120 43728
rect 2037 42232 523200 43448
rect 2037 41952 523120 42232
rect 2037 40872 523200 41952
rect 2037 40592 523120 40872
rect 2037 39376 523200 40592
rect 2037 39096 523120 39376
rect 2037 37880 523200 39096
rect 2037 37600 523120 37880
rect 2037 36384 523200 37600
rect 2037 36104 523120 36384
rect 2037 34888 523200 36104
rect 2037 34608 523120 34888
rect 2037 33392 523200 34608
rect 2037 33112 523120 33392
rect 2037 31896 523200 33112
rect 2037 31616 523120 31896
rect 2037 30400 523200 31616
rect 2037 30120 523120 30400
rect 2037 28904 523200 30120
rect 2037 28624 523120 28904
rect 2037 27544 523200 28624
rect 2037 27264 523120 27544
rect 2037 26048 523200 27264
rect 2037 25768 523120 26048
rect 2037 24552 523200 25768
rect 2037 24272 523120 24552
rect 2037 23056 523200 24272
rect 2037 22776 523120 23056
rect 2037 21560 523200 22776
rect 2037 21280 523120 21560
rect 2037 20064 523200 21280
rect 2037 19784 523120 20064
rect 2037 18568 523200 19784
rect 2037 18288 523120 18568
rect 2037 17072 523200 18288
rect 2037 16792 523120 17072
rect 2037 15576 523200 16792
rect 2037 15296 523120 15576
rect 2037 14216 523200 15296
rect 2037 13936 523120 14216
rect 2037 12720 523200 13936
rect 2037 12440 523120 12720
rect 2037 11224 523200 12440
rect 2037 10944 523120 11224
rect 2037 9728 523200 10944
rect 2037 9448 523120 9728
rect 2037 8232 523200 9448
rect 2037 7952 523120 8232
rect 2037 6736 523200 7952
rect 2037 6456 523120 6736
rect 2037 5240 523200 6456
rect 2037 4960 523120 5240
rect 2037 3744 523200 4960
rect 2037 3464 523120 3744
rect 2037 2248 523200 3464
rect 2037 1968 523120 2248
rect 2037 888 523200 1968
rect 2037 715 523120 888
<< obsm4 >>
rect 1004 2156 518920 149812
<< metal5 >>
rect 1104 143856 2200 144496
rect 109800 143856 120200 144496
rect 517800 143856 522836 144496
rect 1104 130856 2200 131496
rect 109800 130856 120200 131496
rect 517800 130856 522836 131496
rect 1104 117856 2200 118496
rect 109800 117856 120200 118496
rect 517800 117856 522836 118496
rect 1104 104856 2200 105496
rect 109800 104856 120200 105496
rect 517800 104856 522836 105496
rect 1104 91856 2200 92496
rect 109800 91856 120200 92496
rect 517800 91856 522836 92496
rect 1104 78856 2200 79496
rect 109800 78856 120200 79496
rect 517800 78856 522836 79496
rect 1104 65856 2200 66496
rect 109800 65856 120200 66496
rect 517800 65856 522836 66496
rect 1104 52856 2200 53496
rect 109800 52856 120200 53496
rect 517800 52856 522836 53496
rect 1104 39856 2200 40496
rect 109800 39856 120200 40496
rect 517800 39856 522836 40496
rect 1104 26856 2200 27496
rect 109800 26856 120200 27496
rect 517800 26856 522836 27496
rect 1104 13856 2200 14496
rect 109800 13856 120200 14496
rect 517800 13856 522836 14496
<< obsm5 >>
rect 1004 144816 518920 149812
rect 2520 143536 109480 144816
rect 120520 143536 517480 144816
rect 1004 131816 518920 143536
rect 2520 130536 109480 131816
rect 120520 130536 517480 131816
rect 1004 118816 518920 130536
rect 2520 117536 109480 118816
rect 120520 117536 517480 118816
rect 1004 105816 518920 117536
rect 2520 104536 109480 105816
rect 120520 104536 517480 105816
rect 1004 92816 518920 104536
rect 2520 91536 109480 92816
rect 120520 91536 517480 92816
rect 1004 79816 518920 91536
rect 2520 78536 109480 79816
rect 120520 78536 517480 79816
rect 1004 66816 518920 78536
rect 2520 65536 109480 66816
rect 120520 65536 517480 66816
rect 1004 53816 518920 65536
rect 2520 52536 109480 53816
rect 120520 52536 517480 53816
rect 1004 40816 518920 52536
rect 2520 39536 109480 40816
rect 120520 39536 517480 40816
rect 1004 27816 518920 39536
rect 2520 26536 109480 27816
rect 120520 26536 517480 27816
rect 1004 14816 518920 26536
rect 2520 13536 109480 14816
rect 120520 13536 517480 14816
rect 1004 2156 518920 13536
<< labels >>
rlabel metal5 s 1104 26856 2200 27496 6 VGND
port 1 nsew ground input
rlabel metal5 s 109800 26856 120200 27496 6 VGND
port 1 nsew ground input
rlabel metal5 s 517800 26856 522836 27496 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 52856 2200 53496 6 VGND
port 1 nsew ground input
rlabel metal5 s 109800 52856 120200 53496 6 VGND
port 1 nsew ground input
rlabel metal5 s 517800 52856 522836 53496 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 78856 2200 79496 6 VGND
port 1 nsew ground input
rlabel metal5 s 109800 78856 120200 79496 6 VGND
port 1 nsew ground input
rlabel metal5 s 517800 78856 522836 79496 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 104856 2200 105496 6 VGND
port 1 nsew ground input
rlabel metal5 s 109800 104856 120200 105496 6 VGND
port 1 nsew ground input
rlabel metal5 s 517800 104856 522836 105496 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 130856 2200 131496 6 VGND
port 1 nsew ground input
rlabel metal5 s 109800 130856 120200 131496 6 VGND
port 1 nsew ground input
rlabel metal5 s 517800 130856 522836 131496 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 13856 2200 14496 6 VPWR
port 2 nsew power input
rlabel metal5 s 109800 13856 120200 14496 6 VPWR
port 2 nsew power input
rlabel metal5 s 517800 13856 522836 14496 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 39856 2200 40496 6 VPWR
port 2 nsew power input
rlabel metal5 s 109800 39856 120200 40496 6 VPWR
port 2 nsew power input
rlabel metal5 s 517800 39856 522836 40496 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 65856 2200 66496 6 VPWR
port 2 nsew power input
rlabel metal5 s 109800 65856 120200 66496 6 VPWR
port 2 nsew power input
rlabel metal5 s 517800 65856 522836 66496 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 91856 2200 92496 6 VPWR
port 2 nsew power input
rlabel metal5 s 109800 91856 120200 92496 6 VPWR
port 2 nsew power input
rlabel metal5 s 517800 91856 522836 92496 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 117856 2200 118496 6 VPWR
port 2 nsew power input
rlabel metal5 s 109800 117856 120200 118496 6 VPWR
port 2 nsew power input
rlabel metal5 s 517800 117856 522836 118496 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 143856 2200 144496 6 VPWR
port 2 nsew power input
rlabel metal5 s 109800 143856 120200 144496 6 VPWR
port 2 nsew power input
rlabel metal5 s 517800 143856 522836 144496 6 VPWR
port 2 nsew power input
rlabel metal2 s 294786 -400 294842 800 6 core_clk
port 3 nsew signal input
rlabel metal2 s 98274 -400 98330 800 6 core_rstn
port 4 nsew signal input
rlabel metal3 s 523200 62840 524400 62960 6 debug_in
port 5 nsew signal input
rlabel metal3 s 523200 64336 524400 64456 6 debug_mode
port 6 nsew signal output
rlabel metal3 s 523200 65832 524400 65952 6 debug_oeb
port 7 nsew signal output
rlabel metal3 s 523200 67328 524400 67448 6 debug_out
port 8 nsew signal output
rlabel metal3 s 523200 141312 524400 141432 6 flash_clk
port 9 nsew signal output
rlabel metal3 s 523200 139816 524400 139936 6 flash_csb
port 10 nsew signal output
rlabel metal3 s 523200 142808 524400 142928 6 flash_io0_di
port 11 nsew signal input
rlabel metal3 s 523200 144304 524400 144424 6 flash_io0_do
port 12 nsew signal output
rlabel metal3 s 523200 145800 524400 145920 6 flash_io0_oeb
port 13 nsew signal output
rlabel metal3 s 523200 147296 524400 147416 6 flash_io1_di
port 14 nsew signal input
rlabel metal3 s 523200 148656 524400 148776 6 flash_io1_do
port 15 nsew signal output
rlabel metal3 s 523200 150152 524400 150272 6 flash_io1_oeb
port 16 nsew signal output
rlabel metal3 s 523200 151648 524400 151768 6 flash_io2_di
port 17 nsew signal input
rlabel metal3 s 523200 153144 524400 153264 6 flash_io2_do
port 18 nsew signal output
rlabel metal3 s 523200 154640 524400 154760 6 flash_io2_oeb
port 19 nsew signal output
rlabel metal3 s 523200 156136 524400 156256 6 flash_io3_di
port 20 nsew signal input
rlabel metal3 s 523200 157632 524400 157752 6 flash_io3_do
port 21 nsew signal output
rlabel metal3 s 523200 159128 524400 159248 6 flash_io3_oeb
port 22 nsew signal output
rlabel metal2 s 32770 -400 32826 800 6 gpio_in_pad
port 23 nsew signal input
rlabel metal2 s 163778 -400 163834 800 6 gpio_inenb_pad
port 24 nsew signal output
rlabel metal2 s 229282 -400 229338 800 6 gpio_mode0_pad
port 25 nsew signal output
rlabel metal2 s 360290 -400 360346 800 6 gpio_mode1_pad
port 26 nsew signal output
rlabel metal2 s 425794 -400 425850 800 6 gpio_out_pad
port 27 nsew signal output
rlabel metal2 s 491298 -400 491354 800 6 gpio_outenb_pad
port 28 nsew signal output
rlabel metal3 s 523200 89496 524400 89616 6 hk_ack_i
port 29 nsew signal input
rlabel metal2 s 523498 159200 523554 160400 6 hk_cyc_o
port 30 nsew signal output
rlabel metal3 s 523200 92488 524400 92608 6 hk_dat_i[0]
port 31 nsew signal input
rlabel metal3 s 523200 107312 524400 107432 6 hk_dat_i[10]
port 32 nsew signal input
rlabel metal3 s 523200 108672 524400 108792 6 hk_dat_i[11]
port 33 nsew signal input
rlabel metal3 s 523200 110168 524400 110288 6 hk_dat_i[12]
port 34 nsew signal input
rlabel metal3 s 523200 111664 524400 111784 6 hk_dat_i[13]
port 35 nsew signal input
rlabel metal3 s 523200 113160 524400 113280 6 hk_dat_i[14]
port 36 nsew signal input
rlabel metal3 s 523200 114656 524400 114776 6 hk_dat_i[15]
port 37 nsew signal input
rlabel metal3 s 523200 116152 524400 116272 6 hk_dat_i[16]
port 38 nsew signal input
rlabel metal3 s 523200 117648 524400 117768 6 hk_dat_i[17]
port 39 nsew signal input
rlabel metal3 s 523200 119144 524400 119264 6 hk_dat_i[18]
port 40 nsew signal input
rlabel metal3 s 523200 120640 524400 120760 6 hk_dat_i[19]
port 41 nsew signal input
rlabel metal3 s 523200 93984 524400 94104 6 hk_dat_i[1]
port 42 nsew signal input
rlabel metal3 s 523200 122000 524400 122120 6 hk_dat_i[20]
port 43 nsew signal input
rlabel metal3 s 523200 123496 524400 123616 6 hk_dat_i[21]
port 44 nsew signal input
rlabel metal3 s 523200 124992 524400 125112 6 hk_dat_i[22]
port 45 nsew signal input
rlabel metal3 s 523200 126488 524400 126608 6 hk_dat_i[23]
port 46 nsew signal input
rlabel metal3 s 523200 127984 524400 128104 6 hk_dat_i[24]
port 47 nsew signal input
rlabel metal3 s 523200 129480 524400 129600 6 hk_dat_i[25]
port 48 nsew signal input
rlabel metal3 s 523200 130976 524400 131096 6 hk_dat_i[26]
port 49 nsew signal input
rlabel metal3 s 523200 132472 524400 132592 6 hk_dat_i[27]
port 50 nsew signal input
rlabel metal3 s 523200 133968 524400 134088 6 hk_dat_i[28]
port 51 nsew signal input
rlabel metal3 s 523200 135328 524400 135448 6 hk_dat_i[29]
port 52 nsew signal input
rlabel metal3 s 523200 95344 524400 95464 6 hk_dat_i[2]
port 53 nsew signal input
rlabel metal3 s 523200 136824 524400 136944 6 hk_dat_i[30]
port 54 nsew signal input
rlabel metal3 s 523200 138320 524400 138440 6 hk_dat_i[31]
port 55 nsew signal input
rlabel metal3 s 523200 96840 524400 96960 6 hk_dat_i[3]
port 56 nsew signal input
rlabel metal3 s 523200 98336 524400 98456 6 hk_dat_i[4]
port 57 nsew signal input
rlabel metal3 s 523200 99832 524400 99952 6 hk_dat_i[5]
port 58 nsew signal input
rlabel metal3 s 523200 101328 524400 101448 6 hk_dat_i[6]
port 59 nsew signal input
rlabel metal3 s 523200 102824 524400 102944 6 hk_dat_i[7]
port 60 nsew signal input
rlabel metal3 s 523200 104320 524400 104440 6 hk_dat_i[8]
port 61 nsew signal input
rlabel metal3 s 523200 105816 524400 105936 6 hk_dat_i[9]
port 62 nsew signal input
rlabel metal3 s 523200 90992 524400 91112 6 hk_stb_o
port 63 nsew signal output
rlabel metal2 s 521014 159200 521070 160400 6 irq[0]
port 64 nsew signal input
rlabel metal2 s 521842 159200 521898 160400 6 irq[1]
port 65 nsew signal input
rlabel metal2 s 522670 159200 522726 160400 6 irq[2]
port 66 nsew signal input
rlabel metal3 s 523200 73176 524400 73296 6 irq[3]
port 67 nsew signal input
rlabel metal3 s 523200 71680 524400 71800 6 irq[4]
port 68 nsew signal input
rlabel metal3 s 523200 70184 524400 70304 6 irq[5]
port 69 nsew signal input
rlabel metal2 s 386 159200 442 160400 6 la_iena[0]
port 70 nsew signal output
rlabel metal2 s 336278 159200 336334 160400 6 la_iena[100]
port 71 nsew signal output
rlabel metal2 s 339590 159200 339646 160400 6 la_iena[101]
port 72 nsew signal output
rlabel metal2 s 342994 159200 343050 160400 6 la_iena[102]
port 73 nsew signal output
rlabel metal2 s 346306 159200 346362 160400 6 la_iena[103]
port 74 nsew signal output
rlabel metal2 s 349710 159200 349766 160400 6 la_iena[104]
port 75 nsew signal output
rlabel metal2 s 353022 159200 353078 160400 6 la_iena[105]
port 76 nsew signal output
rlabel metal2 s 356426 159200 356482 160400 6 la_iena[106]
port 77 nsew signal output
rlabel metal2 s 359738 159200 359794 160400 6 la_iena[107]
port 78 nsew signal output
rlabel metal2 s 363142 159200 363198 160400 6 la_iena[108]
port 79 nsew signal output
rlabel metal2 s 366454 159200 366510 160400 6 la_iena[109]
port 80 nsew signal output
rlabel metal2 s 33966 159200 34022 160400 6 la_iena[10]
port 81 nsew signal output
rlabel metal2 s 369858 159200 369914 160400 6 la_iena[110]
port 82 nsew signal output
rlabel metal2 s 373170 159200 373226 160400 6 la_iena[111]
port 83 nsew signal output
rlabel metal2 s 376574 159200 376630 160400 6 la_iena[112]
port 84 nsew signal output
rlabel metal2 s 379886 159200 379942 160400 6 la_iena[113]
port 85 nsew signal output
rlabel metal2 s 383290 159200 383346 160400 6 la_iena[114]
port 86 nsew signal output
rlabel metal2 s 386602 159200 386658 160400 6 la_iena[115]
port 87 nsew signal output
rlabel metal2 s 390006 159200 390062 160400 6 la_iena[116]
port 88 nsew signal output
rlabel metal2 s 393410 159200 393466 160400 6 la_iena[117]
port 89 nsew signal output
rlabel metal2 s 396722 159200 396778 160400 6 la_iena[118]
port 90 nsew signal output
rlabel metal2 s 400126 159200 400182 160400 6 la_iena[119]
port 91 nsew signal output
rlabel metal2 s 37278 159200 37334 160400 6 la_iena[11]
port 92 nsew signal output
rlabel metal2 s 403438 159200 403494 160400 6 la_iena[120]
port 93 nsew signal output
rlabel metal2 s 406842 159200 406898 160400 6 la_iena[121]
port 94 nsew signal output
rlabel metal2 s 410154 159200 410210 160400 6 la_iena[122]
port 95 nsew signal output
rlabel metal2 s 413558 159200 413614 160400 6 la_iena[123]
port 96 nsew signal output
rlabel metal2 s 416870 159200 416926 160400 6 la_iena[124]
port 97 nsew signal output
rlabel metal2 s 420274 159200 420330 160400 6 la_iena[125]
port 98 nsew signal output
rlabel metal2 s 423586 159200 423642 160400 6 la_iena[126]
port 99 nsew signal output
rlabel metal2 s 426990 159200 427046 160400 6 la_iena[127]
port 100 nsew signal output
rlabel metal2 s 40682 159200 40738 160400 6 la_iena[12]
port 101 nsew signal output
rlabel metal2 s 43994 159200 44050 160400 6 la_iena[13]
port 102 nsew signal output
rlabel metal2 s 47398 159200 47454 160400 6 la_iena[14]
port 103 nsew signal output
rlabel metal2 s 50710 159200 50766 160400 6 la_iena[15]
port 104 nsew signal output
rlabel metal2 s 54114 159200 54170 160400 6 la_iena[16]
port 105 nsew signal output
rlabel metal2 s 57426 159200 57482 160400 6 la_iena[17]
port 106 nsew signal output
rlabel metal2 s 60830 159200 60886 160400 6 la_iena[18]
port 107 nsew signal output
rlabel metal2 s 64142 159200 64198 160400 6 la_iena[19]
port 108 nsew signal output
rlabel metal2 s 3698 159200 3754 160400 6 la_iena[1]
port 109 nsew signal output
rlabel metal2 s 67546 159200 67602 160400 6 la_iena[20]
port 110 nsew signal output
rlabel metal2 s 70858 159200 70914 160400 6 la_iena[21]
port 111 nsew signal output
rlabel metal2 s 74262 159200 74318 160400 6 la_iena[22]
port 112 nsew signal output
rlabel metal2 s 77574 159200 77630 160400 6 la_iena[23]
port 113 nsew signal output
rlabel metal2 s 80978 159200 81034 160400 6 la_iena[24]
port 114 nsew signal output
rlabel metal2 s 84290 159200 84346 160400 6 la_iena[25]
port 115 nsew signal output
rlabel metal2 s 87694 159200 87750 160400 6 la_iena[26]
port 116 nsew signal output
rlabel metal2 s 91006 159200 91062 160400 6 la_iena[27]
port 117 nsew signal output
rlabel metal2 s 94410 159200 94466 160400 6 la_iena[28]
port 118 nsew signal output
rlabel metal2 s 97722 159200 97778 160400 6 la_iena[29]
port 119 nsew signal output
rlabel metal2 s 7102 159200 7158 160400 6 la_iena[2]
port 120 nsew signal output
rlabel metal2 s 101126 159200 101182 160400 6 la_iena[30]
port 121 nsew signal output
rlabel metal2 s 104438 159200 104494 160400 6 la_iena[31]
port 122 nsew signal output
rlabel metal2 s 107842 159200 107898 160400 6 la_iena[32]
port 123 nsew signal output
rlabel metal2 s 111154 159200 111210 160400 6 la_iena[33]
port 124 nsew signal output
rlabel metal2 s 114558 159200 114614 160400 6 la_iena[34]
port 125 nsew signal output
rlabel metal2 s 117870 159200 117926 160400 6 la_iena[35]
port 126 nsew signal output
rlabel metal2 s 121274 159200 121330 160400 6 la_iena[36]
port 127 nsew signal output
rlabel metal2 s 124586 159200 124642 160400 6 la_iena[37]
port 128 nsew signal output
rlabel metal2 s 127990 159200 128046 160400 6 la_iena[38]
port 129 nsew signal output
rlabel metal2 s 131394 159200 131450 160400 6 la_iena[39]
port 130 nsew signal output
rlabel metal2 s 10414 159200 10470 160400 6 la_iena[3]
port 131 nsew signal output
rlabel metal2 s 134706 159200 134762 160400 6 la_iena[40]
port 132 nsew signal output
rlabel metal2 s 138110 159200 138166 160400 6 la_iena[41]
port 133 nsew signal output
rlabel metal2 s 141422 159200 141478 160400 6 la_iena[42]
port 134 nsew signal output
rlabel metal2 s 144826 159200 144882 160400 6 la_iena[43]
port 135 nsew signal output
rlabel metal2 s 148138 159200 148194 160400 6 la_iena[44]
port 136 nsew signal output
rlabel metal2 s 151542 159200 151598 160400 6 la_iena[45]
port 137 nsew signal output
rlabel metal2 s 154854 159200 154910 160400 6 la_iena[46]
port 138 nsew signal output
rlabel metal2 s 158258 159200 158314 160400 6 la_iena[47]
port 139 nsew signal output
rlabel metal2 s 161570 159200 161626 160400 6 la_iena[48]
port 140 nsew signal output
rlabel metal2 s 164974 159200 165030 160400 6 la_iena[49]
port 141 nsew signal output
rlabel metal2 s 13818 159200 13874 160400 6 la_iena[4]
port 142 nsew signal output
rlabel metal2 s 168286 159200 168342 160400 6 la_iena[50]
port 143 nsew signal output
rlabel metal2 s 171690 159200 171746 160400 6 la_iena[51]
port 144 nsew signal output
rlabel metal2 s 175002 159200 175058 160400 6 la_iena[52]
port 145 nsew signal output
rlabel metal2 s 178406 159200 178462 160400 6 la_iena[53]
port 146 nsew signal output
rlabel metal2 s 181718 159200 181774 160400 6 la_iena[54]
port 147 nsew signal output
rlabel metal2 s 185122 159200 185178 160400 6 la_iena[55]
port 148 nsew signal output
rlabel metal2 s 188434 159200 188490 160400 6 la_iena[56]
port 149 nsew signal output
rlabel metal2 s 191838 159200 191894 160400 6 la_iena[57]
port 150 nsew signal output
rlabel metal2 s 195150 159200 195206 160400 6 la_iena[58]
port 151 nsew signal output
rlabel metal2 s 198554 159200 198610 160400 6 la_iena[59]
port 152 nsew signal output
rlabel metal2 s 17130 159200 17186 160400 6 la_iena[5]
port 153 nsew signal output
rlabel metal2 s 201866 159200 201922 160400 6 la_iena[60]
port 154 nsew signal output
rlabel metal2 s 205270 159200 205326 160400 6 la_iena[61]
port 155 nsew signal output
rlabel metal2 s 208582 159200 208638 160400 6 la_iena[62]
port 156 nsew signal output
rlabel metal2 s 211986 159200 212042 160400 6 la_iena[63]
port 157 nsew signal output
rlabel metal2 s 215298 159200 215354 160400 6 la_iena[64]
port 158 nsew signal output
rlabel metal2 s 218702 159200 218758 160400 6 la_iena[65]
port 159 nsew signal output
rlabel metal2 s 222014 159200 222070 160400 6 la_iena[66]
port 160 nsew signal output
rlabel metal2 s 225418 159200 225474 160400 6 la_iena[67]
port 161 nsew signal output
rlabel metal2 s 228730 159200 228786 160400 6 la_iena[68]
port 162 nsew signal output
rlabel metal2 s 232134 159200 232190 160400 6 la_iena[69]
port 163 nsew signal output
rlabel metal2 s 20534 159200 20590 160400 6 la_iena[6]
port 164 nsew signal output
rlabel metal2 s 235446 159200 235502 160400 6 la_iena[70]
port 165 nsew signal output
rlabel metal2 s 238850 159200 238906 160400 6 la_iena[71]
port 166 nsew signal output
rlabel metal2 s 242162 159200 242218 160400 6 la_iena[72]
port 167 nsew signal output
rlabel metal2 s 245566 159200 245622 160400 6 la_iena[73]
port 168 nsew signal output
rlabel metal2 s 248878 159200 248934 160400 6 la_iena[74]
port 169 nsew signal output
rlabel metal2 s 252282 159200 252338 160400 6 la_iena[75]
port 170 nsew signal output
rlabel metal2 s 255594 159200 255650 160400 6 la_iena[76]
port 171 nsew signal output
rlabel metal2 s 258998 159200 259054 160400 6 la_iena[77]
port 172 nsew signal output
rlabel metal2 s 262402 159200 262458 160400 6 la_iena[78]
port 173 nsew signal output
rlabel metal2 s 265714 159200 265770 160400 6 la_iena[79]
port 174 nsew signal output
rlabel metal2 s 23846 159200 23902 160400 6 la_iena[7]
port 175 nsew signal output
rlabel metal2 s 269118 159200 269174 160400 6 la_iena[80]
port 176 nsew signal output
rlabel metal2 s 272430 159200 272486 160400 6 la_iena[81]
port 177 nsew signal output
rlabel metal2 s 275834 159200 275890 160400 6 la_iena[82]
port 178 nsew signal output
rlabel metal2 s 279146 159200 279202 160400 6 la_iena[83]
port 179 nsew signal output
rlabel metal2 s 282550 159200 282606 160400 6 la_iena[84]
port 180 nsew signal output
rlabel metal2 s 285862 159200 285918 160400 6 la_iena[85]
port 181 nsew signal output
rlabel metal2 s 289266 159200 289322 160400 6 la_iena[86]
port 182 nsew signal output
rlabel metal2 s 292578 159200 292634 160400 6 la_iena[87]
port 183 nsew signal output
rlabel metal2 s 295982 159200 296038 160400 6 la_iena[88]
port 184 nsew signal output
rlabel metal2 s 299294 159200 299350 160400 6 la_iena[89]
port 185 nsew signal output
rlabel metal2 s 27250 159200 27306 160400 6 la_iena[8]
port 186 nsew signal output
rlabel metal2 s 302698 159200 302754 160400 6 la_iena[90]
port 187 nsew signal output
rlabel metal2 s 306010 159200 306066 160400 6 la_iena[91]
port 188 nsew signal output
rlabel metal2 s 309414 159200 309470 160400 6 la_iena[92]
port 189 nsew signal output
rlabel metal2 s 312726 159200 312782 160400 6 la_iena[93]
port 190 nsew signal output
rlabel metal2 s 316130 159200 316186 160400 6 la_iena[94]
port 191 nsew signal output
rlabel metal2 s 319442 159200 319498 160400 6 la_iena[95]
port 192 nsew signal output
rlabel metal2 s 322846 159200 322902 160400 6 la_iena[96]
port 193 nsew signal output
rlabel metal2 s 326158 159200 326214 160400 6 la_iena[97]
port 194 nsew signal output
rlabel metal2 s 329562 159200 329618 160400 6 la_iena[98]
port 195 nsew signal output
rlabel metal2 s 332874 159200 332930 160400 6 la_iena[99]
port 196 nsew signal output
rlabel metal2 s 30562 159200 30618 160400 6 la_iena[9]
port 197 nsew signal output
rlabel metal2 s 1214 159200 1270 160400 6 la_input[0]
port 198 nsew signal input
rlabel metal2 s 337106 159200 337162 160400 6 la_input[100]
port 199 nsew signal input
rlabel metal2 s 340418 159200 340474 160400 6 la_input[101]
port 200 nsew signal input
rlabel metal2 s 343822 159200 343878 160400 6 la_input[102]
port 201 nsew signal input
rlabel metal2 s 347134 159200 347190 160400 6 la_input[103]
port 202 nsew signal input
rlabel metal2 s 350538 159200 350594 160400 6 la_input[104]
port 203 nsew signal input
rlabel metal2 s 353850 159200 353906 160400 6 la_input[105]
port 204 nsew signal input
rlabel metal2 s 357254 159200 357310 160400 6 la_input[106]
port 205 nsew signal input
rlabel metal2 s 360658 159200 360714 160400 6 la_input[107]
port 206 nsew signal input
rlabel metal2 s 363970 159200 364026 160400 6 la_input[108]
port 207 nsew signal input
rlabel metal2 s 367374 159200 367430 160400 6 la_input[109]
port 208 nsew signal input
rlabel metal2 s 34794 159200 34850 160400 6 la_input[10]
port 209 nsew signal input
rlabel metal2 s 370686 159200 370742 160400 6 la_input[110]
port 210 nsew signal input
rlabel metal2 s 374090 159200 374146 160400 6 la_input[111]
port 211 nsew signal input
rlabel metal2 s 377402 159200 377458 160400 6 la_input[112]
port 212 nsew signal input
rlabel metal2 s 380806 159200 380862 160400 6 la_input[113]
port 213 nsew signal input
rlabel metal2 s 384118 159200 384174 160400 6 la_input[114]
port 214 nsew signal input
rlabel metal2 s 387522 159200 387578 160400 6 la_input[115]
port 215 nsew signal input
rlabel metal2 s 390834 159200 390890 160400 6 la_input[116]
port 216 nsew signal input
rlabel metal2 s 394238 159200 394294 160400 6 la_input[117]
port 217 nsew signal input
rlabel metal2 s 397550 159200 397606 160400 6 la_input[118]
port 218 nsew signal input
rlabel metal2 s 400954 159200 401010 160400 6 la_input[119]
port 219 nsew signal input
rlabel metal2 s 38106 159200 38162 160400 6 la_input[11]
port 220 nsew signal input
rlabel metal2 s 404266 159200 404322 160400 6 la_input[120]
port 221 nsew signal input
rlabel metal2 s 407670 159200 407726 160400 6 la_input[121]
port 222 nsew signal input
rlabel metal2 s 410982 159200 411038 160400 6 la_input[122]
port 223 nsew signal input
rlabel metal2 s 414386 159200 414442 160400 6 la_input[123]
port 224 nsew signal input
rlabel metal2 s 417698 159200 417754 160400 6 la_input[124]
port 225 nsew signal input
rlabel metal2 s 421102 159200 421158 160400 6 la_input[125]
port 226 nsew signal input
rlabel metal2 s 424414 159200 424470 160400 6 la_input[126]
port 227 nsew signal input
rlabel metal2 s 427818 159200 427874 160400 6 la_input[127]
port 228 nsew signal input
rlabel metal2 s 41510 159200 41566 160400 6 la_input[12]
port 229 nsew signal input
rlabel metal2 s 44822 159200 44878 160400 6 la_input[13]
port 230 nsew signal input
rlabel metal2 s 48226 159200 48282 160400 6 la_input[14]
port 231 nsew signal input
rlabel metal2 s 51538 159200 51594 160400 6 la_input[15]
port 232 nsew signal input
rlabel metal2 s 54942 159200 54998 160400 6 la_input[16]
port 233 nsew signal input
rlabel metal2 s 58254 159200 58310 160400 6 la_input[17]
port 234 nsew signal input
rlabel metal2 s 61658 159200 61714 160400 6 la_input[18]
port 235 nsew signal input
rlabel metal2 s 64970 159200 65026 160400 6 la_input[19]
port 236 nsew signal input
rlabel metal2 s 4526 159200 4582 160400 6 la_input[1]
port 237 nsew signal input
rlabel metal2 s 68374 159200 68430 160400 6 la_input[20]
port 238 nsew signal input
rlabel metal2 s 71686 159200 71742 160400 6 la_input[21]
port 239 nsew signal input
rlabel metal2 s 75090 159200 75146 160400 6 la_input[22]
port 240 nsew signal input
rlabel metal2 s 78402 159200 78458 160400 6 la_input[23]
port 241 nsew signal input
rlabel metal2 s 81806 159200 81862 160400 6 la_input[24]
port 242 nsew signal input
rlabel metal2 s 85118 159200 85174 160400 6 la_input[25]
port 243 nsew signal input
rlabel metal2 s 88522 159200 88578 160400 6 la_input[26]
port 244 nsew signal input
rlabel metal2 s 91834 159200 91890 160400 6 la_input[27]
port 245 nsew signal input
rlabel metal2 s 95238 159200 95294 160400 6 la_input[28]
port 246 nsew signal input
rlabel metal2 s 98642 159200 98698 160400 6 la_input[29]
port 247 nsew signal input
rlabel metal2 s 7930 159200 7986 160400 6 la_input[2]
port 248 nsew signal input
rlabel metal2 s 101954 159200 102010 160400 6 la_input[30]
port 249 nsew signal input
rlabel metal2 s 105358 159200 105414 160400 6 la_input[31]
port 250 nsew signal input
rlabel metal2 s 108670 159200 108726 160400 6 la_input[32]
port 251 nsew signal input
rlabel metal2 s 112074 159200 112130 160400 6 la_input[33]
port 252 nsew signal input
rlabel metal2 s 115386 159200 115442 160400 6 la_input[34]
port 253 nsew signal input
rlabel metal2 s 118790 159200 118846 160400 6 la_input[35]
port 254 nsew signal input
rlabel metal2 s 122102 159200 122158 160400 6 la_input[36]
port 255 nsew signal input
rlabel metal2 s 125506 159200 125562 160400 6 la_input[37]
port 256 nsew signal input
rlabel metal2 s 128818 159200 128874 160400 6 la_input[38]
port 257 nsew signal input
rlabel metal2 s 132222 159200 132278 160400 6 la_input[39]
port 258 nsew signal input
rlabel metal2 s 11242 159200 11298 160400 6 la_input[3]
port 259 nsew signal input
rlabel metal2 s 135534 159200 135590 160400 6 la_input[40]
port 260 nsew signal input
rlabel metal2 s 138938 159200 138994 160400 6 la_input[41]
port 261 nsew signal input
rlabel metal2 s 142250 159200 142306 160400 6 la_input[42]
port 262 nsew signal input
rlabel metal2 s 145654 159200 145710 160400 6 la_input[43]
port 263 nsew signal input
rlabel metal2 s 148966 159200 149022 160400 6 la_input[44]
port 264 nsew signal input
rlabel metal2 s 152370 159200 152426 160400 6 la_input[45]
port 265 nsew signal input
rlabel metal2 s 155682 159200 155738 160400 6 la_input[46]
port 266 nsew signal input
rlabel metal2 s 159086 159200 159142 160400 6 la_input[47]
port 267 nsew signal input
rlabel metal2 s 162398 159200 162454 160400 6 la_input[48]
port 268 nsew signal input
rlabel metal2 s 165802 159200 165858 160400 6 la_input[49]
port 269 nsew signal input
rlabel metal2 s 14646 159200 14702 160400 6 la_input[4]
port 270 nsew signal input
rlabel metal2 s 169114 159200 169170 160400 6 la_input[50]
port 271 nsew signal input
rlabel metal2 s 172518 159200 172574 160400 6 la_input[51]
port 272 nsew signal input
rlabel metal2 s 175830 159200 175886 160400 6 la_input[52]
port 273 nsew signal input
rlabel metal2 s 179234 159200 179290 160400 6 la_input[53]
port 274 nsew signal input
rlabel metal2 s 182546 159200 182602 160400 6 la_input[54]
port 275 nsew signal input
rlabel metal2 s 185950 159200 186006 160400 6 la_input[55]
port 276 nsew signal input
rlabel metal2 s 189262 159200 189318 160400 6 la_input[56]
port 277 nsew signal input
rlabel metal2 s 192666 159200 192722 160400 6 la_input[57]
port 278 nsew signal input
rlabel metal2 s 195978 159200 196034 160400 6 la_input[58]
port 279 nsew signal input
rlabel metal2 s 199382 159200 199438 160400 6 la_input[59]
port 280 nsew signal input
rlabel metal2 s 17958 159200 18014 160400 6 la_input[5]
port 281 nsew signal input
rlabel metal2 s 202694 159200 202750 160400 6 la_input[60]
port 282 nsew signal input
rlabel metal2 s 206098 159200 206154 160400 6 la_input[61]
port 283 nsew signal input
rlabel metal2 s 209410 159200 209466 160400 6 la_input[62]
port 284 nsew signal input
rlabel metal2 s 212814 159200 212870 160400 6 la_input[63]
port 285 nsew signal input
rlabel metal2 s 216126 159200 216182 160400 6 la_input[64]
port 286 nsew signal input
rlabel metal2 s 219530 159200 219586 160400 6 la_input[65]
port 287 nsew signal input
rlabel metal2 s 222842 159200 222898 160400 6 la_input[66]
port 288 nsew signal input
rlabel metal2 s 226246 159200 226302 160400 6 la_input[67]
port 289 nsew signal input
rlabel metal2 s 229650 159200 229706 160400 6 la_input[68]
port 290 nsew signal input
rlabel metal2 s 232962 159200 233018 160400 6 la_input[69]
port 291 nsew signal input
rlabel metal2 s 21362 159200 21418 160400 6 la_input[6]
port 292 nsew signal input
rlabel metal2 s 236366 159200 236422 160400 6 la_input[70]
port 293 nsew signal input
rlabel metal2 s 239678 159200 239734 160400 6 la_input[71]
port 294 nsew signal input
rlabel metal2 s 243082 159200 243138 160400 6 la_input[72]
port 295 nsew signal input
rlabel metal2 s 246394 159200 246450 160400 6 la_input[73]
port 296 nsew signal input
rlabel metal2 s 249798 159200 249854 160400 6 la_input[74]
port 297 nsew signal input
rlabel metal2 s 253110 159200 253166 160400 6 la_input[75]
port 298 nsew signal input
rlabel metal2 s 256514 159200 256570 160400 6 la_input[76]
port 299 nsew signal input
rlabel metal2 s 259826 159200 259882 160400 6 la_input[77]
port 300 nsew signal input
rlabel metal2 s 263230 159200 263286 160400 6 la_input[78]
port 301 nsew signal input
rlabel metal2 s 266542 159200 266598 160400 6 la_input[79]
port 302 nsew signal input
rlabel metal2 s 24674 159200 24730 160400 6 la_input[7]
port 303 nsew signal input
rlabel metal2 s 269946 159200 270002 160400 6 la_input[80]
port 304 nsew signal input
rlabel metal2 s 273258 159200 273314 160400 6 la_input[81]
port 305 nsew signal input
rlabel metal2 s 276662 159200 276718 160400 6 la_input[82]
port 306 nsew signal input
rlabel metal2 s 279974 159200 280030 160400 6 la_input[83]
port 307 nsew signal input
rlabel metal2 s 283378 159200 283434 160400 6 la_input[84]
port 308 nsew signal input
rlabel metal2 s 286690 159200 286746 160400 6 la_input[85]
port 309 nsew signal input
rlabel metal2 s 290094 159200 290150 160400 6 la_input[86]
port 310 nsew signal input
rlabel metal2 s 293406 159200 293462 160400 6 la_input[87]
port 311 nsew signal input
rlabel metal2 s 296810 159200 296866 160400 6 la_input[88]
port 312 nsew signal input
rlabel metal2 s 300122 159200 300178 160400 6 la_input[89]
port 313 nsew signal input
rlabel metal2 s 28078 159200 28134 160400 6 la_input[8]
port 314 nsew signal input
rlabel metal2 s 303526 159200 303582 160400 6 la_input[90]
port 315 nsew signal input
rlabel metal2 s 306838 159200 306894 160400 6 la_input[91]
port 316 nsew signal input
rlabel metal2 s 310242 159200 310298 160400 6 la_input[92]
port 317 nsew signal input
rlabel metal2 s 313554 159200 313610 160400 6 la_input[93]
port 318 nsew signal input
rlabel metal2 s 316958 159200 317014 160400 6 la_input[94]
port 319 nsew signal input
rlabel metal2 s 320270 159200 320326 160400 6 la_input[95]
port 320 nsew signal input
rlabel metal2 s 323674 159200 323730 160400 6 la_input[96]
port 321 nsew signal input
rlabel metal2 s 326986 159200 327042 160400 6 la_input[97]
port 322 nsew signal input
rlabel metal2 s 330390 159200 330446 160400 6 la_input[98]
port 323 nsew signal input
rlabel metal2 s 333702 159200 333758 160400 6 la_input[99]
port 324 nsew signal input
rlabel metal2 s 31390 159200 31446 160400 6 la_input[9]
port 325 nsew signal input
rlabel metal2 s 2042 159200 2098 160400 6 la_oenb[0]
port 326 nsew signal output
rlabel metal2 s 337934 159200 337990 160400 6 la_oenb[100]
port 327 nsew signal output
rlabel metal2 s 341338 159200 341394 160400 6 la_oenb[101]
port 328 nsew signal output
rlabel metal2 s 344650 159200 344706 160400 6 la_oenb[102]
port 329 nsew signal output
rlabel metal2 s 348054 159200 348110 160400 6 la_oenb[103]
port 330 nsew signal output
rlabel metal2 s 351366 159200 351422 160400 6 la_oenb[104]
port 331 nsew signal output
rlabel metal2 s 354770 159200 354826 160400 6 la_oenb[105]
port 332 nsew signal output
rlabel metal2 s 358082 159200 358138 160400 6 la_oenb[106]
port 333 nsew signal output
rlabel metal2 s 361486 159200 361542 160400 6 la_oenb[107]
port 334 nsew signal output
rlabel metal2 s 364798 159200 364854 160400 6 la_oenb[108]
port 335 nsew signal output
rlabel metal2 s 368202 159200 368258 160400 6 la_oenb[109]
port 336 nsew signal output
rlabel metal2 s 35622 159200 35678 160400 6 la_oenb[10]
port 337 nsew signal output
rlabel metal2 s 371514 159200 371570 160400 6 la_oenb[110]
port 338 nsew signal output
rlabel metal2 s 374918 159200 374974 160400 6 la_oenb[111]
port 339 nsew signal output
rlabel metal2 s 378230 159200 378286 160400 6 la_oenb[112]
port 340 nsew signal output
rlabel metal2 s 381634 159200 381690 160400 6 la_oenb[113]
port 341 nsew signal output
rlabel metal2 s 384946 159200 385002 160400 6 la_oenb[114]
port 342 nsew signal output
rlabel metal2 s 388350 159200 388406 160400 6 la_oenb[115]
port 343 nsew signal output
rlabel metal2 s 391662 159200 391718 160400 6 la_oenb[116]
port 344 nsew signal output
rlabel metal2 s 395066 159200 395122 160400 6 la_oenb[117]
port 345 nsew signal output
rlabel metal2 s 398378 159200 398434 160400 6 la_oenb[118]
port 346 nsew signal output
rlabel metal2 s 401782 159200 401838 160400 6 la_oenb[119]
port 347 nsew signal output
rlabel metal2 s 38934 159200 38990 160400 6 la_oenb[11]
port 348 nsew signal output
rlabel metal2 s 405094 159200 405150 160400 6 la_oenb[120]
port 349 nsew signal output
rlabel metal2 s 408498 159200 408554 160400 6 la_oenb[121]
port 350 nsew signal output
rlabel metal2 s 411810 159200 411866 160400 6 la_oenb[122]
port 351 nsew signal output
rlabel metal2 s 415214 159200 415270 160400 6 la_oenb[123]
port 352 nsew signal output
rlabel metal2 s 418526 159200 418582 160400 6 la_oenb[124]
port 353 nsew signal output
rlabel metal2 s 421930 159200 421986 160400 6 la_oenb[125]
port 354 nsew signal output
rlabel metal2 s 425242 159200 425298 160400 6 la_oenb[126]
port 355 nsew signal output
rlabel metal2 s 428646 159200 428702 160400 6 la_oenb[127]
port 356 nsew signal output
rlabel metal2 s 42338 159200 42394 160400 6 la_oenb[12]
port 357 nsew signal output
rlabel metal2 s 45650 159200 45706 160400 6 la_oenb[13]
port 358 nsew signal output
rlabel metal2 s 49054 159200 49110 160400 6 la_oenb[14]
port 359 nsew signal output
rlabel metal2 s 52366 159200 52422 160400 6 la_oenb[15]
port 360 nsew signal output
rlabel metal2 s 55770 159200 55826 160400 6 la_oenb[16]
port 361 nsew signal output
rlabel metal2 s 59082 159200 59138 160400 6 la_oenb[17]
port 362 nsew signal output
rlabel metal2 s 62486 159200 62542 160400 6 la_oenb[18]
port 363 nsew signal output
rlabel metal2 s 65890 159200 65946 160400 6 la_oenb[19]
port 364 nsew signal output
rlabel metal2 s 5354 159200 5410 160400 6 la_oenb[1]
port 365 nsew signal output
rlabel metal2 s 69202 159200 69258 160400 6 la_oenb[20]
port 366 nsew signal output
rlabel metal2 s 72606 159200 72662 160400 6 la_oenb[21]
port 367 nsew signal output
rlabel metal2 s 75918 159200 75974 160400 6 la_oenb[22]
port 368 nsew signal output
rlabel metal2 s 79322 159200 79378 160400 6 la_oenb[23]
port 369 nsew signal output
rlabel metal2 s 82634 159200 82690 160400 6 la_oenb[24]
port 370 nsew signal output
rlabel metal2 s 86038 159200 86094 160400 6 la_oenb[25]
port 371 nsew signal output
rlabel metal2 s 89350 159200 89406 160400 6 la_oenb[26]
port 372 nsew signal output
rlabel metal2 s 92754 159200 92810 160400 6 la_oenb[27]
port 373 nsew signal output
rlabel metal2 s 96066 159200 96122 160400 6 la_oenb[28]
port 374 nsew signal output
rlabel metal2 s 99470 159200 99526 160400 6 la_oenb[29]
port 375 nsew signal output
rlabel metal2 s 8758 159200 8814 160400 6 la_oenb[2]
port 376 nsew signal output
rlabel metal2 s 102782 159200 102838 160400 6 la_oenb[30]
port 377 nsew signal output
rlabel metal2 s 106186 159200 106242 160400 6 la_oenb[31]
port 378 nsew signal output
rlabel metal2 s 109498 159200 109554 160400 6 la_oenb[32]
port 379 nsew signal output
rlabel metal2 s 112902 159200 112958 160400 6 la_oenb[33]
port 380 nsew signal output
rlabel metal2 s 116214 159200 116270 160400 6 la_oenb[34]
port 381 nsew signal output
rlabel metal2 s 119618 159200 119674 160400 6 la_oenb[35]
port 382 nsew signal output
rlabel metal2 s 122930 159200 122986 160400 6 la_oenb[36]
port 383 nsew signal output
rlabel metal2 s 126334 159200 126390 160400 6 la_oenb[37]
port 384 nsew signal output
rlabel metal2 s 129646 159200 129702 160400 6 la_oenb[38]
port 385 nsew signal output
rlabel metal2 s 133050 159200 133106 160400 6 la_oenb[39]
port 386 nsew signal output
rlabel metal2 s 12070 159200 12126 160400 6 la_oenb[3]
port 387 nsew signal output
rlabel metal2 s 136362 159200 136418 160400 6 la_oenb[40]
port 388 nsew signal output
rlabel metal2 s 139766 159200 139822 160400 6 la_oenb[41]
port 389 nsew signal output
rlabel metal2 s 143078 159200 143134 160400 6 la_oenb[42]
port 390 nsew signal output
rlabel metal2 s 146482 159200 146538 160400 6 la_oenb[43]
port 391 nsew signal output
rlabel metal2 s 149794 159200 149850 160400 6 la_oenb[44]
port 392 nsew signal output
rlabel metal2 s 153198 159200 153254 160400 6 la_oenb[45]
port 393 nsew signal output
rlabel metal2 s 156510 159200 156566 160400 6 la_oenb[46]
port 394 nsew signal output
rlabel metal2 s 159914 159200 159970 160400 6 la_oenb[47]
port 395 nsew signal output
rlabel metal2 s 163226 159200 163282 160400 6 la_oenb[48]
port 396 nsew signal output
rlabel metal2 s 166630 159200 166686 160400 6 la_oenb[49]
port 397 nsew signal output
rlabel metal2 s 15474 159200 15530 160400 6 la_oenb[4]
port 398 nsew signal output
rlabel metal2 s 169942 159200 169998 160400 6 la_oenb[50]
port 399 nsew signal output
rlabel metal2 s 173346 159200 173402 160400 6 la_oenb[51]
port 400 nsew signal output
rlabel metal2 s 176658 159200 176714 160400 6 la_oenb[52]
port 401 nsew signal output
rlabel metal2 s 180062 159200 180118 160400 6 la_oenb[53]
port 402 nsew signal output
rlabel metal2 s 183374 159200 183430 160400 6 la_oenb[54]
port 403 nsew signal output
rlabel metal2 s 186778 159200 186834 160400 6 la_oenb[55]
port 404 nsew signal output
rlabel metal2 s 190090 159200 190146 160400 6 la_oenb[56]
port 405 nsew signal output
rlabel metal2 s 193494 159200 193550 160400 6 la_oenb[57]
port 406 nsew signal output
rlabel metal2 s 196898 159200 196954 160400 6 la_oenb[58]
port 407 nsew signal output
rlabel metal2 s 200210 159200 200266 160400 6 la_oenb[59]
port 408 nsew signal output
rlabel metal2 s 18786 159200 18842 160400 6 la_oenb[5]
port 409 nsew signal output
rlabel metal2 s 203614 159200 203670 160400 6 la_oenb[60]
port 410 nsew signal output
rlabel metal2 s 206926 159200 206982 160400 6 la_oenb[61]
port 411 nsew signal output
rlabel metal2 s 210330 159200 210386 160400 6 la_oenb[62]
port 412 nsew signal output
rlabel metal2 s 213642 159200 213698 160400 6 la_oenb[63]
port 413 nsew signal output
rlabel metal2 s 217046 159200 217102 160400 6 la_oenb[64]
port 414 nsew signal output
rlabel metal2 s 220358 159200 220414 160400 6 la_oenb[65]
port 415 nsew signal output
rlabel metal2 s 223762 159200 223818 160400 6 la_oenb[66]
port 416 nsew signal output
rlabel metal2 s 227074 159200 227130 160400 6 la_oenb[67]
port 417 nsew signal output
rlabel metal2 s 230478 159200 230534 160400 6 la_oenb[68]
port 418 nsew signal output
rlabel metal2 s 233790 159200 233846 160400 6 la_oenb[69]
port 419 nsew signal output
rlabel metal2 s 22190 159200 22246 160400 6 la_oenb[6]
port 420 nsew signal output
rlabel metal2 s 237194 159200 237250 160400 6 la_oenb[70]
port 421 nsew signal output
rlabel metal2 s 240506 159200 240562 160400 6 la_oenb[71]
port 422 nsew signal output
rlabel metal2 s 243910 159200 243966 160400 6 la_oenb[72]
port 423 nsew signal output
rlabel metal2 s 247222 159200 247278 160400 6 la_oenb[73]
port 424 nsew signal output
rlabel metal2 s 250626 159200 250682 160400 6 la_oenb[74]
port 425 nsew signal output
rlabel metal2 s 253938 159200 253994 160400 6 la_oenb[75]
port 426 nsew signal output
rlabel metal2 s 257342 159200 257398 160400 6 la_oenb[76]
port 427 nsew signal output
rlabel metal2 s 260654 159200 260710 160400 6 la_oenb[77]
port 428 nsew signal output
rlabel metal2 s 264058 159200 264114 160400 6 la_oenb[78]
port 429 nsew signal output
rlabel metal2 s 267370 159200 267426 160400 6 la_oenb[79]
port 430 nsew signal output
rlabel metal2 s 25502 159200 25558 160400 6 la_oenb[7]
port 431 nsew signal output
rlabel metal2 s 270774 159200 270830 160400 6 la_oenb[80]
port 432 nsew signal output
rlabel metal2 s 274086 159200 274142 160400 6 la_oenb[81]
port 433 nsew signal output
rlabel metal2 s 277490 159200 277546 160400 6 la_oenb[82]
port 434 nsew signal output
rlabel metal2 s 280802 159200 280858 160400 6 la_oenb[83]
port 435 nsew signal output
rlabel metal2 s 284206 159200 284262 160400 6 la_oenb[84]
port 436 nsew signal output
rlabel metal2 s 287518 159200 287574 160400 6 la_oenb[85]
port 437 nsew signal output
rlabel metal2 s 290922 159200 290978 160400 6 la_oenb[86]
port 438 nsew signal output
rlabel metal2 s 294234 159200 294290 160400 6 la_oenb[87]
port 439 nsew signal output
rlabel metal2 s 297638 159200 297694 160400 6 la_oenb[88]
port 440 nsew signal output
rlabel metal2 s 300950 159200 301006 160400 6 la_oenb[89]
port 441 nsew signal output
rlabel metal2 s 28906 159200 28962 160400 6 la_oenb[8]
port 442 nsew signal output
rlabel metal2 s 304354 159200 304410 160400 6 la_oenb[90]
port 443 nsew signal output
rlabel metal2 s 307666 159200 307722 160400 6 la_oenb[91]
port 444 nsew signal output
rlabel metal2 s 311070 159200 311126 160400 6 la_oenb[92]
port 445 nsew signal output
rlabel metal2 s 314382 159200 314438 160400 6 la_oenb[93]
port 446 nsew signal output
rlabel metal2 s 317786 159200 317842 160400 6 la_oenb[94]
port 447 nsew signal output
rlabel metal2 s 321098 159200 321154 160400 6 la_oenb[95]
port 448 nsew signal output
rlabel metal2 s 324502 159200 324558 160400 6 la_oenb[96]
port 449 nsew signal output
rlabel metal2 s 327906 159200 327962 160400 6 la_oenb[97]
port 450 nsew signal output
rlabel metal2 s 331218 159200 331274 160400 6 la_oenb[98]
port 451 nsew signal output
rlabel metal2 s 334622 159200 334678 160400 6 la_oenb[99]
port 452 nsew signal output
rlabel metal2 s 32218 159200 32274 160400 6 la_oenb[9]
port 453 nsew signal output
rlabel metal2 s 2870 159200 2926 160400 6 la_output[0]
port 454 nsew signal output
rlabel metal2 s 338762 159200 338818 160400 6 la_output[100]
port 455 nsew signal output
rlabel metal2 s 342166 159200 342222 160400 6 la_output[101]
port 456 nsew signal output
rlabel metal2 s 345478 159200 345534 160400 6 la_output[102]
port 457 nsew signal output
rlabel metal2 s 348882 159200 348938 160400 6 la_output[103]
port 458 nsew signal output
rlabel metal2 s 352194 159200 352250 160400 6 la_output[104]
port 459 nsew signal output
rlabel metal2 s 355598 159200 355654 160400 6 la_output[105]
port 460 nsew signal output
rlabel metal2 s 358910 159200 358966 160400 6 la_output[106]
port 461 nsew signal output
rlabel metal2 s 362314 159200 362370 160400 6 la_output[107]
port 462 nsew signal output
rlabel metal2 s 365626 159200 365682 160400 6 la_output[108]
port 463 nsew signal output
rlabel metal2 s 369030 159200 369086 160400 6 la_output[109]
port 464 nsew signal output
rlabel metal2 s 36450 159200 36506 160400 6 la_output[10]
port 465 nsew signal output
rlabel metal2 s 372342 159200 372398 160400 6 la_output[110]
port 466 nsew signal output
rlabel metal2 s 375746 159200 375802 160400 6 la_output[111]
port 467 nsew signal output
rlabel metal2 s 379058 159200 379114 160400 6 la_output[112]
port 468 nsew signal output
rlabel metal2 s 382462 159200 382518 160400 6 la_output[113]
port 469 nsew signal output
rlabel metal2 s 385774 159200 385830 160400 6 la_output[114]
port 470 nsew signal output
rlabel metal2 s 389178 159200 389234 160400 6 la_output[115]
port 471 nsew signal output
rlabel metal2 s 392490 159200 392546 160400 6 la_output[116]
port 472 nsew signal output
rlabel metal2 s 395894 159200 395950 160400 6 la_output[117]
port 473 nsew signal output
rlabel metal2 s 399206 159200 399262 160400 6 la_output[118]
port 474 nsew signal output
rlabel metal2 s 402610 159200 402666 160400 6 la_output[119]
port 475 nsew signal output
rlabel metal2 s 39854 159200 39910 160400 6 la_output[11]
port 476 nsew signal output
rlabel metal2 s 405922 159200 405978 160400 6 la_output[120]
port 477 nsew signal output
rlabel metal2 s 409326 159200 409382 160400 6 la_output[121]
port 478 nsew signal output
rlabel metal2 s 412638 159200 412694 160400 6 la_output[122]
port 479 nsew signal output
rlabel metal2 s 416042 159200 416098 160400 6 la_output[123]
port 480 nsew signal output
rlabel metal2 s 419354 159200 419410 160400 6 la_output[124]
port 481 nsew signal output
rlabel metal2 s 422758 159200 422814 160400 6 la_output[125]
port 482 nsew signal output
rlabel metal2 s 426162 159200 426218 160400 6 la_output[126]
port 483 nsew signal output
rlabel metal2 s 429474 159200 429530 160400 6 la_output[127]
port 484 nsew signal output
rlabel metal2 s 43166 159200 43222 160400 6 la_output[12]
port 485 nsew signal output
rlabel metal2 s 46570 159200 46626 160400 6 la_output[13]
port 486 nsew signal output
rlabel metal2 s 49882 159200 49938 160400 6 la_output[14]
port 487 nsew signal output
rlabel metal2 s 53286 159200 53342 160400 6 la_output[15]
port 488 nsew signal output
rlabel metal2 s 56598 159200 56654 160400 6 la_output[16]
port 489 nsew signal output
rlabel metal2 s 60002 159200 60058 160400 6 la_output[17]
port 490 nsew signal output
rlabel metal2 s 63314 159200 63370 160400 6 la_output[18]
port 491 nsew signal output
rlabel metal2 s 66718 159200 66774 160400 6 la_output[19]
port 492 nsew signal output
rlabel metal2 s 6182 159200 6238 160400 6 la_output[1]
port 493 nsew signal output
rlabel metal2 s 70030 159200 70086 160400 6 la_output[20]
port 494 nsew signal output
rlabel metal2 s 73434 159200 73490 160400 6 la_output[21]
port 495 nsew signal output
rlabel metal2 s 76746 159200 76802 160400 6 la_output[22]
port 496 nsew signal output
rlabel metal2 s 80150 159200 80206 160400 6 la_output[23]
port 497 nsew signal output
rlabel metal2 s 83462 159200 83518 160400 6 la_output[24]
port 498 nsew signal output
rlabel metal2 s 86866 159200 86922 160400 6 la_output[25]
port 499 nsew signal output
rlabel metal2 s 90178 159200 90234 160400 6 la_output[26]
port 500 nsew signal output
rlabel metal2 s 93582 159200 93638 160400 6 la_output[27]
port 501 nsew signal output
rlabel metal2 s 96894 159200 96950 160400 6 la_output[28]
port 502 nsew signal output
rlabel metal2 s 100298 159200 100354 160400 6 la_output[29]
port 503 nsew signal output
rlabel metal2 s 9586 159200 9642 160400 6 la_output[2]
port 504 nsew signal output
rlabel metal2 s 103610 159200 103666 160400 6 la_output[30]
port 505 nsew signal output
rlabel metal2 s 107014 159200 107070 160400 6 la_output[31]
port 506 nsew signal output
rlabel metal2 s 110326 159200 110382 160400 6 la_output[32]
port 507 nsew signal output
rlabel metal2 s 113730 159200 113786 160400 6 la_output[33]
port 508 nsew signal output
rlabel metal2 s 117042 159200 117098 160400 6 la_output[34]
port 509 nsew signal output
rlabel metal2 s 120446 159200 120502 160400 6 la_output[35]
port 510 nsew signal output
rlabel metal2 s 123758 159200 123814 160400 6 la_output[36]
port 511 nsew signal output
rlabel metal2 s 127162 159200 127218 160400 6 la_output[37]
port 512 nsew signal output
rlabel metal2 s 130474 159200 130530 160400 6 la_output[38]
port 513 nsew signal output
rlabel metal2 s 133878 159200 133934 160400 6 la_output[39]
port 514 nsew signal output
rlabel metal2 s 12898 159200 12954 160400 6 la_output[3]
port 515 nsew signal output
rlabel metal2 s 137190 159200 137246 160400 6 la_output[40]
port 516 nsew signal output
rlabel metal2 s 140594 159200 140650 160400 6 la_output[41]
port 517 nsew signal output
rlabel metal2 s 143906 159200 143962 160400 6 la_output[42]
port 518 nsew signal output
rlabel metal2 s 147310 159200 147366 160400 6 la_output[43]
port 519 nsew signal output
rlabel metal2 s 150622 159200 150678 160400 6 la_output[44]
port 520 nsew signal output
rlabel metal2 s 154026 159200 154082 160400 6 la_output[45]
port 521 nsew signal output
rlabel metal2 s 157338 159200 157394 160400 6 la_output[46]
port 522 nsew signal output
rlabel metal2 s 160742 159200 160798 160400 6 la_output[47]
port 523 nsew signal output
rlabel metal2 s 164146 159200 164202 160400 6 la_output[48]
port 524 nsew signal output
rlabel metal2 s 167458 159200 167514 160400 6 la_output[49]
port 525 nsew signal output
rlabel metal2 s 16302 159200 16358 160400 6 la_output[4]
port 526 nsew signal output
rlabel metal2 s 170862 159200 170918 160400 6 la_output[50]
port 527 nsew signal output
rlabel metal2 s 174174 159200 174230 160400 6 la_output[51]
port 528 nsew signal output
rlabel metal2 s 177578 159200 177634 160400 6 la_output[52]
port 529 nsew signal output
rlabel metal2 s 180890 159200 180946 160400 6 la_output[53]
port 530 nsew signal output
rlabel metal2 s 184294 159200 184350 160400 6 la_output[54]
port 531 nsew signal output
rlabel metal2 s 187606 159200 187662 160400 6 la_output[55]
port 532 nsew signal output
rlabel metal2 s 191010 159200 191066 160400 6 la_output[56]
port 533 nsew signal output
rlabel metal2 s 194322 159200 194378 160400 6 la_output[57]
port 534 nsew signal output
rlabel metal2 s 197726 159200 197782 160400 6 la_output[58]
port 535 nsew signal output
rlabel metal2 s 201038 159200 201094 160400 6 la_output[59]
port 536 nsew signal output
rlabel metal2 s 19614 159200 19670 160400 6 la_output[5]
port 537 nsew signal output
rlabel metal2 s 204442 159200 204498 160400 6 la_output[60]
port 538 nsew signal output
rlabel metal2 s 207754 159200 207810 160400 6 la_output[61]
port 539 nsew signal output
rlabel metal2 s 211158 159200 211214 160400 6 la_output[62]
port 540 nsew signal output
rlabel metal2 s 214470 159200 214526 160400 6 la_output[63]
port 541 nsew signal output
rlabel metal2 s 217874 159200 217930 160400 6 la_output[64]
port 542 nsew signal output
rlabel metal2 s 221186 159200 221242 160400 6 la_output[65]
port 543 nsew signal output
rlabel metal2 s 224590 159200 224646 160400 6 la_output[66]
port 544 nsew signal output
rlabel metal2 s 227902 159200 227958 160400 6 la_output[67]
port 545 nsew signal output
rlabel metal2 s 231306 159200 231362 160400 6 la_output[68]
port 546 nsew signal output
rlabel metal2 s 234618 159200 234674 160400 6 la_output[69]
port 547 nsew signal output
rlabel metal2 s 23018 159200 23074 160400 6 la_output[6]
port 548 nsew signal output
rlabel metal2 s 238022 159200 238078 160400 6 la_output[70]
port 549 nsew signal output
rlabel metal2 s 241334 159200 241390 160400 6 la_output[71]
port 550 nsew signal output
rlabel metal2 s 244738 159200 244794 160400 6 la_output[72]
port 551 nsew signal output
rlabel metal2 s 248050 159200 248106 160400 6 la_output[73]
port 552 nsew signal output
rlabel metal2 s 251454 159200 251510 160400 6 la_output[74]
port 553 nsew signal output
rlabel metal2 s 254766 159200 254822 160400 6 la_output[75]
port 554 nsew signal output
rlabel metal2 s 258170 159200 258226 160400 6 la_output[76]
port 555 nsew signal output
rlabel metal2 s 261482 159200 261538 160400 6 la_output[77]
port 556 nsew signal output
rlabel metal2 s 264886 159200 264942 160400 6 la_output[78]
port 557 nsew signal output
rlabel metal2 s 268198 159200 268254 160400 6 la_output[79]
port 558 nsew signal output
rlabel metal2 s 26330 159200 26386 160400 6 la_output[7]
port 559 nsew signal output
rlabel metal2 s 271602 159200 271658 160400 6 la_output[80]
port 560 nsew signal output
rlabel metal2 s 274914 159200 274970 160400 6 la_output[81]
port 561 nsew signal output
rlabel metal2 s 278318 159200 278374 160400 6 la_output[82]
port 562 nsew signal output
rlabel metal2 s 281630 159200 281686 160400 6 la_output[83]
port 563 nsew signal output
rlabel metal2 s 285034 159200 285090 160400 6 la_output[84]
port 564 nsew signal output
rlabel metal2 s 288346 159200 288402 160400 6 la_output[85]
port 565 nsew signal output
rlabel metal2 s 291750 159200 291806 160400 6 la_output[86]
port 566 nsew signal output
rlabel metal2 s 295154 159200 295210 160400 6 la_output[87]
port 567 nsew signal output
rlabel metal2 s 298466 159200 298522 160400 6 la_output[88]
port 568 nsew signal output
rlabel metal2 s 301870 159200 301926 160400 6 la_output[89]
port 569 nsew signal output
rlabel metal2 s 29734 159200 29790 160400 6 la_output[8]
port 570 nsew signal output
rlabel metal2 s 305182 159200 305238 160400 6 la_output[90]
port 571 nsew signal output
rlabel metal2 s 308586 159200 308642 160400 6 la_output[91]
port 572 nsew signal output
rlabel metal2 s 311898 159200 311954 160400 6 la_output[92]
port 573 nsew signal output
rlabel metal2 s 315302 159200 315358 160400 6 la_output[93]
port 574 nsew signal output
rlabel metal2 s 318614 159200 318670 160400 6 la_output[94]
port 575 nsew signal output
rlabel metal2 s 322018 159200 322074 160400 6 la_output[95]
port 576 nsew signal output
rlabel metal2 s 325330 159200 325386 160400 6 la_output[96]
port 577 nsew signal output
rlabel metal2 s 328734 159200 328790 160400 6 la_output[97]
port 578 nsew signal output
rlabel metal2 s 332046 159200 332102 160400 6 la_output[98]
port 579 nsew signal output
rlabel metal2 s 335450 159200 335506 160400 6 la_output[99]
port 580 nsew signal output
rlabel metal2 s 33138 159200 33194 160400 6 la_output[9]
port 581 nsew signal output
rlabel metal2 s 430302 159200 430358 160400 6 mprj_ack_i
port 582 nsew signal input
rlabel metal2 s 434534 159200 434590 160400 6 mprj_adr_o[0]
port 583 nsew signal output
rlabel metal2 s 463054 159200 463110 160400 6 mprj_adr_o[10]
port 584 nsew signal output
rlabel metal2 s 465630 159200 465686 160400 6 mprj_adr_o[11]
port 585 nsew signal output
rlabel metal2 s 468114 159200 468170 160400 6 mprj_adr_o[12]
port 586 nsew signal output
rlabel metal2 s 470598 159200 470654 160400 6 mprj_adr_o[13]
port 587 nsew signal output
rlabel metal2 s 473174 159200 473230 160400 6 mprj_adr_o[14]
port 588 nsew signal output
rlabel metal2 s 475658 159200 475714 160400 6 mprj_adr_o[15]
port 589 nsew signal output
rlabel metal2 s 478142 159200 478198 160400 6 mprj_adr_o[16]
port 590 nsew signal output
rlabel metal2 s 480718 159200 480774 160400 6 mprj_adr_o[17]
port 591 nsew signal output
rlabel metal2 s 483202 159200 483258 160400 6 mprj_adr_o[18]
port 592 nsew signal output
rlabel metal2 s 485778 159200 485834 160400 6 mprj_adr_o[19]
port 593 nsew signal output
rlabel metal2 s 437846 159200 437902 160400 6 mprj_adr_o[1]
port 594 nsew signal output
rlabel metal2 s 488262 159200 488318 160400 6 mprj_adr_o[20]
port 595 nsew signal output
rlabel metal2 s 490746 159200 490802 160400 6 mprj_adr_o[21]
port 596 nsew signal output
rlabel metal2 s 493322 159200 493378 160400 6 mprj_adr_o[22]
port 597 nsew signal output
rlabel metal2 s 495806 159200 495862 160400 6 mprj_adr_o[23]
port 598 nsew signal output
rlabel metal2 s 498382 159200 498438 160400 6 mprj_adr_o[24]
port 599 nsew signal output
rlabel metal2 s 500866 159200 500922 160400 6 mprj_adr_o[25]
port 600 nsew signal output
rlabel metal2 s 503350 159200 503406 160400 6 mprj_adr_o[26]
port 601 nsew signal output
rlabel metal2 s 505926 159200 505982 160400 6 mprj_adr_o[27]
port 602 nsew signal output
rlabel metal2 s 508410 159200 508466 160400 6 mprj_adr_o[28]
port 603 nsew signal output
rlabel metal2 s 510894 159200 510950 160400 6 mprj_adr_o[29]
port 604 nsew signal output
rlabel metal2 s 441250 159200 441306 160400 6 mprj_adr_o[2]
port 605 nsew signal output
rlabel metal2 s 513470 159200 513526 160400 6 mprj_adr_o[30]
port 606 nsew signal output
rlabel metal2 s 515954 159200 516010 160400 6 mprj_adr_o[31]
port 607 nsew signal output
rlabel metal2 s 444562 159200 444618 160400 6 mprj_adr_o[3]
port 608 nsew signal output
rlabel metal2 s 447966 159200 448022 160400 6 mprj_adr_o[4]
port 609 nsew signal output
rlabel metal2 s 450450 159200 450506 160400 6 mprj_adr_o[5]
port 610 nsew signal output
rlabel metal2 s 453026 159200 453082 160400 6 mprj_adr_o[6]
port 611 nsew signal output
rlabel metal2 s 455510 159200 455566 160400 6 mprj_adr_o[7]
port 612 nsew signal output
rlabel metal2 s 457994 159200 458050 160400 6 mprj_adr_o[8]
port 613 nsew signal output
rlabel metal2 s 460570 159200 460626 160400 6 mprj_adr_o[9]
port 614 nsew signal output
rlabel metal2 s 431130 159200 431186 160400 6 mprj_cyc_o
port 615 nsew signal output
rlabel metal2 s 435362 159200 435418 160400 6 mprj_dat_i[0]
port 616 nsew signal input
rlabel metal2 s 463882 159200 463938 160400 6 mprj_dat_i[10]
port 617 nsew signal input
rlabel metal2 s 466458 159200 466514 160400 6 mprj_dat_i[11]
port 618 nsew signal input
rlabel metal2 s 468942 159200 468998 160400 6 mprj_dat_i[12]
port 619 nsew signal input
rlabel metal2 s 471426 159200 471482 160400 6 mprj_dat_i[13]
port 620 nsew signal input
rlabel metal2 s 474002 159200 474058 160400 6 mprj_dat_i[14]
port 621 nsew signal input
rlabel metal2 s 476486 159200 476542 160400 6 mprj_dat_i[15]
port 622 nsew signal input
rlabel metal2 s 479062 159200 479118 160400 6 mprj_dat_i[16]
port 623 nsew signal input
rlabel metal2 s 481546 159200 481602 160400 6 mprj_dat_i[17]
port 624 nsew signal input
rlabel metal2 s 484030 159200 484086 160400 6 mprj_dat_i[18]
port 625 nsew signal input
rlabel metal2 s 486606 159200 486662 160400 6 mprj_dat_i[19]
port 626 nsew signal input
rlabel metal2 s 438674 159200 438730 160400 6 mprj_dat_i[1]
port 627 nsew signal input
rlabel metal2 s 489090 159200 489146 160400 6 mprj_dat_i[20]
port 628 nsew signal input
rlabel metal2 s 491666 159200 491722 160400 6 mprj_dat_i[21]
port 629 nsew signal input
rlabel metal2 s 494150 159200 494206 160400 6 mprj_dat_i[22]
port 630 nsew signal input
rlabel metal2 s 496634 159200 496690 160400 6 mprj_dat_i[23]
port 631 nsew signal input
rlabel metal2 s 499210 159200 499266 160400 6 mprj_dat_i[24]
port 632 nsew signal input
rlabel metal2 s 501694 159200 501750 160400 6 mprj_dat_i[25]
port 633 nsew signal input
rlabel metal2 s 504178 159200 504234 160400 6 mprj_dat_i[26]
port 634 nsew signal input
rlabel metal2 s 506754 159200 506810 160400 6 mprj_dat_i[27]
port 635 nsew signal input
rlabel metal2 s 509238 159200 509294 160400 6 mprj_dat_i[28]
port 636 nsew signal input
rlabel metal2 s 511814 159200 511870 160400 6 mprj_dat_i[29]
port 637 nsew signal input
rlabel metal2 s 442078 159200 442134 160400 6 mprj_dat_i[2]
port 638 nsew signal input
rlabel metal2 s 514298 159200 514354 160400 6 mprj_dat_i[30]
port 639 nsew signal input
rlabel metal2 s 516782 159200 516838 160400 6 mprj_dat_i[31]
port 640 nsew signal input
rlabel metal2 s 445390 159200 445446 160400 6 mprj_dat_i[3]
port 641 nsew signal input
rlabel metal2 s 448794 159200 448850 160400 6 mprj_dat_i[4]
port 642 nsew signal input
rlabel metal2 s 451278 159200 451334 160400 6 mprj_dat_i[5]
port 643 nsew signal input
rlabel metal2 s 453854 159200 453910 160400 6 mprj_dat_i[6]
port 644 nsew signal input
rlabel metal2 s 456338 159200 456394 160400 6 mprj_dat_i[7]
port 645 nsew signal input
rlabel metal2 s 458914 159200 458970 160400 6 mprj_dat_i[8]
port 646 nsew signal input
rlabel metal2 s 461398 159200 461454 160400 6 mprj_dat_i[9]
port 647 nsew signal input
rlabel metal2 s 436190 159200 436246 160400 6 mprj_dat_o[0]
port 648 nsew signal output
rlabel metal2 s 464710 159200 464766 160400 6 mprj_dat_o[10]
port 649 nsew signal output
rlabel metal2 s 467286 159200 467342 160400 6 mprj_dat_o[11]
port 650 nsew signal output
rlabel metal2 s 469770 159200 469826 160400 6 mprj_dat_o[12]
port 651 nsew signal output
rlabel metal2 s 472346 159200 472402 160400 6 mprj_dat_o[13]
port 652 nsew signal output
rlabel metal2 s 474830 159200 474886 160400 6 mprj_dat_o[14]
port 653 nsew signal output
rlabel metal2 s 477314 159200 477370 160400 6 mprj_dat_o[15]
port 654 nsew signal output
rlabel metal2 s 479890 159200 479946 160400 6 mprj_dat_o[16]
port 655 nsew signal output
rlabel metal2 s 482374 159200 482430 160400 6 mprj_dat_o[17]
port 656 nsew signal output
rlabel metal2 s 484858 159200 484914 160400 6 mprj_dat_o[18]
port 657 nsew signal output
rlabel metal2 s 487434 159200 487490 160400 6 mprj_dat_o[19]
port 658 nsew signal output
rlabel metal2 s 439594 159200 439650 160400 6 mprj_dat_o[1]
port 659 nsew signal output
rlabel metal2 s 489918 159200 489974 160400 6 mprj_dat_o[20]
port 660 nsew signal output
rlabel metal2 s 492494 159200 492550 160400 6 mprj_dat_o[21]
port 661 nsew signal output
rlabel metal2 s 494978 159200 495034 160400 6 mprj_dat_o[22]
port 662 nsew signal output
rlabel metal2 s 497462 159200 497518 160400 6 mprj_dat_o[23]
port 663 nsew signal output
rlabel metal2 s 500038 159200 500094 160400 6 mprj_dat_o[24]
port 664 nsew signal output
rlabel metal2 s 502522 159200 502578 160400 6 mprj_dat_o[25]
port 665 nsew signal output
rlabel metal2 s 505098 159200 505154 160400 6 mprj_dat_o[26]
port 666 nsew signal output
rlabel metal2 s 507582 159200 507638 160400 6 mprj_dat_o[27]
port 667 nsew signal output
rlabel metal2 s 510066 159200 510122 160400 6 mprj_dat_o[28]
port 668 nsew signal output
rlabel metal2 s 512642 159200 512698 160400 6 mprj_dat_o[29]
port 669 nsew signal output
rlabel metal2 s 442906 159200 442962 160400 6 mprj_dat_o[2]
port 670 nsew signal output
rlabel metal2 s 515126 159200 515182 160400 6 mprj_dat_o[30]
port 671 nsew signal output
rlabel metal2 s 517610 159200 517666 160400 6 mprj_dat_o[31]
port 672 nsew signal output
rlabel metal2 s 446310 159200 446366 160400 6 mprj_dat_o[3]
port 673 nsew signal output
rlabel metal2 s 449622 159200 449678 160400 6 mprj_dat_o[4]
port 674 nsew signal output
rlabel metal2 s 452106 159200 452162 160400 6 mprj_dat_o[5]
port 675 nsew signal output
rlabel metal2 s 454682 159200 454738 160400 6 mprj_dat_o[6]
port 676 nsew signal output
rlabel metal2 s 457166 159200 457222 160400 6 mprj_dat_o[7]
port 677 nsew signal output
rlabel metal2 s 459742 159200 459798 160400 6 mprj_dat_o[8]
port 678 nsew signal output
rlabel metal2 s 462226 159200 462282 160400 6 mprj_dat_o[9]
port 679 nsew signal output
rlabel metal2 s 437018 159200 437074 160400 6 mprj_sel_o[0]
port 680 nsew signal output
rlabel metal2 s 440422 159200 440478 160400 6 mprj_sel_o[1]
port 681 nsew signal output
rlabel metal2 s 443734 159200 443790 160400 6 mprj_sel_o[2]
port 682 nsew signal output
rlabel metal2 s 447138 159200 447194 160400 6 mprj_sel_o[3]
port 683 nsew signal output
rlabel metal2 s 431958 159200 432014 160400 6 mprj_stb_o
port 684 nsew signal output
rlabel metal2 s 432878 159200 432934 160400 6 mprj_wb_iena
port 685 nsew signal output
rlabel metal2 s 433706 159200 433762 160400 6 mprj_we_o
port 686 nsew signal output
rlabel metal3 s 523200 88000 524400 88120 6 qspi_enabled
port 687 nsew signal output
rlabel metal3 s 523200 82016 524400 82136 6 ser_rx
port 688 nsew signal input
rlabel metal3 s 523200 83512 524400 83632 6 ser_tx
port 689 nsew signal output
rlabel metal3 s 523200 79160 524400 79280 6 spi_csb
port 690 nsew signal output
rlabel metal3 s 523200 85008 524400 85128 6 spi_enabled
port 691 nsew signal output
rlabel metal3 s 523200 77664 524400 77784 6 spi_sck
port 692 nsew signal output
rlabel metal3 s 523200 80656 524400 80776 6 spi_sdi
port 693 nsew signal input
rlabel metal3 s 523200 76168 524400 76288 6 spi_sdo
port 694 nsew signal output
rlabel metal3 s 523200 74672 524400 74792 6 spi_sdoenb
port 695 nsew signal output
rlabel metal3 s 523200 2048 524400 2168 6 sram_ro_addr[0]
port 696 nsew signal input
rlabel metal3 s 523200 3544 524400 3664 6 sram_ro_addr[1]
port 697 nsew signal input
rlabel metal3 s 523200 5040 524400 5160 6 sram_ro_addr[2]
port 698 nsew signal input
rlabel metal3 s 523200 6536 524400 6656 6 sram_ro_addr[3]
port 699 nsew signal input
rlabel metal3 s 523200 8032 524400 8152 6 sram_ro_addr[4]
port 700 nsew signal input
rlabel metal3 s 523200 9528 524400 9648 6 sram_ro_addr[5]
port 701 nsew signal input
rlabel metal3 s 523200 11024 524400 11144 6 sram_ro_addr[6]
port 702 nsew signal input
rlabel metal3 s 523200 12520 524400 12640 6 sram_ro_addr[7]
port 703 nsew signal input
rlabel metal3 s 523200 14016 524400 14136 6 sram_ro_clk
port 704 nsew signal input
rlabel metal3 s 523200 688 524400 808 6 sram_ro_csb
port 705 nsew signal input
rlabel metal3 s 523200 15376 524400 15496 6 sram_ro_data[0]
port 706 nsew signal output
rlabel metal3 s 523200 30200 524400 30320 6 sram_ro_data[10]
port 707 nsew signal output
rlabel metal3 s 523200 31696 524400 31816 6 sram_ro_data[11]
port 708 nsew signal output
rlabel metal3 s 523200 33192 524400 33312 6 sram_ro_data[12]
port 709 nsew signal output
rlabel metal3 s 523200 34688 524400 34808 6 sram_ro_data[13]
port 710 nsew signal output
rlabel metal3 s 523200 36184 524400 36304 6 sram_ro_data[14]
port 711 nsew signal output
rlabel metal3 s 523200 37680 524400 37800 6 sram_ro_data[15]
port 712 nsew signal output
rlabel metal3 s 523200 39176 524400 39296 6 sram_ro_data[16]
port 713 nsew signal output
rlabel metal3 s 523200 40672 524400 40792 6 sram_ro_data[17]
port 714 nsew signal output
rlabel metal3 s 523200 42032 524400 42152 6 sram_ro_data[18]
port 715 nsew signal output
rlabel metal3 s 523200 43528 524400 43648 6 sram_ro_data[19]
port 716 nsew signal output
rlabel metal3 s 523200 16872 524400 16992 6 sram_ro_data[1]
port 717 nsew signal output
rlabel metal3 s 523200 45024 524400 45144 6 sram_ro_data[20]
port 718 nsew signal output
rlabel metal3 s 523200 46520 524400 46640 6 sram_ro_data[21]
port 719 nsew signal output
rlabel metal3 s 523200 48016 524400 48136 6 sram_ro_data[22]
port 720 nsew signal output
rlabel metal3 s 523200 49512 524400 49632 6 sram_ro_data[23]
port 721 nsew signal output
rlabel metal3 s 523200 51008 524400 51128 6 sram_ro_data[24]
port 722 nsew signal output
rlabel metal3 s 523200 52504 524400 52624 6 sram_ro_data[25]
port 723 nsew signal output
rlabel metal3 s 523200 54000 524400 54120 6 sram_ro_data[26]
port 724 nsew signal output
rlabel metal3 s 523200 55360 524400 55480 6 sram_ro_data[27]
port 725 nsew signal output
rlabel metal3 s 523200 56856 524400 56976 6 sram_ro_data[28]
port 726 nsew signal output
rlabel metal3 s 523200 58352 524400 58472 6 sram_ro_data[29]
port 727 nsew signal output
rlabel metal3 s 523200 18368 524400 18488 6 sram_ro_data[2]
port 728 nsew signal output
rlabel metal3 s 523200 59848 524400 59968 6 sram_ro_data[30]
port 729 nsew signal output
rlabel metal3 s 523200 61344 524400 61464 6 sram_ro_data[31]
port 730 nsew signal output
rlabel metal3 s 523200 19864 524400 19984 6 sram_ro_data[3]
port 731 nsew signal output
rlabel metal3 s 523200 21360 524400 21480 6 sram_ro_data[4]
port 732 nsew signal output
rlabel metal3 s 523200 22856 524400 22976 6 sram_ro_data[5]
port 733 nsew signal output
rlabel metal3 s 523200 24352 524400 24472 6 sram_ro_data[6]
port 734 nsew signal output
rlabel metal3 s 523200 25848 524400 25968 6 sram_ro_data[7]
port 735 nsew signal output
rlabel metal3 s 523200 27344 524400 27464 6 sram_ro_data[8]
port 736 nsew signal output
rlabel metal3 s 523200 28704 524400 28824 6 sram_ro_data[9]
port 737 nsew signal output
rlabel metal3 s 523200 68688 524400 68808 6 trap
port 738 nsew signal output
rlabel metal3 s 523200 86504 524400 86624 6 uart_enabled
port 739 nsew signal output
rlabel metal2 s 518530 159200 518586 160400 6 user_irq_ena[0]
port 740 nsew signal output
rlabel metal2 s 519358 159200 519414 160400 6 user_irq_ena[1]
port 741 nsew signal output
rlabel metal2 s 520186 159200 520242 160400 6 user_irq_ena[2]
port 742 nsew signal output
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 524000 160000
string LEFview TRUE
string GDS_FILE /project/openlane/mgmt_core_wrapper/runs/mgmt_core_wrapper/results/magic/mgmt_core_wrapper.gds
string GDS_END 170568968
string GDS_START 169345058
<< end >>

