magic
tech sky130A
magscale 1 2
timestamp 1665629310
<< obsli1 >>
rect 552 527 159068 79985
<< obsm1 >>
rect 290 76 159606 80504
<< metal2 >>
rect 2778 80112 2834 80512
rect 7746 80112 7802 80512
rect 12714 80112 12770 80512
rect 17682 80112 17738 80512
rect 22650 80112 22706 80512
rect 27618 80112 27674 80512
rect 32586 80112 32642 80512
rect 37554 80112 37610 80512
rect 42522 80112 42578 80512
rect 47490 80112 47546 80512
rect 52458 80112 52514 80512
rect 57426 80112 57482 80512
rect 62394 80112 62450 80512
rect 67362 80112 67418 80512
rect 72330 80112 72386 80512
rect 77298 80112 77354 80512
rect 82266 80112 82322 80512
rect 87234 80112 87290 80512
rect 92202 80112 92258 80512
rect 97170 80112 97226 80512
rect 102138 80112 102194 80512
rect 107106 80112 107162 80512
rect 112074 80112 112130 80512
rect 117042 80112 117098 80512
rect 122010 80112 122066 80512
rect 126978 80112 127034 80512
rect 131946 80112 132002 80512
rect 136914 80112 136970 80512
rect 141882 80112 141938 80512
rect 146850 80112 146906 80512
rect 151818 80112 151874 80512
rect 156786 80112 156842 80512
rect 2778 0 2834 400
rect 7746 0 7802 400
rect 12714 0 12770 400
rect 17682 0 17738 400
rect 22650 0 22706 400
rect 27618 0 27674 400
rect 32586 0 32642 400
rect 37554 0 37610 400
rect 42522 0 42578 400
rect 47490 0 47546 400
rect 52458 0 52514 400
rect 57426 0 57482 400
rect 62394 0 62450 400
rect 67362 0 67418 400
rect 72330 0 72386 400
rect 77298 0 77354 400
rect 82266 0 82322 400
rect 87234 0 87290 400
rect 92202 0 92258 400
rect 97170 0 97226 400
rect 102138 0 102194 400
rect 107106 0 107162 400
rect 112074 0 112130 400
rect 117042 0 117098 400
rect 122010 0 122066 400
rect 126978 0 127034 400
rect 131946 0 132002 400
rect 136914 0 136970 400
rect 141882 0 141938 400
rect 146850 0 146906 400
rect 151818 0 151874 400
rect 156786 0 156842 400
<< obsm2 >>
rect 294 80056 2722 80510
rect 2890 80056 7690 80510
rect 7858 80056 12658 80510
rect 12826 80056 17626 80510
rect 17794 80056 22594 80510
rect 22762 80056 27562 80510
rect 27730 80056 32530 80510
rect 32698 80056 37498 80510
rect 37666 80056 42466 80510
rect 42634 80056 47434 80510
rect 47602 80056 52402 80510
rect 52570 80056 57370 80510
rect 57538 80056 62338 80510
rect 62506 80056 67306 80510
rect 67474 80056 72274 80510
rect 72442 80056 77242 80510
rect 77410 80056 82210 80510
rect 82378 80056 87178 80510
rect 87346 80056 92146 80510
rect 92314 80056 97114 80510
rect 97282 80056 102082 80510
rect 102250 80056 107050 80510
rect 107218 80056 112018 80510
rect 112186 80056 116986 80510
rect 117154 80056 121954 80510
rect 122122 80056 126922 80510
rect 127090 80056 131890 80510
rect 132058 80056 136858 80510
rect 137026 80056 141826 80510
rect 141994 80056 146794 80510
rect 146962 80056 151762 80510
rect 151930 80056 156730 80510
rect 156898 80056 159600 80510
rect 294 456 159600 80056
rect 294 31 2722 456
rect 2890 31 7690 456
rect 7858 31 12658 456
rect 12826 31 17626 456
rect 17794 31 22594 456
rect 22762 31 27562 456
rect 27730 31 32530 456
rect 32698 31 37498 456
rect 37666 31 42466 456
rect 42634 31 47434 456
rect 47602 31 52402 456
rect 52570 31 57370 456
rect 57538 31 62338 456
rect 62506 31 67306 456
rect 67474 31 72274 456
rect 72442 31 77242 456
rect 77410 31 82210 456
rect 82378 31 87178 456
rect 87346 31 92146 456
rect 92314 31 97114 456
rect 97282 31 102082 456
rect 102250 31 107050 456
rect 107218 31 112018 456
rect 112186 31 116986 456
rect 117154 31 121954 456
rect 122122 31 126922 456
rect 127090 31 131890 456
rect 132058 31 136858 456
rect 137026 31 141826 456
rect 141994 31 146794 456
rect 146962 31 151762 456
rect 151930 31 156730 456
rect 156898 31 159600 456
<< metal3 >>
rect 159220 76848 159620 76968
rect 159220 70728 159620 70848
rect 159220 64608 159620 64728
rect 159220 58488 159620 58608
rect 159220 52368 159620 52488
rect 159220 46248 159620 46368
rect 0 40128 400 40248
rect 159220 40128 159620 40248
rect 159220 34008 159620 34128
rect 159220 27888 159620 28008
rect 159220 21768 159620 21888
rect 159220 15648 159620 15768
rect 159220 9528 159620 9648
rect 159220 3408 159620 3528
<< obsm3 >>
rect 289 77048 159515 80477
rect 289 76768 159140 77048
rect 289 70928 159515 76768
rect 289 70648 159140 70928
rect 289 64808 159515 70648
rect 289 64528 159140 64808
rect 289 58688 159515 64528
rect 289 58408 159140 58688
rect 289 52568 159515 58408
rect 289 52288 159140 52568
rect 289 46448 159515 52288
rect 289 46168 159140 46448
rect 289 40328 159515 46168
rect 480 40048 159140 40328
rect 289 34208 159515 40048
rect 289 33928 159140 34208
rect 289 28088 159515 33928
rect 289 27808 159140 28088
rect 289 21968 159515 27808
rect 289 21688 159140 21968
rect 289 15848 159515 21688
rect 289 15568 159140 15848
rect 289 9728 159515 15568
rect 289 9448 159140 9728
rect 289 3608 159515 9448
rect 289 3328 159140 3608
rect 289 35 159515 3328
<< metal4 >>
rect 3656 496 3976 80016
rect 19016 496 19336 80016
rect 34376 496 34696 80016
rect 49736 496 50056 80016
rect 65096 496 65416 80016
rect 80456 496 80776 80016
rect 95816 496 96136 80016
rect 111176 496 111496 80016
rect 126536 496 126856 80016
rect 141896 496 142216 80016
rect 157256 496 157576 80016
<< obsm4 >>
rect 1163 80096 157077 80477
rect 1163 851 3576 80096
rect 4056 851 18936 80096
rect 19416 851 34296 80096
rect 34776 851 49656 80096
rect 50136 851 65016 80096
rect 65496 851 80376 80096
rect 80856 851 95736 80096
rect 96216 851 111096 80096
rect 111576 851 126456 80096
rect 126936 851 141816 80096
rect 142296 851 157077 80096
<< labels >>
rlabel metal3 s 159220 34008 159620 34128 6 A0[0]
port 1 nsew signal input
rlabel metal3 s 159220 40128 159620 40248 6 A0[1]
port 2 nsew signal input
rlabel metal3 s 159220 46248 159620 46368 6 A0[2]
port 3 nsew signal input
rlabel metal3 s 159220 52368 159620 52488 6 A0[3]
port 4 nsew signal input
rlabel metal3 s 159220 58488 159620 58608 6 A0[4]
port 5 nsew signal input
rlabel metal3 s 159220 64608 159620 64728 6 A0[5]
port 6 nsew signal input
rlabel metal3 s 159220 70728 159620 70848 6 A0[6]
port 7 nsew signal input
rlabel metal3 s 159220 76848 159620 76968 6 A0[7]
port 8 nsew signal input
rlabel metal3 s 0 40128 400 40248 6 CLK
port 9 nsew signal input
rlabel metal2 s 2778 0 2834 400 6 Di0[0]
port 10 nsew signal input
rlabel metal2 s 52458 0 52514 400 6 Di0[10]
port 11 nsew signal input
rlabel metal2 s 57426 0 57482 400 6 Di0[11]
port 12 nsew signal input
rlabel metal2 s 62394 0 62450 400 6 Di0[12]
port 13 nsew signal input
rlabel metal2 s 67362 0 67418 400 6 Di0[13]
port 14 nsew signal input
rlabel metal2 s 72330 0 72386 400 6 Di0[14]
port 15 nsew signal input
rlabel metal2 s 77298 0 77354 400 6 Di0[15]
port 16 nsew signal input
rlabel metal2 s 82266 0 82322 400 6 Di0[16]
port 17 nsew signal input
rlabel metal2 s 87234 0 87290 400 6 Di0[17]
port 18 nsew signal input
rlabel metal2 s 92202 0 92258 400 6 Di0[18]
port 19 nsew signal input
rlabel metal2 s 97170 0 97226 400 6 Di0[19]
port 20 nsew signal input
rlabel metal2 s 7746 0 7802 400 6 Di0[1]
port 21 nsew signal input
rlabel metal2 s 102138 0 102194 400 6 Di0[20]
port 22 nsew signal input
rlabel metal2 s 107106 0 107162 400 6 Di0[21]
port 23 nsew signal input
rlabel metal2 s 112074 0 112130 400 6 Di0[22]
port 24 nsew signal input
rlabel metal2 s 117042 0 117098 400 6 Di0[23]
port 25 nsew signal input
rlabel metal2 s 122010 0 122066 400 6 Di0[24]
port 26 nsew signal input
rlabel metal2 s 126978 0 127034 400 6 Di0[25]
port 27 nsew signal input
rlabel metal2 s 131946 0 132002 400 6 Di0[26]
port 28 nsew signal input
rlabel metal2 s 136914 0 136970 400 6 Di0[27]
port 29 nsew signal input
rlabel metal2 s 141882 0 141938 400 6 Di0[28]
port 30 nsew signal input
rlabel metal2 s 146850 0 146906 400 6 Di0[29]
port 31 nsew signal input
rlabel metal2 s 12714 0 12770 400 6 Di0[2]
port 32 nsew signal input
rlabel metal2 s 151818 0 151874 400 6 Di0[30]
port 33 nsew signal input
rlabel metal2 s 156786 0 156842 400 6 Di0[31]
port 34 nsew signal input
rlabel metal2 s 17682 0 17738 400 6 Di0[3]
port 35 nsew signal input
rlabel metal2 s 22650 0 22706 400 6 Di0[4]
port 36 nsew signal input
rlabel metal2 s 27618 0 27674 400 6 Di0[5]
port 37 nsew signal input
rlabel metal2 s 32586 0 32642 400 6 Di0[6]
port 38 nsew signal input
rlabel metal2 s 37554 0 37610 400 6 Di0[7]
port 39 nsew signal input
rlabel metal2 s 42522 0 42578 400 6 Di0[8]
port 40 nsew signal input
rlabel metal2 s 47490 0 47546 400 6 Di0[9]
port 41 nsew signal input
rlabel metal2 s 2778 80112 2834 80512 6 Do0[0]
port 42 nsew signal output
rlabel metal2 s 52458 80112 52514 80512 6 Do0[10]
port 43 nsew signal output
rlabel metal2 s 57426 80112 57482 80512 6 Do0[11]
port 44 nsew signal output
rlabel metal2 s 62394 80112 62450 80512 6 Do0[12]
port 45 nsew signal output
rlabel metal2 s 67362 80112 67418 80512 6 Do0[13]
port 46 nsew signal output
rlabel metal2 s 72330 80112 72386 80512 6 Do0[14]
port 47 nsew signal output
rlabel metal2 s 77298 80112 77354 80512 6 Do0[15]
port 48 nsew signal output
rlabel metal2 s 82266 80112 82322 80512 6 Do0[16]
port 49 nsew signal output
rlabel metal2 s 87234 80112 87290 80512 6 Do0[17]
port 50 nsew signal output
rlabel metal2 s 92202 80112 92258 80512 6 Do0[18]
port 51 nsew signal output
rlabel metal2 s 97170 80112 97226 80512 6 Do0[19]
port 52 nsew signal output
rlabel metal2 s 7746 80112 7802 80512 6 Do0[1]
port 53 nsew signal output
rlabel metal2 s 102138 80112 102194 80512 6 Do0[20]
port 54 nsew signal output
rlabel metal2 s 107106 80112 107162 80512 6 Do0[21]
port 55 nsew signal output
rlabel metal2 s 112074 80112 112130 80512 6 Do0[22]
port 56 nsew signal output
rlabel metal2 s 117042 80112 117098 80512 6 Do0[23]
port 57 nsew signal output
rlabel metal2 s 122010 80112 122066 80512 6 Do0[24]
port 58 nsew signal output
rlabel metal2 s 126978 80112 127034 80512 6 Do0[25]
port 59 nsew signal output
rlabel metal2 s 131946 80112 132002 80512 6 Do0[26]
port 60 nsew signal output
rlabel metal2 s 136914 80112 136970 80512 6 Do0[27]
port 61 nsew signal output
rlabel metal2 s 141882 80112 141938 80512 6 Do0[28]
port 62 nsew signal output
rlabel metal2 s 146850 80112 146906 80512 6 Do0[29]
port 63 nsew signal output
rlabel metal2 s 12714 80112 12770 80512 6 Do0[2]
port 64 nsew signal output
rlabel metal2 s 151818 80112 151874 80512 6 Do0[30]
port 65 nsew signal output
rlabel metal2 s 156786 80112 156842 80512 6 Do0[31]
port 66 nsew signal output
rlabel metal2 s 17682 80112 17738 80512 6 Do0[3]
port 67 nsew signal output
rlabel metal2 s 22650 80112 22706 80512 6 Do0[4]
port 68 nsew signal output
rlabel metal2 s 27618 80112 27674 80512 6 Do0[5]
port 69 nsew signal output
rlabel metal2 s 32586 80112 32642 80512 6 Do0[6]
port 70 nsew signal output
rlabel metal2 s 37554 80112 37610 80512 6 Do0[7]
port 71 nsew signal output
rlabel metal2 s 42522 80112 42578 80512 6 Do0[8]
port 72 nsew signal output
rlabel metal2 s 47490 80112 47546 80512 6 Do0[9]
port 73 nsew signal output
rlabel metal3 s 159220 3408 159620 3528 6 EN0
port 74 nsew signal input
rlabel metal4 s 19016 496 19336 80016 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 49736 496 50056 80016 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 80456 496 80776 80016 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 111176 496 111496 80016 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 141896 496 142216 80016 6 VGND
port 75 nsew ground bidirectional
rlabel metal4 s 3656 496 3976 80016 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 34376 496 34696 80016 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 65096 496 65416 80016 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 95816 496 96136 80016 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 126536 496 126856 80016 6 VPWR
port 76 nsew power bidirectional
rlabel metal4 s 157256 496 157576 80016 6 VPWR
port 76 nsew power bidirectional
rlabel metal3 s 159220 9528 159620 9648 6 WE0[0]
port 77 nsew signal input
rlabel metal3 s 159220 15648 159620 15768 6 WE0[1]
port 78 nsew signal input
rlabel metal3 s 159220 21768 159620 21888 6 WE0[2]
port 79 nsew signal input
rlabel metal3 s 159220 27888 159620 28008 6 WE0[3]
port 80 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 159620 80512
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 44017104
string GDS_FILE /mnt/dffram/build/256x32_DEFAULT/openlane/runs/RUN_2022.10.13_02.18.37/results/signoff/RAM256.magic.gds
string GDS_START 183640
<< end >>

