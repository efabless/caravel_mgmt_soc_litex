magic
tech sky130A
magscale 1 2
timestamp 1638229739
<< metal1 >>
rect 277136 160160 277394 160188
rect 144914 160120 144920 160132
rect 141804 160092 144920 160120
rect 63402 160012 63408 160064
rect 63460 160052 63466 160064
rect 141804 160052 141832 160092
rect 144914 160080 144920 160092
rect 144972 160080 144978 160132
rect 63460 160024 141832 160052
rect 63460 160012 63466 160024
rect 141878 160012 141884 160064
rect 141936 160052 141942 160064
rect 154482 160052 154488 160064
rect 141936 160024 154488 160052
rect 141936 160012 141942 160024
rect 154482 160012 154488 160024
rect 154540 160012 154546 160064
rect 156782 160012 156788 160064
rect 156840 160052 156846 160064
rect 191742 160052 191748 160064
rect 156840 160024 191748 160052
rect 156840 160012 156846 160024
rect 191742 160012 191748 160024
rect 191800 160012 191806 160064
rect 197170 160012 197176 160064
rect 197228 160052 197234 160064
rect 207106 160052 207112 160064
rect 197228 160024 207112 160052
rect 197228 160012 197234 160024
rect 207106 160012 207112 160024
rect 207164 160012 207170 160064
rect 211430 160012 211436 160064
rect 211488 160052 211494 160064
rect 277136 160052 277164 160160
rect 211488 160024 277164 160052
rect 277366 160052 277394 160160
rect 330662 160120 330668 160132
rect 327368 160092 330668 160120
rect 280338 160052 280344 160064
rect 277366 160024 280344 160052
rect 211488 160012 211494 160024
rect 280338 160012 280344 160024
rect 280396 160012 280402 160064
rect 281258 160012 281264 160064
rect 281316 160052 281322 160064
rect 327368 160052 327396 160092
rect 330662 160080 330668 160092
rect 330720 160080 330726 160132
rect 336090 160120 336096 160132
rect 335004 160092 336096 160120
rect 281316 160024 327396 160052
rect 281316 160012 281322 160024
rect 327442 160012 327448 160064
rect 327500 160052 327506 160064
rect 333974 160052 333980 160064
rect 327500 160024 333980 160052
rect 327500 160012 327506 160024
rect 333974 160012 333980 160024
rect 334032 160012 334038 160064
rect 334250 160012 334256 160064
rect 334308 160052 334314 160064
rect 335004 160052 335032 160092
rect 336090 160080 336096 160092
rect 336148 160080 336154 160132
rect 338408 160092 339632 160120
rect 334308 160024 335032 160052
rect 334308 160012 334314 160024
rect 335078 160012 335084 160064
rect 335136 160052 335142 160064
rect 338408 160052 338436 160092
rect 335136 160024 338436 160052
rect 335136 160012 335142 160024
rect 338482 160012 338488 160064
rect 338540 160052 338546 160064
rect 339494 160052 339500 160064
rect 338540 160024 339500 160052
rect 338540 160012 338546 160024
rect 339494 160012 339500 160024
rect 339552 160012 339558 160064
rect 339604 160052 339632 160092
rect 374454 160052 374460 160064
rect 339604 160024 374460 160052
rect 374454 160012 374460 160024
rect 374512 160012 374518 160064
rect 378870 160012 378876 160064
rect 378928 160052 378934 160064
rect 398098 160052 398104 160064
rect 378928 160024 398104 160052
rect 378928 160012 378934 160024
rect 398098 160012 398104 160024
rect 398156 160012 398162 160064
rect 455414 160012 455420 160064
rect 455472 160052 455478 160064
rect 466638 160052 466644 160064
rect 455472 160024 466644 160052
rect 455472 160012 455478 160024
rect 466638 160012 466644 160024
rect 466696 160012 466702 160064
rect 468018 160012 468024 160064
rect 468076 160052 468082 160064
rect 476022 160052 476028 160064
rect 468076 160024 476028 160052
rect 468076 160012 468082 160024
rect 476022 160012 476028 160024
rect 476080 160012 476086 160064
rect 25590 159944 25596 159996
rect 25648 159984 25654 159996
rect 109954 159984 109960 159996
rect 25648 159956 109960 159984
rect 25648 159944 25654 159956
rect 109954 159944 109960 159956
rect 110012 159944 110018 159996
rect 117222 159944 117228 159996
rect 117280 159984 117286 159996
rect 191650 159984 191656 159996
rect 117280 159956 191656 159984
rect 117280 159944 117286 159956
rect 191650 159944 191656 159956
rect 191708 159944 191714 159996
rect 197998 159944 198004 159996
rect 198056 159984 198062 159996
rect 269758 159984 269764 159996
rect 198056 159956 269764 159984
rect 198056 159944 198062 159956
rect 269758 159944 269764 159956
rect 269816 159944 269822 159996
rect 271230 159944 271236 159996
rect 271288 159984 271294 159996
rect 272518 159984 272524 159996
rect 271288 159956 272524 159984
rect 271288 159944 271294 159956
rect 272518 159944 272524 159956
rect 272576 159944 272582 159996
rect 275370 159944 275376 159996
rect 275428 159984 275434 159996
rect 328822 159984 328828 159996
rect 275428 159956 328828 159984
rect 275428 159944 275434 159956
rect 328822 159944 328828 159956
rect 328880 159944 328886 159996
rect 329190 159944 329196 159996
rect 329248 159984 329254 159996
rect 370038 159984 370044 159996
rect 329248 159956 370044 159984
rect 329248 159944 329254 159956
rect 370038 159944 370044 159956
rect 370096 159944 370102 159996
rect 372154 159944 372160 159996
rect 372212 159984 372218 159996
rect 396258 159984 396264 159996
rect 372212 159956 396264 159984
rect 372212 159944 372218 159956
rect 396258 159944 396264 159956
rect 396316 159944 396322 159996
rect 403250 159944 403256 159996
rect 403308 159984 403314 159996
rect 416590 159984 416596 159996
rect 403308 159956 416596 159984
rect 403308 159944 403314 159956
rect 416590 159944 416596 159956
rect 416648 159944 416654 159996
rect 467190 159944 467196 159996
rect 467248 159984 467254 159996
rect 473354 159984 473360 159996
rect 467248 159956 473360 159984
rect 467248 159944 467254 159956
rect 473354 159944 473360 159956
rect 473412 159944 473418 159996
rect 76926 159876 76932 159928
rect 76984 159916 76990 159928
rect 162486 159916 162492 159928
rect 76984 159888 162492 159916
rect 76984 159876 76990 159888
rect 162486 159876 162492 159888
rect 162544 159876 162550 159928
rect 166902 159876 166908 159928
rect 166960 159916 166966 159928
rect 186406 159916 186412 159928
rect 166960 159888 186412 159916
rect 166960 159876 166966 159888
rect 186406 159876 186412 159888
rect 186464 159876 186470 159928
rect 191282 159876 191288 159928
rect 191340 159916 191346 159928
rect 264882 159916 264888 159928
rect 191340 159888 264888 159916
rect 191340 159876 191346 159888
rect 264882 159876 264888 159888
rect 264940 159876 264946 159928
rect 268654 159876 268660 159928
rect 268712 159916 268718 159928
rect 323670 159916 323676 159928
rect 268712 159888 323676 159916
rect 268712 159876 268718 159888
rect 323670 159876 323676 159888
rect 323728 159876 323734 159928
rect 328362 159876 328368 159928
rect 328420 159916 328426 159928
rect 369210 159916 369216 159928
rect 328420 159888 369216 159916
rect 328420 159876 328426 159888
rect 369210 159876 369216 159888
rect 369268 159876 369274 159928
rect 373626 159876 373632 159928
rect 373684 159916 373690 159928
rect 379422 159916 379428 159928
rect 373684 159888 379428 159916
rect 373684 159876 373690 159888
rect 379422 159876 379428 159888
rect 379480 159876 379486 159928
rect 379698 159876 379704 159928
rect 379756 159916 379762 159928
rect 405826 159916 405832 159928
rect 379756 159888 405832 159916
rect 379756 159876 379762 159888
rect 405826 159876 405832 159888
rect 405884 159876 405890 159928
rect 409966 159876 409972 159928
rect 410024 159916 410030 159928
rect 417602 159916 417608 159928
rect 410024 159888 417608 159916
rect 410024 159876 410030 159888
rect 417602 159876 417608 159888
rect 417660 159876 417666 159928
rect 480622 159876 480628 159928
rect 480680 159916 480686 159928
rect 485866 159916 485872 159928
rect 480680 159888 485872 159916
rect 480680 159876 480686 159888
rect 485866 159876 485872 159888
rect 485924 159876 485930 159928
rect 70118 159808 70124 159860
rect 70176 159848 70182 159860
rect 156874 159848 156880 159860
rect 70176 159820 156880 159848
rect 70176 159808 70182 159820
rect 156874 159808 156880 159820
rect 156932 159808 156938 159860
rect 166258 159808 166264 159860
rect 166316 159848 166322 159860
rect 172422 159848 172428 159860
rect 166316 159820 172428 159848
rect 166316 159808 166322 159820
rect 172422 159808 172428 159820
rect 172480 159808 172486 159860
rect 180702 159848 180708 159860
rect 175936 159820 180708 159848
rect 56686 159740 56692 159792
rect 56744 159780 56750 159792
rect 137278 159780 137284 159792
rect 56744 159752 137284 159780
rect 56744 159740 56750 159752
rect 137278 159740 137284 159752
rect 137336 159740 137342 159792
rect 137370 159740 137376 159792
rect 137428 159780 137434 159792
rect 139578 159780 139584 159792
rect 137428 159752 139584 159780
rect 137428 159740 137434 159752
rect 139578 159740 139584 159752
rect 139636 159740 139642 159792
rect 139854 159740 139860 159792
rect 139912 159780 139918 159792
rect 144822 159780 144828 159792
rect 139912 159752 144828 159780
rect 139912 159740 139918 159752
rect 144822 159740 144828 159752
rect 144880 159740 144886 159792
rect 144914 159740 144920 159792
rect 144972 159780 144978 159792
rect 146478 159780 146484 159792
rect 144972 159752 146484 159780
rect 144972 159740 144978 159752
rect 146478 159740 146484 159752
rect 146536 159740 146542 159792
rect 146662 159740 146668 159792
rect 146720 159780 146726 159792
rect 153286 159780 153292 159792
rect 146720 159752 153292 159780
rect 146720 159740 146726 159752
rect 153286 159740 153292 159752
rect 153344 159740 153350 159792
rect 153470 159740 153476 159792
rect 153528 159780 153534 159792
rect 175936 159780 175964 159820
rect 180702 159808 180708 159820
rect 180760 159808 180766 159860
rect 184566 159808 184572 159860
rect 184624 159848 184630 159860
rect 259638 159848 259644 159860
rect 184624 159820 259644 159848
rect 184624 159808 184630 159820
rect 259638 159808 259644 159820
rect 259696 159808 259702 159860
rect 261938 159808 261944 159860
rect 261996 159848 262002 159860
rect 318978 159848 318984 159860
rect 261996 159820 318984 159848
rect 261996 159808 262002 159820
rect 318978 159808 318984 159820
rect 319036 159808 319042 159860
rect 320818 159808 320824 159860
rect 320876 159848 320882 159860
rect 356054 159848 356060 159860
rect 320876 159820 356060 159848
rect 320876 159808 320882 159820
rect 356054 159808 356060 159820
rect 356112 159808 356118 159860
rect 359734 159848 359740 159860
rect 356256 159820 359740 159848
rect 153528 159752 175964 159780
rect 153528 159740 153534 159752
rect 177850 159740 177856 159792
rect 177908 159780 177914 159792
rect 254302 159780 254308 159792
rect 177908 159752 254308 159780
rect 177908 159740 177914 159752
rect 254302 159740 254308 159752
rect 254360 159740 254366 159792
rect 255222 159740 255228 159792
rect 255280 159780 255286 159792
rect 313366 159780 313372 159792
rect 255280 159752 313372 159780
rect 255280 159740 255286 159752
rect 313366 159740 313372 159752
rect 313424 159740 313430 159792
rect 314102 159740 314108 159792
rect 314160 159780 314166 159792
rect 355962 159780 355968 159792
rect 314160 159752 355968 159780
rect 314160 159740 314166 159752
rect 355962 159740 355968 159752
rect 356020 159740 356026 159792
rect 18874 159672 18880 159724
rect 18932 159712 18938 159724
rect 109126 159712 109132 159724
rect 18932 159684 109132 159712
rect 18932 159672 18938 159684
rect 109126 159672 109132 159684
rect 109184 159672 109190 159724
rect 113082 159672 113088 159724
rect 113140 159712 113146 159724
rect 126422 159712 126428 159724
rect 113140 159684 126428 159712
rect 113140 159672 113146 159684
rect 126422 159672 126428 159684
rect 126480 159672 126486 159724
rect 126514 159672 126520 159724
rect 126572 159712 126578 159724
rect 156322 159712 156328 159724
rect 126572 159684 156328 159712
rect 126572 159672 126578 159684
rect 156322 159672 156328 159684
rect 156380 159672 156386 159724
rect 164142 159712 164148 159724
rect 156524 159684 164148 159712
rect 49970 159604 49976 159656
rect 50028 159644 50034 159656
rect 143258 159644 143264 159656
rect 50028 159616 143264 159644
rect 50028 159604 50034 159616
rect 143258 159604 143264 159616
rect 143316 159604 143322 159656
rect 143350 159604 143356 159656
rect 143408 159644 143414 159656
rect 156414 159644 156420 159656
rect 143408 159616 156420 159644
rect 143408 159604 143414 159616
rect 156414 159604 156420 159616
rect 156472 159604 156478 159656
rect 43254 159536 43260 159588
rect 43312 159576 43318 159588
rect 137094 159576 137100 159588
rect 43312 159548 137100 159576
rect 43312 159536 43318 159548
rect 137094 159536 137100 159548
rect 137152 159536 137158 159588
rect 137278 159536 137284 159588
rect 137336 159576 137342 159588
rect 139854 159576 139860 159588
rect 137336 159548 139860 159576
rect 137336 159536 137342 159548
rect 139854 159536 139860 159548
rect 139912 159536 139918 159588
rect 139946 159536 139952 159588
rect 140004 159576 140010 159588
rect 156524 159576 156552 159684
rect 164142 159672 164148 159684
rect 164200 159672 164206 159724
rect 167730 159672 167736 159724
rect 167788 159712 167794 159724
rect 246666 159712 246672 159724
rect 167788 159684 246672 159712
rect 167788 159672 167794 159684
rect 246666 159672 246672 159684
rect 246724 159672 246730 159724
rect 250990 159672 250996 159724
rect 251048 159712 251054 159724
rect 310606 159712 310612 159724
rect 251048 159684 310612 159712
rect 251048 159672 251054 159684
rect 310606 159672 310612 159684
rect 310664 159672 310670 159724
rect 315758 159672 315764 159724
rect 315816 159712 315822 159724
rect 356256 159712 356284 159820
rect 359734 159808 359740 159820
rect 359792 159808 359798 159860
rect 376294 159808 376300 159860
rect 376352 159848 376358 159860
rect 405918 159848 405924 159860
rect 376352 159820 405924 159848
rect 376352 159808 376358 159820
rect 405918 159808 405924 159820
rect 405976 159808 405982 159860
rect 449526 159808 449532 159860
rect 449584 159848 449590 159860
rect 459554 159848 459560 159860
rect 449584 159820 459560 159848
rect 449584 159808 449590 159820
rect 459554 159808 459560 159820
rect 459612 159808 459618 159860
rect 461302 159808 461308 159860
rect 461360 159848 461366 159860
rect 468018 159848 468024 159860
rect 461360 159820 468024 159848
rect 461360 159808 461366 159820
rect 468018 159808 468024 159820
rect 468076 159808 468082 159860
rect 478966 159808 478972 159860
rect 479024 159848 479030 159860
rect 484578 159848 484584 159860
rect 479024 159820 484584 159848
rect 479024 159808 479030 159820
rect 484578 159808 484584 159820
rect 484636 159808 484642 159860
rect 357802 159740 357808 159792
rect 357860 159780 357866 159792
rect 365346 159780 365352 159792
rect 357860 159752 365352 159780
rect 357860 159740 357866 159752
rect 365346 159740 365352 159752
rect 365404 159740 365410 159792
rect 365438 159740 365444 159792
rect 365496 159780 365502 159792
rect 395154 159780 395160 159792
rect 365496 159752 395160 159780
rect 365496 159740 365502 159752
rect 395154 159740 395160 159752
rect 395212 159740 395218 159792
rect 396534 159740 396540 159792
rect 396592 159780 396598 159792
rect 413738 159780 413744 159792
rect 396592 159752 413744 159780
rect 396592 159740 396598 159752
rect 413738 159740 413744 159752
rect 413796 159740 413802 159792
rect 420914 159740 420920 159792
rect 420972 159780 420978 159792
rect 440418 159780 440424 159792
rect 420972 159752 440424 159780
rect 420972 159740 420978 159752
rect 440418 159740 440424 159752
rect 440476 159740 440482 159792
rect 453758 159740 453764 159792
rect 453816 159780 453822 159792
rect 464982 159780 464988 159792
rect 453816 159752 464988 159780
rect 453816 159740 453822 159752
rect 464982 159740 464988 159752
rect 465040 159740 465046 159792
rect 471422 159740 471428 159792
rect 471480 159780 471486 159792
rect 478414 159780 478420 159792
rect 471480 159752 478420 159780
rect 471480 159740 471486 159752
rect 478414 159740 478420 159752
rect 478472 159740 478478 159792
rect 315816 159684 356284 159712
rect 315816 159672 315822 159684
rect 369578 159672 369584 159724
rect 369636 159712 369642 159724
rect 400674 159712 400680 159724
rect 369636 159684 400680 159712
rect 369636 159672 369642 159684
rect 400674 159672 400680 159684
rect 400732 159672 400738 159724
rect 407482 159672 407488 159724
rect 407540 159712 407546 159724
rect 429562 159712 429568 159724
rect 407540 159684 429568 159712
rect 407540 159672 407546 159684
rect 429562 159672 429568 159684
rect 429620 159672 429626 159724
rect 450354 159672 450360 159724
rect 450412 159712 450418 159724
rect 462222 159712 462228 159724
rect 450412 159684 462228 159712
rect 450412 159672 450418 159684
rect 462222 159672 462228 159684
rect 462280 159672 462286 159724
rect 468846 159672 468852 159724
rect 468904 159712 468910 159724
rect 474826 159712 474832 159724
rect 468904 159684 474832 159712
rect 468904 159672 468910 159684
rect 474826 159672 474832 159684
rect 474884 159672 474890 159724
rect 156782 159604 156788 159656
rect 156840 159644 156846 159656
rect 160094 159644 160100 159656
rect 156840 159616 160100 159644
rect 156840 159604 156846 159616
rect 160094 159604 160100 159616
rect 160152 159604 160158 159656
rect 161014 159604 161020 159656
rect 161072 159644 161078 159656
rect 241422 159644 241428 159656
rect 161072 159616 241428 159644
rect 161072 159604 161078 159616
rect 241422 159604 241428 159616
rect 241480 159604 241486 159656
rect 244274 159604 244280 159656
rect 244332 159644 244338 159656
rect 297818 159644 297824 159656
rect 244332 159616 297824 159644
rect 244332 159604 244338 159616
rect 297818 159604 297824 159616
rect 297876 159604 297882 159656
rect 303062 159644 303068 159656
rect 297928 159616 303068 159644
rect 140004 159548 156552 159576
rect 140004 159536 140010 159548
rect 157610 159536 157616 159588
rect 157668 159576 157674 159588
rect 238938 159576 238944 159588
rect 157668 159548 238944 159576
rect 157668 159536 157674 159548
rect 238938 159536 238944 159548
rect 238996 159536 239002 159588
rect 241790 159536 241796 159588
rect 241848 159576 241854 159588
rect 297928 159576 297956 159616
rect 303062 159604 303068 159616
rect 303120 159604 303126 159656
rect 309042 159604 309048 159656
rect 309100 159644 309106 159656
rect 354858 159644 354864 159656
rect 309100 159616 354864 159644
rect 309100 159604 309106 159616
rect 354858 159604 354864 159616
rect 354916 159604 354922 159656
rect 356146 159604 356152 159656
rect 356204 159644 356210 159656
rect 359642 159644 359648 159656
rect 356204 159616 359648 159644
rect 356204 159604 356210 159616
rect 359642 159604 359648 159616
rect 359700 159604 359706 159656
rect 362862 159604 362868 159656
rect 362920 159644 362926 159656
rect 395246 159644 395252 159656
rect 362920 159616 395252 159644
rect 362920 159604 362926 159616
rect 395246 159604 395252 159616
rect 395304 159604 395310 159656
rect 399018 159604 399024 159656
rect 399076 159644 399082 159656
rect 408586 159644 408592 159656
rect 399076 159616 408592 159644
rect 399076 159604 399082 159616
rect 408586 159604 408592 159616
rect 408644 159604 408650 159656
rect 410794 159604 410800 159656
rect 410852 159644 410858 159656
rect 432138 159644 432144 159656
rect 410852 159616 432144 159644
rect 410852 159604 410858 159616
rect 432138 159604 432144 159616
rect 432196 159604 432202 159656
rect 451182 159604 451188 159656
rect 451240 159644 451246 159656
rect 461854 159644 461860 159656
rect 451240 159616 461860 159644
rect 451240 159604 451246 159616
rect 461854 159604 461860 159616
rect 461912 159604 461918 159656
rect 476114 159644 476120 159656
rect 470566 159616 476120 159644
rect 470566 159588 470594 159616
rect 476114 159604 476120 159616
rect 476172 159604 476178 159656
rect 482278 159604 482284 159656
rect 482336 159644 482342 159656
rect 487430 159644 487436 159656
rect 482336 159616 487436 159644
rect 482336 159604 482342 159616
rect 487430 159604 487436 159616
rect 487488 159604 487494 159656
rect 241848 159548 297956 159576
rect 241848 159536 241854 159548
rect 302326 159536 302332 159588
rect 302384 159576 302390 159588
rect 347130 159576 347136 159588
rect 302384 159548 347136 159576
rect 302384 159536 302390 159548
rect 347130 159536 347136 159548
rect 347188 159536 347194 159588
rect 347774 159536 347780 159588
rect 347832 159576 347838 159588
rect 347832 159548 349936 159576
rect 347832 159536 347838 159548
rect 36538 159468 36544 159520
rect 36596 159508 36602 159520
rect 126330 159508 126336 159520
rect 36596 159480 126336 159508
rect 36596 159468 36602 159480
rect 126330 159468 126336 159480
rect 126388 159468 126394 159520
rect 126422 159468 126428 159520
rect 126480 159508 126486 159520
rect 127618 159508 127624 159520
rect 126480 159480 127624 159508
rect 126480 159468 126486 159480
rect 127618 159468 127624 159480
rect 127676 159468 127682 159520
rect 129918 159468 129924 159520
rect 129976 159508 129982 159520
rect 141878 159508 141884 159520
rect 129976 159480 141884 159508
rect 129976 159468 129982 159480
rect 141878 159468 141884 159480
rect 141936 159468 141942 159520
rect 144178 159468 144184 159520
rect 144236 159508 144242 159520
rect 225138 159508 225144 159520
rect 144236 159480 225144 159508
rect 144236 159468 144242 159480
rect 225138 159468 225144 159480
rect 225196 159468 225202 159520
rect 231670 159468 231676 159520
rect 231728 159508 231734 159520
rect 295518 159508 295524 159520
rect 231728 159480 295524 159508
rect 231728 159468 231734 159480
rect 295518 159468 295524 159480
rect 295576 159468 295582 159520
rect 295610 159468 295616 159520
rect 295668 159508 295674 159520
rect 335906 159508 335912 159520
rect 295668 159480 335912 159508
rect 295668 159468 295674 159480
rect 335906 159468 335912 159480
rect 335964 159468 335970 159520
rect 336090 159468 336096 159520
rect 336148 159508 336154 159520
rect 339126 159508 339132 159520
rect 336148 159480 339132 159508
rect 336148 159468 336154 159480
rect 339126 159468 339132 159480
rect 339184 159468 339190 159520
rect 339310 159468 339316 159520
rect 339368 159508 339374 159520
rect 349798 159508 349804 159520
rect 339368 159480 349804 159508
rect 339368 159468 339374 159480
rect 349798 159468 349804 159480
rect 349856 159468 349862 159520
rect 349908 159508 349936 159548
rect 351914 159536 351920 159588
rect 351972 159576 351978 159588
rect 385494 159576 385500 159588
rect 351972 159548 385500 159576
rect 351972 159536 351978 159548
rect 385494 159536 385500 159548
rect 385552 159536 385558 159588
rect 389818 159536 389824 159588
rect 389876 159576 389882 159588
rect 413830 159576 413836 159588
rect 389876 159548 413836 159576
rect 389876 159536 389882 159548
rect 413830 159536 413836 159548
rect 413888 159536 413894 159588
rect 414198 159536 414204 159588
rect 414256 159576 414262 159588
rect 434806 159576 434812 159588
rect 414256 159548 434812 159576
rect 414256 159536 414262 159548
rect 434806 159536 434812 159548
rect 434864 159536 434870 159588
rect 452010 159536 452016 159588
rect 452068 159576 452074 159588
rect 463602 159576 463608 159588
rect 452068 159548 463608 159576
rect 452068 159536 452074 159548
rect 463602 159536 463608 159548
rect 463660 159536 463666 159588
rect 470502 159536 470508 159588
rect 470560 159548 470594 159588
rect 470560 159536 470566 159548
rect 472250 159536 472256 159588
rect 472308 159576 472314 159588
rect 479058 159576 479064 159588
rect 472308 159548 479064 159576
rect 472308 159536 472314 159548
rect 479058 159536 479064 159548
rect 479116 159536 479122 159588
rect 479794 159536 479800 159588
rect 479852 159576 479858 159588
rect 484762 159576 484768 159588
rect 479852 159548 484768 159576
rect 479852 159536 479858 159548
rect 484762 159536 484768 159548
rect 484820 159536 484826 159588
rect 359458 159508 359464 159520
rect 349908 159480 359464 159508
rect 359458 159468 359464 159480
rect 359516 159468 359522 159520
rect 392394 159508 392400 159520
rect 359568 159480 392400 159508
rect 32306 159400 32312 159452
rect 32364 159440 32370 159452
rect 32364 159412 123064 159440
rect 32364 159400 32370 159412
rect 6270 159332 6276 159384
rect 6328 159372 6334 159384
rect 122742 159372 122748 159384
rect 6328 159344 122748 159372
rect 6328 159332 6334 159344
rect 122742 159332 122748 159344
rect 122800 159332 122806 159384
rect 123036 159372 123064 159412
rect 123110 159400 123116 159452
rect 123168 159440 123174 159452
rect 147398 159440 147404 159452
rect 123168 159412 147404 159440
rect 123168 159400 123174 159412
rect 147398 159400 147404 159412
rect 147456 159400 147462 159452
rect 150894 159400 150900 159452
rect 150952 159440 150958 159452
rect 233786 159440 233792 159452
rect 150952 159412 233792 159440
rect 150952 159400 150958 159412
rect 233786 159400 233792 159412
rect 233844 159400 233850 159452
rect 234982 159400 234988 159452
rect 235040 159440 235046 159452
rect 298002 159440 298008 159452
rect 235040 159412 298008 159440
rect 235040 159400 235046 159412
rect 298002 159400 298008 159412
rect 298060 159400 298066 159452
rect 301498 159400 301504 159452
rect 301556 159440 301562 159452
rect 348786 159440 348792 159452
rect 301556 159412 348792 159440
rect 301556 159400 301562 159412
rect 348786 159400 348792 159412
rect 348844 159400 348850 159452
rect 348970 159400 348976 159452
rect 349028 159440 349034 159452
rect 353846 159440 353852 159452
rect 349028 159412 353852 159440
rect 349028 159400 349034 159412
rect 353846 159400 353852 159412
rect 353904 159400 353910 159452
rect 355962 159400 355968 159452
rect 356020 159440 356026 159452
rect 357986 159440 357992 159452
rect 356020 159412 357992 159440
rect 356020 159400 356026 159412
rect 357986 159400 357992 159412
rect 358044 159400 358050 159452
rect 358630 159400 358636 159452
rect 358688 159440 358694 159452
rect 359568 159440 359596 159480
rect 392394 159468 392400 159480
rect 392452 159468 392458 159520
rect 424318 159468 424324 159520
rect 424376 159508 424382 159520
rect 442442 159508 442448 159520
rect 424376 159480 442448 159508
rect 424376 159468 424382 159480
rect 442442 159468 442448 159480
rect 442500 159468 442506 159520
rect 446122 159468 446128 159520
rect 446180 159508 446186 159520
rect 456794 159508 456800 159520
rect 446180 159480 456800 159508
rect 446180 159468 446186 159480
rect 456794 159468 456800 159480
rect 456852 159468 456858 159520
rect 458726 159468 458732 159520
rect 458784 159508 458790 159520
rect 465074 159508 465080 159520
rect 458784 159480 465080 159508
rect 458784 159468 458790 159480
rect 465074 159468 465080 159480
rect 465132 159468 465138 159520
rect 469674 159468 469680 159520
rect 469732 159508 469738 159520
rect 477402 159508 477408 159520
rect 469732 159480 477408 159508
rect 469732 159468 469738 159480
rect 477402 159468 477408 159480
rect 477460 159468 477466 159520
rect 478138 159468 478144 159520
rect 478196 159508 478202 159520
rect 483658 159508 483664 159520
rect 478196 159480 483664 159508
rect 478196 159468 478202 159480
rect 483658 159468 483664 159480
rect 483716 159468 483722 159520
rect 518342 159468 518348 159520
rect 518400 159508 518406 159520
rect 522666 159508 522672 159520
rect 518400 159480 522672 159508
rect 518400 159468 518406 159480
rect 522666 159468 522672 159480
rect 522724 159468 522730 159520
rect 358688 159412 359596 159440
rect 358688 159400 358694 159412
rect 359642 159400 359648 159452
rect 359700 159440 359706 159452
rect 390738 159440 390744 159452
rect 359700 159412 390744 159440
rect 359700 159400 359706 159412
rect 390738 159400 390744 159412
rect 390796 159400 390802 159452
rect 400766 159400 400772 159452
rect 400824 159440 400830 159452
rect 424502 159440 424508 159452
rect 400824 159412 424508 159440
rect 400824 159400 400830 159412
rect 424502 159400 424508 159412
rect 424560 159400 424566 159452
rect 427630 159400 427636 159452
rect 427688 159440 427694 159452
rect 445018 159440 445024 159452
rect 427688 159412 445024 159440
rect 427688 159400 427694 159412
rect 445018 159400 445024 159412
rect 445076 159400 445082 159452
rect 447870 159400 447876 159452
rect 447928 159440 447934 159452
rect 460106 159440 460112 159452
rect 447928 159412 460112 159440
rect 447928 159400 447934 159412
rect 460106 159400 460112 159412
rect 460164 159400 460170 159452
rect 462130 159400 462136 159452
rect 462188 159440 462194 159452
rect 467834 159440 467840 159452
rect 462188 159412 467840 159440
rect 462188 159400 462194 159412
rect 467834 159400 467840 159412
rect 467892 159400 467898 159452
rect 477310 159400 477316 159452
rect 477368 159440 477374 159452
rect 483290 159440 483296 159452
rect 477368 159412 483296 159440
rect 477368 159400 477374 159412
rect 483290 159400 483296 159412
rect 483348 159400 483354 159452
rect 126882 159372 126888 159384
rect 123036 159344 126888 159372
rect 126882 159332 126888 159344
rect 126940 159332 126946 159384
rect 126974 159332 126980 159384
rect 127032 159372 127038 159384
rect 130654 159372 130660 159384
rect 127032 159344 130660 159372
rect 127032 159332 127038 159344
rect 130654 159332 130660 159344
rect 130712 159332 130718 159384
rect 133138 159332 133144 159384
rect 133196 159372 133202 159384
rect 137370 159372 137376 159384
rect 133196 159344 137376 159372
rect 133196 159332 133202 159344
rect 137370 159332 137376 159344
rect 137428 159332 137434 159384
rect 137462 159332 137468 159384
rect 137520 159372 137526 159384
rect 223574 159372 223580 159384
rect 137520 159344 223580 159372
rect 137520 159332 137526 159344
rect 223574 159332 223580 159344
rect 223632 159332 223638 159384
rect 224954 159332 224960 159384
rect 225012 159372 225018 159384
rect 290274 159372 290280 159384
rect 225012 159344 290280 159372
rect 225012 159332 225018 159344
rect 290274 159332 290280 159344
rect 290332 159332 290338 159384
rect 294782 159332 294788 159384
rect 294840 159372 294846 159384
rect 343450 159372 343456 159384
rect 294840 159344 343456 159372
rect 294840 159332 294846 159344
rect 343450 159332 343456 159344
rect 343508 159332 343514 159384
rect 346026 159332 346032 159384
rect 346084 159372 346090 159384
rect 346084 159344 374684 159372
rect 346084 159332 346090 159344
rect 73522 159264 73528 159316
rect 73580 159304 73586 159316
rect 80054 159304 80060 159316
rect 73580 159276 80060 159304
rect 73580 159264 73586 159276
rect 80054 159264 80060 159276
rect 80112 159264 80118 159316
rect 83642 159264 83648 159316
rect 83700 159304 83706 159316
rect 166994 159304 167000 159316
rect 83700 159276 167000 159304
rect 83700 159264 83706 159276
rect 166994 159264 167000 159276
rect 167052 159264 167058 159316
rect 170214 159264 170220 159316
rect 170272 159304 170278 159316
rect 199286 159304 199292 159316
rect 170272 159276 199292 159304
rect 170272 159264 170278 159276
rect 199286 159264 199292 159276
rect 199344 159264 199350 159316
rect 201402 159264 201408 159316
rect 201460 159304 201466 159316
rect 213086 159304 213092 159316
rect 201460 159276 213092 159304
rect 201460 159264 201466 159276
rect 213086 159264 213092 159276
rect 213144 159264 213150 159316
rect 214006 159264 214012 159316
rect 214064 159304 214070 159316
rect 281994 159304 282000 159316
rect 214064 159276 282000 159304
rect 214064 159264 214070 159276
rect 281994 159264 282000 159276
rect 282052 159264 282058 159316
rect 282086 159264 282092 159316
rect 282144 159304 282150 159316
rect 327442 159304 327448 159316
rect 282144 159276 327448 159304
rect 282144 159264 282150 159276
rect 327442 159264 327448 159276
rect 327500 159264 327506 159316
rect 327534 159264 327540 159316
rect 327592 159304 327598 159316
rect 330570 159304 330576 159316
rect 327592 159276 330576 159304
rect 327592 159264 327598 159276
rect 330570 159264 330576 159276
rect 330628 159264 330634 159316
rect 330662 159264 330668 159316
rect 330720 159304 330726 159316
rect 333330 159304 333336 159316
rect 330720 159276 333336 159304
rect 330720 159264 330726 159276
rect 333330 159264 333336 159276
rect 333388 159264 333394 159316
rect 333514 159264 333520 159316
rect 333572 159304 333578 159316
rect 339034 159304 339040 159316
rect 333572 159276 339040 159304
rect 333572 159264 333578 159276
rect 339034 159264 339040 159276
rect 339092 159264 339098 159316
rect 339126 159264 339132 159316
rect 339184 159304 339190 159316
rect 374086 159304 374092 159316
rect 339184 159276 374092 159304
rect 339184 159264 339190 159276
rect 374086 159264 374092 159276
rect 374144 159264 374150 159316
rect 80238 159196 80244 159248
rect 80296 159236 80302 159248
rect 91094 159236 91100 159248
rect 80296 159208 91100 159236
rect 80296 159196 80302 159208
rect 91094 159196 91100 159208
rect 91152 159196 91158 159248
rect 100478 159196 100484 159248
rect 100536 159236 100542 159248
rect 184658 159236 184664 159248
rect 100536 159208 184664 159236
rect 100536 159196 100542 159208
rect 184658 159196 184664 159208
rect 184716 159196 184722 159248
rect 187050 159196 187056 159248
rect 187108 159236 187114 159248
rect 214098 159236 214104 159248
rect 187108 159208 214104 159236
rect 187108 159196 187114 159208
rect 214098 159196 214104 159208
rect 214156 159196 214162 159248
rect 218238 159196 218244 159248
rect 218296 159236 218302 159248
rect 285122 159236 285128 159248
rect 218296 159208 285128 159236
rect 218296 159196 218302 159208
rect 285122 159196 285128 159208
rect 285180 159196 285186 159248
rect 287974 159196 287980 159248
rect 288032 159236 288038 159248
rect 288032 159208 335124 159236
rect 288032 159196 288038 159208
rect 86954 159128 86960 159180
rect 87012 159168 87018 159180
rect 169938 159168 169944 159180
rect 87012 159140 169944 159168
rect 87012 159128 87018 159140
rect 169938 159128 169944 159140
rect 169996 159128 170002 159180
rect 171134 159128 171140 159180
rect 171192 159168 171198 159180
rect 172514 159168 172520 159180
rect 171192 159140 172520 159168
rect 171192 159128 171198 159140
rect 172514 159128 172520 159140
rect 172572 159128 172578 159180
rect 173618 159128 173624 159180
rect 173676 159168 173682 159180
rect 197354 159168 197360 159180
rect 173676 159140 197360 159168
rect 173676 159128 173682 159140
rect 197354 159128 197360 159140
rect 197412 159128 197418 159180
rect 203886 159128 203892 159180
rect 203944 159168 203950 159180
rect 213638 159168 213644 159180
rect 203944 159140 213644 159168
rect 203944 159128 203950 159140
rect 213638 159128 213644 159140
rect 213696 159128 213702 159180
rect 220722 159128 220728 159180
rect 220780 159168 220786 159180
rect 283006 159168 283012 159180
rect 220780 159140 283012 159168
rect 220780 159128 220786 159140
rect 283006 159128 283012 159140
rect 283064 159128 283070 159180
rect 284662 159128 284668 159180
rect 284720 159168 284726 159180
rect 285766 159168 285772 159180
rect 284720 159140 285772 159168
rect 284720 159128 284726 159140
rect 285766 159128 285772 159140
rect 285824 159128 285830 159180
rect 288342 159168 288348 159180
rect 287026 159140 288348 159168
rect 93670 159060 93676 159112
rect 93728 159100 93734 159112
rect 166258 159100 166264 159112
rect 93728 159072 166264 159100
rect 93728 159060 93734 159072
rect 166258 159060 166264 159072
rect 166316 159060 166322 159112
rect 183462 159100 183468 159112
rect 171106 159072 183468 159100
rect 107194 158992 107200 159044
rect 107252 159032 107258 159044
rect 171106 159032 171134 159072
rect 183462 159060 183468 159072
rect 183520 159060 183526 159112
rect 193766 159060 193772 159112
rect 193824 159100 193830 159112
rect 218054 159100 218060 159112
rect 193824 159072 218060 159100
rect 193824 159060 193830 159072
rect 218054 159060 218060 159072
rect 218112 159060 218118 159112
rect 224126 159060 224132 159112
rect 224184 159100 224190 159112
rect 287026 159100 287054 159140
rect 288342 159128 288348 159140
rect 288400 159128 288406 159180
rect 288894 159128 288900 159180
rect 288952 159168 288958 159180
rect 333514 159168 333520 159180
rect 288952 159140 333520 159168
rect 288952 159128 288958 159140
rect 333514 159128 333520 159140
rect 333572 159128 333578 159180
rect 335096 159168 335124 159208
rect 335906 159196 335912 159248
rect 335964 159236 335970 159248
rect 342438 159236 342444 159248
rect 335964 159208 342444 159236
rect 335964 159196 335970 159208
rect 342438 159196 342444 159208
rect 342496 159196 342502 159248
rect 342714 159196 342720 159248
rect 342772 159236 342778 159248
rect 343818 159236 343824 159248
rect 342772 159208 343824 159236
rect 342772 159196 342778 159208
rect 343818 159196 343824 159208
rect 343876 159196 343882 159248
rect 347130 159196 347136 159248
rect 347188 159236 347194 159248
rect 349338 159236 349344 159248
rect 347188 159208 349344 159236
rect 347188 159196 347194 159208
rect 349338 159196 349344 159208
rect 349396 159196 349402 159248
rect 349798 159196 349804 159248
rect 349856 159236 349862 159248
rect 374656 159236 374684 159344
rect 374730 159332 374736 159384
rect 374788 159372 374794 159384
rect 385862 159372 385868 159384
rect 374788 159344 385868 159372
rect 374788 159332 374794 159344
rect 385862 159332 385868 159344
rect 385920 159332 385926 159384
rect 388990 159332 388996 159384
rect 389048 159372 389054 159384
rect 403894 159372 403900 159384
rect 389048 159344 403900 159372
rect 389048 159332 389054 159344
rect 403894 159332 403900 159344
rect 403952 159332 403958 159384
rect 417510 159332 417516 159384
rect 417568 159372 417574 159384
rect 437658 159372 437664 159384
rect 417568 159344 437664 159372
rect 417568 159332 417574 159344
rect 437658 159332 437664 159344
rect 437716 159332 437722 159384
rect 448698 159332 448704 159384
rect 448756 159372 448762 159384
rect 461118 159372 461124 159384
rect 448756 159344 461124 159372
rect 448756 159332 448762 159344
rect 461118 159332 461124 159344
rect 461176 159332 461182 159384
rect 463786 159332 463792 159384
rect 463844 159372 463850 159384
rect 471698 159372 471704 159384
rect 463844 159344 471704 159372
rect 463844 159332 463850 159344
rect 471698 159332 471704 159344
rect 471756 159332 471762 159384
rect 518710 159332 518716 159384
rect 518768 159372 518774 159384
rect 523494 159372 523500 159384
rect 518768 159344 523500 159372
rect 518768 159332 518774 159344
rect 523494 159332 523500 159344
rect 523552 159332 523558 159384
rect 378042 159264 378048 159316
rect 378100 159304 378106 159316
rect 388346 159304 388352 159316
rect 378100 159276 388352 159304
rect 378100 159264 378106 159276
rect 388346 159264 388352 159276
rect 388404 159264 388410 159316
rect 404078 159264 404084 159316
rect 404136 159304 404142 159316
rect 426986 159304 426992 159316
rect 404136 159276 426992 159304
rect 404136 159264 404142 159276
rect 426986 159264 426992 159276
rect 427044 159264 427050 159316
rect 454586 159264 454592 159316
rect 454644 159304 454650 159316
rect 465442 159304 465448 159316
rect 454644 159276 465448 159304
rect 454644 159264 454650 159276
rect 465442 159264 465448 159276
rect 465500 159264 465506 159316
rect 465534 159264 465540 159316
rect 465592 159304 465598 159316
rect 472250 159304 472256 159316
rect 465592 159276 472256 159304
rect 465592 159264 465598 159276
rect 472250 159264 472256 159276
rect 472308 159264 472314 159316
rect 382734 159236 382740 159248
rect 349856 159208 373764 159236
rect 374656 159208 382740 159236
rect 349856 159196 349862 159208
rect 338390 159168 338396 159180
rect 335096 159140 338396 159168
rect 338390 159128 338396 159140
rect 338448 159128 338454 159180
rect 341886 159128 341892 159180
rect 341944 159168 341950 159180
rect 373626 159168 373632 159180
rect 341944 159140 373632 159168
rect 341944 159128 341950 159140
rect 373626 159128 373632 159140
rect 373684 159128 373690 159180
rect 373736 159168 373764 159208
rect 382734 159196 382740 159208
rect 382792 159196 382798 159248
rect 385586 159196 385592 159248
rect 385644 159236 385650 159248
rect 399570 159236 399576 159248
rect 385644 159208 399576 159236
rect 385644 159196 385650 159208
rect 399570 159196 399576 159208
rect 399628 159196 399634 159248
rect 457898 159196 457904 159248
rect 457956 159236 457962 159248
rect 468110 159236 468116 159248
rect 457956 159208 468116 159236
rect 457956 159196 457962 159208
rect 468110 159196 468116 159208
rect 468168 159196 468174 159248
rect 377582 159168 377588 159180
rect 373736 159140 377588 159168
rect 377582 159128 377588 159140
rect 377640 159128 377646 159180
rect 392302 159128 392308 159180
rect 392360 159168 392366 159180
rect 404262 159168 404268 159180
rect 392360 159140 404268 159168
rect 392360 159128 392366 159140
rect 404262 159128 404268 159140
rect 404320 159128 404326 159180
rect 457070 159128 457076 159180
rect 457128 159168 457134 159180
rect 467926 159168 467932 159180
rect 457128 159140 467932 159168
rect 457128 159128 457134 159140
rect 467926 159128 467932 159140
rect 467984 159128 467990 159180
rect 224184 159072 287054 159100
rect 224184 159060 224190 159072
rect 297818 159060 297824 159112
rect 297876 159100 297882 159112
rect 305178 159100 305184 159112
rect 297876 159072 305184 159100
rect 297876 159060 297882 159072
rect 305178 159060 305184 159072
rect 305236 159060 305242 159112
rect 307386 159060 307392 159112
rect 307444 159100 307450 159112
rect 307444 159072 349200 159100
rect 307444 159060 307450 159072
rect 107252 159004 171134 159032
rect 107252 158992 107258 159004
rect 174354 158992 174360 159044
rect 174412 159032 174418 159044
rect 176654 159032 176660 159044
rect 174412 159004 176660 159032
rect 174412 158992 174418 159004
rect 176654 158992 176660 159004
rect 176712 158992 176718 159044
rect 183738 158992 183744 159044
rect 183796 159032 183802 159044
rect 200482 159032 200488 159044
rect 183796 159004 200488 159032
rect 183796 158992 183802 159004
rect 200482 158992 200488 159004
rect 200540 158992 200546 159044
rect 200574 158992 200580 159044
rect 200632 159032 200638 159044
rect 224954 159032 224960 159044
rect 200632 159004 224960 159032
rect 200632 158992 200638 159004
rect 224954 158992 224960 159004
rect 225012 158992 225018 159044
rect 230842 158992 230848 159044
rect 230900 159032 230906 159044
rect 294782 159032 294788 159044
rect 230900 159004 294788 159032
rect 230900 158992 230906 159004
rect 294782 158992 294788 159004
rect 294840 158992 294846 159044
rect 298094 158992 298100 159044
rect 298152 159032 298158 159044
rect 299934 159032 299940 159044
rect 298152 159004 299940 159032
rect 298152 158992 298158 159004
rect 299934 158992 299940 159004
rect 299992 158992 299998 159044
rect 308214 158992 308220 159044
rect 308272 159032 308278 159044
rect 348970 159032 348976 159044
rect 308272 159004 348976 159032
rect 308272 158992 308278 159004
rect 348970 158992 348976 159004
rect 349028 158992 349034 159044
rect 349172 159032 349200 159072
rect 351086 159060 351092 159112
rect 351144 159100 351150 159112
rect 382366 159100 382372 159112
rect 351144 159072 382372 159100
rect 351144 159060 351150 159072
rect 382366 159060 382372 159072
rect 382424 159060 382430 159112
rect 395706 159060 395712 159112
rect 395764 159100 395770 159112
rect 405642 159100 405648 159112
rect 395764 159072 405648 159100
rect 395764 159060 395770 159072
rect 405642 159060 405648 159072
rect 405700 159060 405706 159112
rect 412542 159060 412548 159112
rect 412600 159100 412606 159112
rect 413922 159100 413928 159112
rect 412600 159072 413928 159100
rect 412600 159060 412606 159072
rect 413922 159060 413928 159072
rect 413980 159060 413986 159112
rect 459646 159060 459652 159112
rect 459704 159100 459710 159112
rect 466454 159100 466460 159112
rect 459704 159072 466460 159100
rect 459704 159060 459710 159072
rect 466454 159060 466460 159072
rect 466512 159060 466518 159112
rect 353202 159032 353208 159044
rect 349172 159004 353208 159032
rect 353202 158992 353208 159004
rect 353260 158992 353266 159044
rect 356054 158992 356060 159044
rect 356112 159032 356118 159044
rect 356112 159004 358860 159032
rect 356112 158992 356118 159004
rect 96246 158924 96252 158976
rect 96304 158964 96310 158976
rect 121638 158964 121644 158976
rect 96304 158936 121644 158964
rect 96304 158924 96310 158936
rect 121638 158924 121644 158936
rect 121696 158924 121702 158976
rect 124030 158924 124036 158976
rect 124088 158964 124094 158976
rect 194502 158964 194508 158976
rect 124088 158936 194508 158964
rect 124088 158924 124094 158936
rect 194502 158924 194508 158936
rect 194560 158924 194566 158976
rect 194686 158924 194692 158976
rect 194744 158964 194750 158976
rect 203702 158964 203708 158976
rect 194744 158936 203708 158964
rect 194744 158924 194750 158936
rect 203702 158924 203708 158936
rect 203760 158924 203766 158976
rect 208118 158924 208124 158976
rect 208176 158964 208182 158976
rect 212442 158964 212448 158976
rect 208176 158936 212448 158964
rect 208176 158924 208182 158936
rect 212442 158924 212448 158936
rect 212500 158924 212506 158976
rect 231026 158964 231032 158976
rect 214576 158936 231032 158964
rect 125502 158896 125508 158908
rect 103486 158868 125508 158896
rect 102962 158788 102968 158840
rect 103020 158828 103026 158840
rect 103486 158828 103514 158868
rect 125502 158856 125508 158868
rect 125560 158856 125566 158908
rect 127342 158856 127348 158908
rect 127400 158896 127406 158908
rect 127986 158896 127992 158908
rect 127400 158868 127992 158896
rect 127400 158856 127406 158868
rect 127986 158856 127992 158868
rect 128044 158856 128050 158908
rect 130746 158856 130752 158908
rect 130804 158896 130810 158908
rect 194962 158896 194968 158908
rect 130804 158868 194968 158896
rect 130804 158856 130810 158868
rect 194962 158856 194968 158868
rect 195020 158856 195026 158908
rect 113818 158828 113824 158840
rect 103020 158800 103514 158828
rect 108316 158800 113824 158828
rect 103020 158788 103026 158800
rect 90358 158720 90364 158772
rect 90416 158760 90422 158772
rect 92474 158760 92480 158772
rect 90416 158732 92480 158760
rect 90416 158720 90422 158732
rect 92474 158720 92480 158732
rect 92532 158720 92538 158772
rect 92842 158720 92848 158772
rect 92900 158760 92906 158772
rect 108316 158760 108344 158800
rect 113818 158788 113824 158800
rect 113876 158788 113882 158840
rect 133138 158828 133144 158840
rect 117976 158800 133144 158828
rect 92900 158732 108344 158760
rect 92900 158720 92906 158732
rect 109678 158720 109684 158772
rect 109736 158760 109742 158772
rect 117976 158760 118004 158800
rect 133138 158788 133144 158800
rect 133196 158788 133202 158840
rect 133230 158788 133236 158840
rect 133288 158828 133294 158840
rect 158714 158828 158720 158840
rect 133288 158800 158720 158828
rect 133288 158788 133294 158800
rect 158714 158788 158720 158800
rect 158772 158788 158778 158840
rect 163498 158788 163504 158840
rect 163556 158828 163562 158840
rect 196066 158828 196072 158840
rect 163556 158800 196072 158828
rect 163556 158788 163562 158800
rect 196066 158788 196072 158800
rect 196124 158788 196130 158840
rect 207290 158788 207296 158840
rect 207348 158828 207354 158840
rect 214576 158828 214604 158936
rect 231026 158924 231032 158936
rect 231084 158924 231090 158976
rect 237558 158924 237564 158976
rect 237616 158964 237622 158976
rect 300026 158964 300032 158976
rect 237616 158936 300032 158964
rect 237616 158924 237622 158936
rect 300026 158924 300032 158936
rect 300084 158924 300090 158976
rect 301516 158936 308260 158964
rect 217318 158856 217324 158908
rect 217376 158896 217382 158908
rect 220722 158896 220728 158908
rect 217376 158868 220728 158896
rect 217376 158856 217382 158868
rect 220722 158856 220728 158868
rect 220780 158856 220786 158908
rect 248506 158856 248512 158908
rect 248564 158896 248570 158908
rect 301516 158896 301544 158936
rect 308232 158908 308260 158936
rect 314930 158924 314936 158976
rect 314988 158964 314994 158976
rect 358722 158964 358728 158976
rect 314988 158936 358728 158964
rect 314988 158924 314994 158936
rect 358722 158924 358728 158936
rect 358780 158924 358786 158976
rect 358832 158964 358860 159004
rect 359458 158992 359464 159044
rect 359516 159032 359522 159044
rect 378778 159032 378784 159044
rect 359516 159004 378784 159032
rect 359516 158992 359522 159004
rect 378778 158992 378784 159004
rect 378836 158992 378842 159044
rect 383102 158992 383108 159044
rect 383160 159032 383166 159044
rect 411438 159032 411444 159044
rect 383160 159004 411444 159032
rect 383160 158992 383166 159004
rect 411438 158992 411444 159004
rect 411496 158992 411502 159044
rect 462958 158992 462964 159044
rect 463016 159032 463022 159044
rect 469214 159032 469220 159044
rect 463016 159004 469220 159032
rect 463016 158992 463022 159004
rect 469214 158992 469220 159004
rect 469272 158992 469278 159044
rect 473906 158992 473912 159044
rect 473964 159032 473970 159044
rect 480254 159032 480260 159044
rect 473964 159004 480260 159032
rect 473964 158992 473970 159004
rect 480254 158992 480260 159004
rect 480312 158992 480318 159044
rect 363506 158964 363512 158976
rect 358832 158936 363512 158964
rect 363506 158924 363512 158936
rect 363564 158924 363570 158976
rect 364794 158964 364800 158976
rect 364306 158936 364800 158964
rect 248564 158868 301544 158896
rect 248564 158856 248570 158868
rect 305638 158856 305644 158908
rect 305696 158896 305702 158908
rect 307662 158896 307668 158908
rect 305696 158868 307668 158896
rect 305696 158856 305702 158868
rect 307662 158856 307668 158868
rect 307720 158856 307726 158908
rect 308214 158856 308220 158908
rect 308272 158856 308278 158908
rect 310698 158856 310704 158908
rect 310756 158896 310762 158908
rect 311986 158896 311992 158908
rect 310756 158868 311992 158896
rect 310756 158856 310762 158868
rect 311986 158856 311992 158868
rect 312044 158856 312050 158908
rect 312446 158856 312452 158908
rect 312504 158896 312510 158908
rect 313458 158896 313464 158908
rect 312504 158868 313464 158896
rect 312504 158856 312510 158868
rect 313458 158856 313464 158868
rect 313516 158856 313522 158908
rect 319162 158856 319168 158908
rect 319220 158896 319226 158908
rect 322842 158896 322848 158908
rect 319220 158868 322848 158896
rect 319220 158856 319226 158868
rect 322842 158856 322848 158868
rect 322900 158856 322906 158908
rect 364306 158896 364334 158936
rect 364794 158924 364800 158936
rect 364852 158924 364858 158976
rect 365346 158924 365352 158976
rect 365404 158964 365410 158976
rect 371878 158964 371884 158976
rect 365404 158936 371884 158964
rect 365404 158924 365410 158936
rect 371878 158924 371884 158936
rect 371936 158924 371942 158976
rect 374546 158924 374552 158976
rect 374604 158964 374610 158976
rect 386322 158964 386328 158976
rect 374604 158936 386328 158964
rect 374604 158924 374610 158936
rect 386322 158924 386328 158936
rect 386380 158924 386386 158976
rect 391474 158924 391480 158976
rect 391532 158964 391538 158976
rect 394602 158964 394608 158976
rect 391532 158936 394608 158964
rect 391532 158924 391538 158936
rect 394602 158924 394608 158936
rect 394660 158924 394666 158976
rect 409138 158924 409144 158976
rect 409196 158964 409202 158976
rect 410886 158964 410892 158976
rect 409196 158936 410892 158964
rect 409196 158924 409202 158936
rect 410886 158924 410892 158936
rect 410944 158924 410950 158976
rect 420086 158924 420092 158976
rect 420144 158964 420150 158976
rect 423582 158964 423588 158976
rect 420144 158936 423588 158964
rect 420144 158924 420150 158936
rect 423582 158924 423588 158936
rect 423640 158924 423646 158976
rect 460474 158924 460480 158976
rect 460532 158964 460538 158976
rect 466546 158964 466552 158976
rect 460532 158936 466552 158964
rect 460532 158924 460538 158936
rect 466546 158924 466552 158936
rect 466604 158924 466610 158976
rect 475562 158924 475568 158976
rect 475620 158964 475626 158976
rect 481726 158964 481732 158976
rect 475620 158936 481732 158964
rect 475620 158924 475626 158936
rect 481726 158924 481732 158936
rect 481784 158924 481790 158976
rect 329668 158868 364334 158896
rect 374564 158868 379514 158896
rect 207348 158800 214604 158828
rect 207348 158788 207354 158800
rect 214834 158788 214840 158840
rect 214892 158828 214898 158840
rect 221734 158828 221740 158840
rect 214892 158800 221740 158828
rect 214892 158788 214898 158800
rect 221734 158788 221740 158800
rect 221792 158788 221798 158840
rect 238386 158788 238392 158840
rect 238444 158828 238450 158840
rect 242802 158828 242808 158840
rect 238444 158800 242808 158828
rect 238444 158788 238450 158800
rect 242802 158788 242808 158800
rect 242860 158788 242866 158840
rect 261110 158788 261116 158840
rect 261168 158828 261174 158840
rect 316954 158828 316960 158840
rect 261168 158800 316960 158828
rect 261168 158788 261174 158800
rect 316954 158788 316960 158800
rect 317012 158788 317018 158840
rect 322474 158788 322480 158840
rect 322532 158828 322538 158840
rect 329668 158828 329696 158868
rect 361114 158828 361120 158840
rect 322532 158800 329696 158828
rect 330496 158800 361120 158828
rect 322532 158788 322538 158800
rect 109736 158732 118004 158760
rect 109736 158720 109742 158732
rect 118970 158720 118976 158772
rect 119028 158760 119034 158772
rect 119614 158760 119620 158772
rect 119028 158732 119620 158760
rect 119028 158720 119034 158732
rect 119614 158720 119620 158732
rect 119672 158720 119678 158772
rect 119798 158720 119804 158772
rect 119856 158760 119862 158772
rect 147398 158760 147404 158772
rect 119856 158732 147404 158760
rect 119856 158720 119862 158732
rect 147398 158720 147404 158732
rect 147456 158720 147462 158772
rect 147490 158720 147496 158772
rect 147548 158760 147554 158772
rect 149054 158760 149060 158772
rect 147548 158732 149060 158760
rect 147548 158720 147554 158732
rect 149054 158720 149060 158732
rect 149112 158720 149118 158772
rect 153286 158720 153292 158772
rect 153344 158760 153350 158772
rect 174354 158760 174360 158772
rect 153344 158732 174360 158760
rect 153344 158720 153350 158732
rect 174354 158720 174360 158732
rect 174412 158720 174418 158772
rect 174446 158720 174452 158772
rect 174504 158760 174510 158772
rect 174906 158760 174912 158772
rect 174504 158732 174912 158760
rect 174504 158720 174510 158732
rect 174906 158720 174912 158732
rect 174964 158720 174970 158772
rect 180334 158720 180340 158772
rect 180392 158760 180398 158772
rect 204898 158760 204904 158772
rect 180392 158732 204904 158760
rect 180392 158720 180398 158732
rect 204898 158720 204904 158732
rect 204956 158720 204962 158772
rect 210602 158720 210608 158772
rect 210660 158760 210666 158772
rect 215294 158760 215300 158772
rect 210660 158732 215300 158760
rect 210660 158720 210666 158732
rect 215294 158720 215300 158732
rect 215352 158720 215358 158772
rect 221550 158720 221556 158772
rect 221608 158760 221614 158772
rect 223850 158760 223856 158772
rect 221608 158732 223856 158760
rect 221608 158720 221614 158732
rect 223850 158720 223856 158732
rect 223908 158720 223914 158772
rect 240870 158720 240876 158772
rect 240928 158760 240934 158772
rect 243354 158760 243360 158772
rect 240928 158732 243360 158760
rect 240928 158720 240934 158732
rect 243354 158720 243360 158732
rect 243412 158720 243418 158772
rect 254394 158720 254400 158772
rect 254452 158760 254458 158772
rect 255314 158760 255320 158772
rect 254452 158732 255320 158760
rect 254452 158720 254458 158732
rect 255314 158720 255320 158732
rect 255372 158720 255378 158772
rect 258534 158720 258540 158772
rect 258592 158760 258598 158772
rect 260926 158760 260932 158772
rect 258592 158732 260932 158760
rect 258592 158720 258598 158732
rect 260926 158720 260932 158732
rect 260984 158720 260990 158772
rect 264422 158720 264428 158772
rect 264480 158760 264486 158772
rect 267090 158760 267096 158772
rect 264480 158732 267096 158760
rect 264480 158720 264486 158732
rect 267090 158720 267096 158732
rect 267148 158720 267154 158772
rect 267826 158720 267832 158772
rect 267884 158760 267890 158772
rect 320266 158760 320272 158772
rect 267884 158732 320272 158760
rect 267884 158720 267890 158732
rect 320266 158720 320272 158732
rect 320324 158720 320330 158772
rect 321646 158720 321652 158772
rect 321704 158760 321710 158772
rect 330496 158760 330524 158800
rect 361114 158788 361120 158800
rect 361172 158788 361178 158840
rect 361206 158788 361212 158840
rect 361264 158828 361270 158840
rect 361264 158800 367876 158828
rect 361264 158788 361270 158800
rect 321704 158732 330524 158760
rect 321704 158720 321710 158732
rect 330570 158720 330576 158772
rect 330628 158760 330634 158772
rect 367186 158760 367192 158772
rect 330628 158732 367192 158760
rect 330628 158720 330634 158732
rect 367186 158720 367192 158732
rect 367244 158720 367250 158772
rect 81066 158652 81072 158704
rect 81124 158692 81130 158704
rect 180794 158692 180800 158704
rect 81124 158664 180800 158692
rect 81124 158652 81130 158664
rect 180794 158652 180800 158664
rect 180852 158652 180858 158704
rect 180886 158652 180892 158704
rect 180944 158692 180950 158704
rect 181898 158692 181904 158704
rect 180944 158664 181904 158692
rect 180944 158652 180950 158664
rect 181898 158652 181904 158664
rect 181956 158652 181962 158704
rect 181990 158652 181996 158704
rect 182048 158692 182054 158704
rect 257522 158692 257528 158704
rect 182048 158664 257528 158692
rect 182048 158652 182054 158664
rect 257522 158652 257528 158664
rect 257580 158652 257586 158704
rect 367848 158692 367876 158800
rect 371878 158788 371884 158840
rect 371936 158828 371942 158840
rect 374564 158828 374592 158868
rect 371936 158800 374592 158828
rect 371936 158788 371942 158800
rect 374822 158788 374828 158840
rect 374880 158828 374886 158840
rect 379486 158828 379514 158868
rect 384758 158856 384764 158908
rect 384816 158896 384822 158908
rect 389174 158896 389180 158908
rect 384816 158868 389180 158896
rect 384816 158856 384822 158868
rect 389174 158856 389180 158868
rect 389232 158856 389238 158908
rect 405734 158856 405740 158908
rect 405792 158896 405798 158908
rect 409322 158896 409328 158908
rect 405792 158868 409328 158896
rect 405792 158856 405798 158868
rect 409322 158856 409328 158868
rect 409380 158856 409386 158908
rect 416682 158856 416688 158908
rect 416740 158896 416746 158908
rect 419626 158896 419632 158908
rect 416740 158868 419632 158896
rect 416740 158856 416746 158868
rect 419626 158856 419632 158868
rect 419684 158856 419690 158908
rect 452838 158856 452844 158908
rect 452896 158896 452902 158908
rect 464246 158896 464252 158908
rect 452896 158868 464252 158896
rect 452896 158856 452902 158868
rect 464246 158856 464252 158868
rect 464304 158856 464310 158908
rect 466362 158856 466368 158908
rect 466420 158896 466426 158908
rect 472342 158896 472348 158908
rect 466420 158868 472348 158896
rect 466420 158856 466426 158868
rect 472342 158856 472348 158868
rect 472400 158856 472406 158908
rect 474734 158856 474740 158908
rect 474792 158896 474798 158908
rect 480990 158896 480996 158908
rect 474792 158868 480996 158896
rect 474792 158856 474798 158868
rect 480990 158856 480996 158868
rect 481048 158856 481054 158908
rect 508682 158856 508688 158908
rect 508740 158896 508746 158908
rect 510062 158896 510068 158908
rect 508740 158868 510068 158896
rect 508740 158856 508746 158868
rect 510062 158856 510068 158868
rect 510120 158856 510126 158908
rect 383654 158828 383660 158840
rect 374880 158800 379376 158828
rect 379486 158800 383660 158828
rect 374880 158788 374886 158800
rect 367922 158720 367928 158772
rect 367980 158760 367986 158772
rect 374730 158760 374736 158772
rect 367980 158732 374736 158760
rect 367980 158720 367986 158732
rect 374730 158720 374736 158732
rect 374788 158720 374794 158772
rect 379348 158760 379376 158800
rect 383654 158788 383660 158800
rect 383712 158788 383718 158840
rect 387886 158828 387892 158840
rect 384776 158800 387892 158828
rect 384776 158760 384804 158800
rect 387886 158788 387892 158800
rect 387944 158788 387950 158840
rect 388070 158788 388076 158840
rect 388128 158828 388134 158840
rect 390370 158828 390376 158840
rect 388128 158800 390376 158828
rect 388128 158788 388134 158800
rect 390370 158788 390376 158800
rect 390428 158788 390434 158840
rect 456242 158788 456248 158840
rect 456300 158828 456306 158840
rect 466822 158828 466828 158840
rect 456300 158800 466828 158828
rect 456300 158788 456306 158800
rect 466822 158788 466828 158800
rect 466880 158788 466886 158840
rect 476390 158788 476396 158840
rect 476448 158828 476454 158840
rect 482370 158828 482376 158840
rect 476448 158800 482376 158828
rect 476448 158788 476454 158800
rect 482370 158788 482376 158800
rect 482428 158788 482434 158840
rect 506382 158788 506388 158840
rect 506440 158828 506446 158840
rect 507578 158828 507584 158840
rect 506440 158800 507584 158828
rect 506440 158788 506446 158800
rect 507578 158788 507584 158800
rect 507636 158788 507642 158840
rect 379348 158732 384804 158760
rect 413370 158720 413376 158772
rect 413428 158760 413434 158772
rect 419718 158760 419724 158772
rect 413428 158732 419724 158760
rect 413428 158720 413434 158732
rect 419718 158720 419724 158732
rect 419776 158720 419782 158772
rect 464614 158720 464620 158772
rect 464672 158760 464678 158772
rect 471238 158760 471244 158772
rect 464672 158732 471244 158760
rect 464672 158720 464678 158732
rect 471238 158720 471244 158732
rect 471296 158720 471302 158772
rect 473078 158720 473084 158772
rect 473136 158760 473142 158772
rect 479702 158760 479708 158772
rect 473136 158732 479708 158760
rect 473136 158720 473142 158732
rect 479702 158720 479708 158732
rect 479760 158720 479766 158772
rect 481450 158720 481456 158772
rect 481508 158760 481514 158772
rect 486142 158760 486148 158772
rect 481508 158732 486148 158760
rect 481508 158720 481514 158732
rect 486142 158720 486148 158732
rect 486200 158720 486206 158772
rect 504082 158720 504088 158772
rect 504140 158760 504146 158772
rect 505002 158760 505008 158772
rect 504140 158732 505008 158760
rect 504140 158720 504146 158732
rect 505002 158720 505008 158732
rect 505060 158720 505066 158772
rect 506198 158720 506204 158772
rect 506256 158760 506262 158772
rect 506750 158760 506756 158772
rect 506256 158732 506756 158760
rect 506256 158720 506262 158732
rect 506750 158720 506756 158732
rect 506808 158720 506814 158772
rect 507486 158720 507492 158772
rect 507544 158760 507550 158772
rect 508406 158760 508412 158772
rect 507544 158732 508412 158760
rect 507544 158720 507550 158732
rect 508406 158720 508412 158732
rect 508464 158720 508470 158772
rect 509970 158720 509976 158772
rect 510028 158760 510034 158772
rect 511718 158760 511724 158772
rect 510028 158732 511724 158760
rect 510028 158720 510034 158732
rect 511718 158720 511724 158732
rect 511776 158720 511782 158772
rect 515122 158720 515128 158772
rect 515180 158760 515186 158772
rect 518526 158760 518532 158772
rect 515180 158732 518532 158760
rect 515180 158720 515186 158732
rect 518526 158720 518532 158732
rect 518584 158720 518590 158772
rect 374546 158692 374552 158704
rect 367848 158664 374552 158692
rect 374546 158652 374552 158664
rect 374604 158652 374610 158704
rect 74350 158584 74356 158636
rect 74408 158624 74414 158636
rect 175182 158624 175188 158636
rect 74408 158596 175188 158624
rect 74408 158584 74414 158596
rect 175182 158584 175188 158596
rect 175240 158584 175246 158636
rect 175274 158584 175280 158636
rect 175332 158624 175338 158636
rect 252554 158624 252560 158636
rect 175332 158596 252560 158624
rect 175332 158584 175338 158596
rect 252554 158584 252560 158596
rect 252612 158584 252618 158636
rect 71038 158516 71044 158568
rect 71096 158556 71102 158568
rect 172698 158556 172704 158568
rect 71096 158528 172704 158556
rect 71096 158516 71102 158528
rect 172698 158516 172704 158528
rect 172756 158516 172762 158568
rect 178678 158516 178684 158568
rect 178736 158556 178742 158568
rect 255406 158556 255412 158568
rect 178736 158528 255412 158556
rect 178736 158516 178742 158528
rect 255406 158516 255412 158528
rect 255464 158516 255470 158568
rect 361114 158516 361120 158568
rect 361172 158556 361178 158568
rect 362954 158556 362960 158568
rect 361172 158528 362960 158556
rect 361172 158516 361178 158528
rect 362954 158516 362960 158528
rect 363012 158516 363018 158568
rect 67634 158448 67640 158500
rect 67692 158488 67698 158500
rect 170214 158488 170220 158500
rect 67692 158460 170220 158488
rect 67692 158448 67698 158460
rect 170214 158448 170220 158460
rect 170272 158448 170278 158500
rect 171962 158448 171968 158500
rect 172020 158488 172026 158500
rect 249794 158488 249800 158500
rect 172020 158460 249800 158488
rect 172020 158448 172026 158460
rect 249794 158448 249800 158460
rect 249852 158448 249858 158500
rect 60918 158380 60924 158432
rect 60976 158420 60982 158432
rect 165062 158420 165068 158432
rect 60976 158392 165068 158420
rect 60976 158380 60982 158392
rect 165062 158380 165068 158392
rect 165120 158380 165126 158432
rect 165246 158380 165252 158432
rect 165304 158420 165310 158432
rect 244642 158420 244648 158432
rect 165304 158392 244648 158420
rect 165304 158380 165310 158392
rect 244642 158380 244648 158392
rect 244700 158380 244706 158432
rect 64230 158312 64236 158364
rect 64288 158352 64294 158364
rect 167546 158352 167552 158364
rect 64288 158324 167552 158352
rect 64288 158312 64294 158324
rect 167546 158312 167552 158324
rect 167604 158312 167610 158364
rect 168558 158312 168564 158364
rect 168616 158352 168622 158364
rect 247218 158352 247224 158364
rect 168616 158324 247224 158352
rect 168616 158312 168622 158324
rect 247218 158312 247224 158324
rect 247276 158312 247282 158364
rect 54202 158244 54208 158296
rect 54260 158284 54266 158296
rect 160278 158284 160284 158296
rect 54260 158256 160284 158284
rect 54260 158244 54266 158256
rect 160278 158244 160284 158256
rect 160336 158244 160342 158296
rect 161842 158244 161848 158296
rect 161900 158284 161906 158296
rect 242066 158284 242072 158296
rect 161900 158256 242072 158284
rect 161900 158244 161906 158256
rect 242066 158244 242072 158256
rect 242124 158244 242130 158296
rect 50798 158176 50804 158228
rect 50856 158216 50862 158228
rect 157334 158216 157340 158228
rect 50856 158188 157340 158216
rect 50856 158176 50862 158188
rect 157334 158176 157340 158188
rect 157392 158176 157398 158228
rect 158438 158176 158444 158228
rect 158496 158216 158502 158228
rect 239674 158216 239680 158228
rect 158496 158188 239680 158216
rect 158496 158176 158502 158188
rect 239674 158176 239680 158188
rect 239732 158176 239738 158228
rect 256878 158176 256884 158228
rect 256936 158216 256942 158228
rect 314746 158216 314752 158228
rect 256936 158188 314752 158216
rect 256936 158176 256942 158188
rect 314746 158176 314752 158188
rect 314804 158176 314810 158228
rect 47486 158108 47492 158160
rect 47544 158148 47550 158160
rect 154758 158148 154764 158160
rect 47544 158120 154764 158148
rect 47544 158108 47550 158120
rect 154758 158108 154764 158120
rect 154816 158108 154822 158160
rect 155126 158108 155132 158160
rect 155184 158148 155190 158160
rect 237374 158148 237380 158160
rect 155184 158120 237380 158148
rect 155184 158108 155190 158120
rect 237374 158108 237380 158120
rect 237432 158108 237438 158160
rect 246758 158108 246764 158160
rect 246816 158148 246822 158160
rect 306926 158148 306932 158160
rect 246816 158120 306932 158148
rect 246816 158108 246822 158120
rect 306926 158108 306932 158120
rect 306984 158108 306990 158160
rect 37366 158040 37372 158092
rect 37424 158080 37430 158092
rect 147122 158080 147128 158092
rect 37424 158052 147128 158080
rect 37424 158040 37430 158052
rect 147122 158040 147128 158052
rect 147180 158040 147186 158092
rect 148410 158040 148416 158092
rect 148468 158080 148474 158092
rect 231854 158080 231860 158092
rect 148468 158052 231860 158080
rect 148468 158040 148474 158052
rect 231854 158040 231860 158052
rect 231912 158040 231918 158092
rect 243446 158040 243452 158092
rect 243504 158080 243510 158092
rect 304350 158080 304356 158092
rect 243504 158052 304356 158080
rect 243504 158040 243510 158052
rect 304350 158040 304356 158052
rect 304408 158040 304414 158092
rect 382 157972 388 158024
rect 440 158012 446 158024
rect 118878 158012 118884 158024
rect 440 157984 118884 158012
rect 440 157972 446 157984
rect 118878 157972 118884 157984
rect 118936 157972 118942 158024
rect 122742 157972 122748 158024
rect 122800 158012 122806 158024
rect 123386 158012 123392 158024
rect 122800 157984 123392 158012
rect 122800 157972 122806 157984
rect 123386 157972 123392 157984
rect 123444 157972 123450 158024
rect 131574 157972 131580 158024
rect 131632 158012 131638 158024
rect 218974 158012 218980 158024
rect 131632 157984 218980 158012
rect 131632 157972 131638 157984
rect 218974 157972 218980 157984
rect 219032 157972 219038 158024
rect 236730 157972 236736 158024
rect 236788 158012 236794 158024
rect 299566 158012 299572 158024
rect 236788 157984 299572 158012
rect 236788 157972 236794 157984
rect 299566 157972 299572 157984
rect 299624 157972 299630 158024
rect 77754 157904 77760 157956
rect 77812 157944 77818 157956
rect 77812 157916 176056 157944
rect 77812 157904 77818 157916
rect 84470 157836 84476 157888
rect 84528 157876 84534 157888
rect 175918 157876 175924 157888
rect 84528 157848 175924 157876
rect 84528 157836 84534 157848
rect 175918 157836 175924 157848
rect 175976 157836 175982 157888
rect 176028 157876 176056 157916
rect 176194 157904 176200 157956
rect 176252 157944 176258 157956
rect 182818 157944 182824 157956
rect 176252 157916 182824 157944
rect 176252 157904 176258 157916
rect 182818 157904 182824 157916
rect 182876 157904 182882 157956
rect 185394 157904 185400 157956
rect 185452 157944 185458 157956
rect 260190 157944 260196 157956
rect 185452 157916 260196 157944
rect 185452 157904 185458 157916
rect 260190 157904 260196 157916
rect 260248 157904 260254 157956
rect 178034 157876 178040 157888
rect 176028 157848 178040 157876
rect 178034 157836 178040 157848
rect 178092 157836 178098 157888
rect 181530 157836 181536 157888
rect 181588 157876 181594 157888
rect 188154 157876 188160 157888
rect 181588 157848 188160 157876
rect 181588 157836 181594 157848
rect 188154 157836 188160 157848
rect 188212 157836 188218 157888
rect 188798 157836 188804 157888
rect 188856 157876 188862 157888
rect 262674 157876 262680 157888
rect 188856 157848 262680 157876
rect 188856 157836 188862 157848
rect 262674 157836 262680 157848
rect 262732 157836 262738 157888
rect 87782 157768 87788 157820
rect 87840 157808 87846 157820
rect 181622 157808 181628 157820
rect 87840 157780 181628 157808
rect 87840 157768 87846 157780
rect 181622 157768 181628 157780
rect 181680 157768 181686 157820
rect 181806 157768 181812 157820
rect 181864 157808 181870 157820
rect 190638 157808 190644 157820
rect 181864 157780 190644 157808
rect 181864 157768 181870 157780
rect 190638 157768 190644 157780
rect 190696 157768 190702 157820
rect 195514 157768 195520 157820
rect 195572 157808 195578 157820
rect 267734 157808 267740 157820
rect 195572 157780 267740 157808
rect 195572 157768 195578 157780
rect 267734 157768 267740 157780
rect 267792 157768 267798 157820
rect 91186 157700 91192 157752
rect 91244 157740 91250 157752
rect 181254 157740 181260 157752
rect 91244 157712 181260 157740
rect 91244 157700 91250 157712
rect 181254 157700 181260 157712
rect 181312 157700 181318 157752
rect 181898 157700 181904 157752
rect 181956 157740 181962 157752
rect 181956 157712 186314 157740
rect 181956 157700 181962 157712
rect 94590 157632 94596 157684
rect 94648 157672 94654 157684
rect 181530 157672 181536 157684
rect 94648 157644 181536 157672
rect 94648 157632 94654 157644
rect 181530 157632 181536 157644
rect 181588 157632 181594 157684
rect 181714 157632 181720 157684
rect 181772 157672 181778 157684
rect 185578 157672 185584 157684
rect 181772 157644 185584 157672
rect 181772 157632 181778 157644
rect 185578 157632 185584 157644
rect 185636 157632 185642 157684
rect 186286 157672 186314 157712
rect 190454 157700 190460 157752
rect 190512 157740 190518 157752
rect 264054 157740 264060 157752
rect 190512 157712 264060 157740
rect 190512 157700 190518 157712
rect 264054 157700 264060 157712
rect 264112 157700 264118 157752
rect 236086 157672 236092 157684
rect 186286 157644 236092 157672
rect 236086 157632 236092 157644
rect 236144 157632 236150 157684
rect 97902 157564 97908 157616
rect 97960 157604 97966 157616
rect 193214 157604 193220 157616
rect 97960 157576 193220 157604
rect 97960 157564 97966 157576
rect 193214 157564 193220 157576
rect 193272 157564 193278 157616
rect 197354 157564 197360 157616
rect 197412 157604 197418 157616
rect 251266 157604 251272 157616
rect 197412 157576 251272 157604
rect 197412 157564 197418 157576
rect 251266 157564 251272 157576
rect 251324 157564 251330 157616
rect 111334 157496 111340 157548
rect 111392 157536 111398 157548
rect 203426 157536 203432 157548
rect 111392 157508 203432 157536
rect 111392 157496 111398 157508
rect 203426 157496 203432 157508
rect 203484 157496 203490 157548
rect 204898 157496 204904 157548
rect 204956 157536 204962 157548
rect 256326 157536 256332 157548
rect 204956 157508 256332 157536
rect 204956 157496 204962 157508
rect 256326 157496 256332 157508
rect 256384 157496 256390 157548
rect 114738 157428 114744 157480
rect 114796 157468 114802 157480
rect 206186 157468 206192 157480
rect 114796 157440 206192 157468
rect 114796 157428 114802 157440
rect 206186 157428 206192 157440
rect 206244 157428 206250 157480
rect 141694 157360 141700 157412
rect 141752 157400 141758 157412
rect 226702 157400 226708 157412
rect 141752 157372 226708 157400
rect 141752 157360 141758 157372
rect 226702 157360 226708 157372
rect 226760 157360 226766 157412
rect 49142 157292 49148 157344
rect 49200 157332 49206 157344
rect 156046 157332 156052 157344
rect 49200 157304 156052 157332
rect 49200 157292 49206 157304
rect 156046 157292 156052 157304
rect 156104 157292 156110 157344
rect 156322 157292 156328 157344
rect 156380 157332 156386 157344
rect 212534 157332 212540 157344
rect 156380 157304 212540 157332
rect 156380 157292 156386 157304
rect 212534 157292 212540 157304
rect 212592 157292 212598 157344
rect 213178 157292 213184 157344
rect 213236 157332 213242 157344
rect 281626 157332 281632 157344
rect 213236 157304 281632 157332
rect 213236 157292 213242 157304
rect 281626 157292 281632 157304
rect 281684 157292 281690 157344
rect 45738 157224 45744 157276
rect 45796 157264 45802 157276
rect 153470 157264 153476 157276
rect 45796 157236 153476 157264
rect 45796 157224 45802 157236
rect 153470 157224 153476 157236
rect 153528 157224 153534 157276
rect 192110 157224 192116 157276
rect 192168 157264 192174 157276
rect 265158 157264 265164 157276
rect 192168 157236 265164 157264
rect 192168 157224 192174 157236
rect 265158 157224 265164 157236
rect 265216 157224 265222 157276
rect 39022 157156 39028 157208
rect 39080 157196 39086 157208
rect 148226 157196 148232 157208
rect 39080 157168 148232 157196
rect 39080 157156 39086 157168
rect 148226 157156 148232 157168
rect 148284 157156 148290 157208
rect 160094 157156 160100 157208
rect 160152 157196 160158 157208
rect 164050 157196 164056 157208
rect 160152 157168 164056 157196
rect 160152 157156 160158 157168
rect 164050 157156 164056 157168
rect 164108 157156 164114 157208
rect 164142 157156 164148 157208
rect 164200 157196 164206 157208
rect 171594 157196 171600 157208
rect 164200 157168 171600 157196
rect 164200 157156 164206 157168
rect 171594 157156 171600 157168
rect 171652 157156 171658 157208
rect 177022 157156 177028 157208
rect 177080 157196 177086 157208
rect 254026 157196 254032 157208
rect 177080 157168 254032 157196
rect 177080 157156 177086 157168
rect 254026 157156 254032 157168
rect 254084 157156 254090 157208
rect 290550 157156 290556 157208
rect 290608 157196 290614 157208
rect 339954 157196 339960 157208
rect 290608 157168 339960 157196
rect 290608 157156 290614 157168
rect 339954 157156 339960 157168
rect 340012 157156 340018 157208
rect 42426 157088 42432 157140
rect 42484 157128 42490 157140
rect 150894 157128 150900 157140
rect 42484 157100 150900 157128
rect 42484 157088 42490 157100
rect 150894 157088 150900 157100
rect 150952 157088 150958 157140
rect 151722 157088 151728 157140
rect 151780 157128 151786 157140
rect 234614 157128 234620 157140
rect 151780 157100 234620 157128
rect 151780 157088 151786 157100
rect 234614 157088 234620 157100
rect 234672 157088 234678 157140
rect 287146 157088 287152 157140
rect 287204 157128 287210 157140
rect 338114 157128 338120 157140
rect 287204 157100 338120 157128
rect 287204 157088 287210 157100
rect 338114 157088 338120 157100
rect 338172 157088 338178 157140
rect 35710 157020 35716 157072
rect 35768 157060 35774 157072
rect 35768 157032 138014 157060
rect 35768 157020 35774 157032
rect 24762 156952 24768 157004
rect 24820 156992 24826 157004
rect 137554 156992 137560 157004
rect 24820 156964 137560 156992
rect 24820 156952 24826 156964
rect 137554 156952 137560 156964
rect 137612 156952 137618 157004
rect 137986 156992 138014 157032
rect 145006 157020 145012 157072
rect 145064 157060 145070 157072
rect 229278 157060 229284 157072
rect 145064 157032 229284 157060
rect 145064 157020 145070 157032
rect 229278 157020 229284 157032
rect 229336 157020 229342 157072
rect 231026 157020 231032 157072
rect 231084 157060 231090 157072
rect 276842 157060 276848 157072
rect 231084 157032 276848 157060
rect 231084 157020 231090 157032
rect 276842 157020 276848 157032
rect 276900 157020 276906 157072
rect 280430 157020 280436 157072
rect 280488 157060 280494 157072
rect 332686 157060 332692 157072
rect 280488 157032 332692 157060
rect 280488 157020 280494 157032
rect 332686 157020 332692 157032
rect 332744 157020 332750 157072
rect 146018 156992 146024 157004
rect 137986 156964 146024 156992
rect 146018 156952 146024 156964
rect 146076 156952 146082 157004
rect 150066 156952 150072 157004
rect 150124 156992 150130 157004
rect 233234 156992 233240 157004
rect 150124 156964 233240 156992
rect 150124 156952 150130 156964
rect 233234 156952 233240 156964
rect 233292 156952 233298 157004
rect 283834 156952 283840 157004
rect 283892 156992 283898 157004
rect 335446 156992 335452 157004
rect 283892 156964 335452 156992
rect 283892 156952 283898 156964
rect 335446 156952 335452 156964
rect 335504 156952 335510 157004
rect 18046 156884 18052 156936
rect 18104 156924 18110 156936
rect 132494 156924 132500 156936
rect 18104 156896 132500 156924
rect 18104 156884 18110 156896
rect 132494 156884 132500 156896
rect 132552 156884 132558 156936
rect 138290 156884 138296 156936
rect 138348 156924 138354 156936
rect 224126 156924 224132 156936
rect 138348 156896 224132 156924
rect 138348 156884 138354 156896
rect 224126 156884 224132 156896
rect 224184 156884 224190 156936
rect 273714 156884 273720 156936
rect 273772 156924 273778 156936
rect 327534 156924 327540 156936
rect 273772 156896 327540 156924
rect 273772 156884 273778 156896
rect 327534 156884 327540 156896
rect 327592 156884 327598 156936
rect 21358 156816 21364 156868
rect 21416 156856 21422 156868
rect 135254 156856 135260 156868
rect 21416 156828 135260 156856
rect 21416 156816 21422 156828
rect 135254 156816 135260 156828
rect 135312 156816 135318 156868
rect 135806 156816 135812 156868
rect 135864 156856 135870 156868
rect 222194 156856 222200 156868
rect 135864 156828 222200 156856
rect 135864 156816 135870 156828
rect 222194 156816 222200 156828
rect 222252 156816 222258 156868
rect 224954 156816 224960 156868
rect 225012 156856 225018 156868
rect 271966 156856 271972 156868
rect 225012 156828 271972 156856
rect 225012 156816 225018 156828
rect 271966 156816 271972 156828
rect 272024 156816 272030 156868
rect 277118 156816 277124 156868
rect 277176 156856 277182 156868
rect 330018 156856 330024 156868
rect 277176 156828 330024 156856
rect 277176 156816 277182 156828
rect 330018 156816 330024 156828
rect 330076 156816 330082 156868
rect 11238 156748 11244 156800
rect 11296 156788 11302 156800
rect 127158 156788 127164 156800
rect 11296 156760 127164 156788
rect 11296 156748 11302 156760
rect 127158 156748 127164 156760
rect 127216 156748 127222 156800
rect 139118 156748 139124 156800
rect 139176 156788 139182 156800
rect 225046 156788 225052 156800
rect 139176 156760 225052 156788
rect 139176 156748 139182 156760
rect 225046 156748 225052 156760
rect 225104 156748 225110 156800
rect 226610 156748 226616 156800
rect 226668 156788 226674 156800
rect 291562 156788 291568 156800
rect 226668 156760 291568 156788
rect 226668 156748 226674 156760
rect 291562 156748 291568 156760
rect 291620 156748 291626 156800
rect 297266 156748 297272 156800
rect 297324 156788 297330 156800
rect 345566 156788 345572 156800
rect 297324 156760 345572 156788
rect 297324 156748 297330 156760
rect 345566 156748 345572 156760
rect 345624 156748 345630 156800
rect 14642 156680 14648 156732
rect 14700 156720 14706 156732
rect 129826 156720 129832 156732
rect 14700 156692 129832 156720
rect 14700 156680 14706 156692
rect 129826 156680 129832 156692
rect 129884 156680 129890 156732
rect 134886 156680 134892 156732
rect 134944 156720 134950 156732
rect 221366 156720 221372 156732
rect 134944 156692 221372 156720
rect 134944 156680 134950 156692
rect 221366 156680 221372 156692
rect 221424 156680 221430 156732
rect 230014 156680 230020 156732
rect 230072 156720 230078 156732
rect 294046 156720 294052 156732
rect 230072 156692 294052 156720
rect 230072 156680 230078 156692
rect 294046 156680 294052 156692
rect 294104 156680 294110 156732
rect 300670 156680 300676 156732
rect 300728 156720 300734 156732
rect 348050 156720 348056 156732
rect 300728 156692 348056 156720
rect 300728 156680 300734 156692
rect 348050 156680 348056 156692
rect 348108 156680 348114 156732
rect 2038 156612 2044 156664
rect 2096 156652 2102 156664
rect 120166 156652 120172 156664
rect 2096 156624 120172 156652
rect 2096 156612 2102 156624
rect 120166 156612 120172 156624
rect 120224 156612 120230 156664
rect 128170 156612 128176 156664
rect 128228 156652 128234 156664
rect 216674 156652 216680 156664
rect 128228 156624 216680 156652
rect 128228 156612 128234 156624
rect 216674 156612 216680 156624
rect 216732 156612 216738 156664
rect 223206 156612 223212 156664
rect 223264 156652 223270 156664
rect 288986 156652 288992 156664
rect 223264 156624 288992 156652
rect 223264 156612 223270 156624
rect 288986 156612 288992 156624
rect 289044 156612 289050 156664
rect 293862 156612 293868 156664
rect 293920 156652 293926 156664
rect 342254 156652 342260 156664
rect 293920 156624 342260 156652
rect 293920 156612 293926 156624
rect 342254 156612 342260 156624
rect 342312 156612 342318 156664
rect 52454 156544 52460 156596
rect 52512 156584 52518 156596
rect 158622 156584 158628 156596
rect 52512 156556 158628 156584
rect 52512 156544 52518 156556
rect 158622 156544 158628 156556
rect 158680 156544 158686 156596
rect 158714 156544 158720 156596
rect 158772 156584 158778 156596
rect 219986 156584 219992 156596
rect 158772 156556 219992 156584
rect 158772 156544 158778 156556
rect 219986 156544 219992 156556
rect 220044 156544 220050 156596
rect 59262 156476 59268 156528
rect 59320 156516 59326 156528
rect 163774 156516 163780 156528
rect 59320 156488 163780 156516
rect 59320 156476 59326 156488
rect 163774 156476 163780 156488
rect 163832 156476 163838 156528
rect 164050 156476 164056 156528
rect 164108 156516 164114 156528
rect 164108 156488 164280 156516
rect 164108 156476 164114 156488
rect 69290 156408 69296 156460
rect 69348 156448 69354 156460
rect 164142 156448 164148 156460
rect 69348 156420 164148 156448
rect 69348 156408 69354 156420
rect 164142 156408 164148 156420
rect 164200 156408 164206 156460
rect 164252 156448 164280 156488
rect 164326 156476 164332 156528
rect 164384 156516 164390 156528
rect 225506 156516 225512 156528
rect 164384 156488 225512 156516
rect 164384 156476 164390 156488
rect 225506 156476 225512 156488
rect 225564 156476 225570 156528
rect 227990 156448 227996 156460
rect 164252 156420 227996 156448
rect 227990 156408 227996 156420
rect 228048 156408 228054 156460
rect 82814 156340 82820 156392
rect 82872 156380 82878 156392
rect 181806 156380 181812 156392
rect 82872 156352 181812 156380
rect 82872 156340 82878 156352
rect 181806 156340 181812 156352
rect 181864 156340 181870 156392
rect 198826 156340 198832 156392
rect 198884 156380 198890 156392
rect 200942 156380 200948 156392
rect 198884 156352 200948 156380
rect 198884 156340 198890 156352
rect 200942 156340 200948 156352
rect 201000 156340 201006 156392
rect 209774 156340 209780 156392
rect 209832 156380 209838 156392
rect 278866 156380 278872 156392
rect 209832 156352 278872 156380
rect 209832 156340 209838 156352
rect 278866 156340 278872 156352
rect 278924 156340 278930 156392
rect 101306 156272 101312 156324
rect 101364 156312 101370 156324
rect 196158 156312 196164 156324
rect 101364 156284 196164 156312
rect 101364 156272 101370 156284
rect 196158 156272 196164 156284
rect 196216 156272 196222 156324
rect 200758 156272 200764 156324
rect 200816 156312 200822 156324
rect 211338 156312 211344 156324
rect 200816 156284 211344 156312
rect 200816 156272 200822 156284
rect 211338 156272 211344 156284
rect 211396 156272 211402 156324
rect 212534 156272 212540 156324
rect 212592 156312 212598 156324
rect 215386 156312 215392 156324
rect 212592 156284 215392 156312
rect 212592 156272 212598 156284
rect 215386 156272 215392 156284
rect 215444 156272 215450 156324
rect 216490 156272 216496 156324
rect 216548 156312 216554 156324
rect 283466 156312 283472 156324
rect 216548 156284 283472 156312
rect 216548 156272 216554 156284
rect 283466 156272 283472 156284
rect 283524 156272 283530 156324
rect 99558 156204 99564 156256
rect 99616 156244 99622 156256
rect 194686 156244 194692 156256
rect 99616 156216 194692 156244
rect 99616 156204 99622 156216
rect 194686 156204 194692 156216
rect 194744 156204 194750 156256
rect 200776 156216 200988 156244
rect 108022 156136 108028 156188
rect 108080 156176 108086 156188
rect 200666 156176 200672 156188
rect 108080 156148 200672 156176
rect 108080 156136 108086 156148
rect 200666 156136 200672 156148
rect 200724 156136 200730 156188
rect 118142 156068 118148 156120
rect 118200 156108 118206 156120
rect 200776 156108 200804 156216
rect 200960 156176 200988 156216
rect 203058 156204 203064 156256
rect 203116 156244 203122 156256
rect 203116 156216 214604 156244
rect 203116 156204 203122 156216
rect 208762 156176 208768 156188
rect 200960 156148 208768 156176
rect 208762 156136 208768 156148
rect 208820 156136 208826 156188
rect 118200 156080 200804 156108
rect 118200 156068 118206 156080
rect 200942 156068 200948 156120
rect 201000 156108 201006 156120
rect 214576 156108 214604 156216
rect 219894 156204 219900 156256
rect 219952 156244 219958 156256
rect 285674 156244 285680 156256
rect 219952 156216 285680 156244
rect 219952 156204 219958 156216
rect 285674 156204 285680 156216
rect 285732 156204 285738 156256
rect 218054 156136 218060 156188
rect 218112 156176 218118 156188
rect 266538 156176 266544 156188
rect 218112 156148 266544 156176
rect 218112 156136 218118 156148
rect 266538 156136 266544 156148
rect 266596 156136 266602 156188
rect 273530 156108 273536 156120
rect 201000 156080 214512 156108
rect 214576 156080 273536 156108
rect 201000 156068 201006 156080
rect 121454 156000 121460 156052
rect 121512 156040 121518 156052
rect 200758 156040 200764 156052
rect 121512 156012 200764 156040
rect 121512 156000 121518 156012
rect 200758 156000 200764 156012
rect 200816 156000 200822 156052
rect 202230 156000 202236 156052
rect 202288 156040 202294 156052
rect 214282 156040 214288 156052
rect 202288 156012 214288 156040
rect 202288 156000 202294 156012
rect 214282 156000 214288 156012
rect 214340 156000 214346 156052
rect 124858 155932 124864 155984
rect 124916 155972 124922 155984
rect 213914 155972 213920 155984
rect 124916 155944 213920 155972
rect 124916 155932 124922 155944
rect 213914 155932 213920 155944
rect 213972 155932 213978 155984
rect 214484 155972 214512 156080
rect 273530 156068 273536 156080
rect 273588 156068 273594 156120
rect 214558 156000 214564 156052
rect 214616 156040 214622 156052
rect 273254 156040 273260 156052
rect 214616 156012 273260 156040
rect 214616 156000 214622 156012
rect 273254 156000 273260 156012
rect 273312 156000 273318 156052
rect 270494 155972 270500 155984
rect 214484 155944 270500 155972
rect 270494 155932 270500 155944
rect 270552 155932 270558 155984
rect 89530 155864 89536 155916
rect 89588 155904 89594 155916
rect 186958 155904 186964 155916
rect 89588 155876 186964 155904
rect 89588 155864 89594 155876
rect 186958 155864 186964 155876
rect 187016 155864 187022 155916
rect 192938 155864 192944 155916
rect 192996 155904 193002 155916
rect 265894 155904 265900 155916
rect 192996 155876 265900 155904
rect 192996 155864 193002 155876
rect 265894 155864 265900 155876
rect 265952 155864 265958 155916
rect 293034 155864 293040 155916
rect 293092 155904 293098 155916
rect 342346 155904 342352 155916
rect 293092 155876 342352 155904
rect 293092 155864 293098 155876
rect 342346 155864 342352 155876
rect 342404 155864 342410 155916
rect 53374 155796 53380 155848
rect 53432 155836 53438 155848
rect 66714 155836 66720 155848
rect 53432 155808 66720 155836
rect 53432 155796 53438 155808
rect 66714 155796 66720 155808
rect 66772 155796 66778 155848
rect 66806 155796 66812 155848
rect 66864 155836 66870 155848
rect 82906 155836 82912 155848
rect 66864 155808 82912 155836
rect 66864 155796 66870 155808
rect 82906 155796 82912 155808
rect 82964 155796 82970 155848
rect 88702 155796 88708 155848
rect 88760 155836 88766 155848
rect 186406 155836 186412 155848
rect 88760 155808 186412 155836
rect 88760 155796 88766 155808
rect 186406 155796 186412 155808
rect 186464 155796 186470 155848
rect 189626 155796 189632 155848
rect 189684 155836 189690 155848
rect 263686 155836 263692 155848
rect 189684 155808 263692 155836
rect 189684 155796 189690 155808
rect 263686 155796 263692 155808
rect 263744 155796 263750 155848
rect 296438 155796 296444 155848
rect 296496 155836 296502 155848
rect 345106 155836 345112 155848
rect 296496 155808 345112 155836
rect 296496 155796 296502 155808
rect 345106 155796 345112 155808
rect 345164 155796 345170 155848
rect 12158 155728 12164 155780
rect 12216 155768 12222 155780
rect 109770 155768 109776 155780
rect 12216 155740 109776 155768
rect 12216 155728 12222 155740
rect 109770 155728 109776 155740
rect 109828 155728 109834 155780
rect 112254 155728 112260 155780
rect 112312 155768 112318 155780
rect 204346 155768 204352 155780
rect 112312 155740 204352 155768
rect 112312 155728 112318 155740
rect 204346 155728 204352 155740
rect 204404 155728 204410 155780
rect 206462 155728 206468 155780
rect 206520 155768 206526 155780
rect 276106 155768 276112 155780
rect 206520 155740 276112 155768
rect 206520 155728 206526 155740
rect 276106 155728 276112 155740
rect 276164 155728 276170 155780
rect 289722 155728 289728 155780
rect 289780 155768 289786 155780
rect 339586 155768 339592 155780
rect 289780 155740 339592 155768
rect 289780 155728 289786 155740
rect 339586 155728 339592 155740
rect 339644 155728 339650 155780
rect 60090 155660 60096 155712
rect 60148 155700 60154 155712
rect 78858 155700 78864 155712
rect 60148 155672 78864 155700
rect 60148 155660 60154 155672
rect 78858 155660 78864 155672
rect 78916 155660 78922 155712
rect 81894 155660 81900 155712
rect 81952 155700 81958 155712
rect 181162 155700 181168 155712
rect 81952 155672 181168 155700
rect 81952 155660 81958 155672
rect 181162 155660 181168 155672
rect 181220 155660 181226 155712
rect 186222 155660 186228 155712
rect 186280 155700 186286 155712
rect 260834 155700 260840 155712
rect 186280 155672 260840 155700
rect 186280 155660 186286 155672
rect 260834 155660 260840 155672
rect 260892 155660 260898 155712
rect 266998 155660 267004 155712
rect 267056 155700 267062 155712
rect 322106 155700 322112 155712
rect 267056 155672 322112 155700
rect 267056 155660 267062 155672
rect 322106 155660 322112 155672
rect 322164 155660 322170 155712
rect 340966 155660 340972 155712
rect 341024 155700 341030 155712
rect 378686 155700 378692 155712
rect 341024 155672 378692 155700
rect 341024 155660 341030 155672
rect 378686 155660 378692 155672
rect 378744 155660 378750 155712
rect 46566 155592 46572 155644
rect 46624 155632 46630 155644
rect 75086 155632 75092 155644
rect 46624 155604 75092 155632
rect 46624 155592 46630 155604
rect 75086 155592 75092 155604
rect 75144 155592 75150 155644
rect 75178 155592 75184 155644
rect 75236 155632 75242 155644
rect 176010 155632 176016 155644
rect 75236 155604 176016 155632
rect 75236 155592 75242 155604
rect 176010 155592 176016 155604
rect 176068 155592 176074 155644
rect 179506 155592 179512 155644
rect 179564 155632 179570 155644
rect 255590 155632 255596 155644
rect 179564 155604 255596 155632
rect 179564 155592 179570 155604
rect 255590 155592 255596 155604
rect 255648 155592 255654 155644
rect 270310 155592 270316 155644
rect 270368 155632 270374 155644
rect 324958 155632 324964 155644
rect 270368 155604 324964 155632
rect 270368 155592 270374 155604
rect 324958 155592 324964 155604
rect 325016 155592 325022 155644
rect 344370 155592 344376 155644
rect 344428 155632 344434 155644
rect 381446 155632 381452 155644
rect 344428 155604 381452 155632
rect 344428 155592 344434 155604
rect 381446 155592 381452 155604
rect 381504 155592 381510 155644
rect 39850 155524 39856 155576
rect 39908 155564 39914 155576
rect 68922 155564 68928 155576
rect 39908 155536 68928 155564
rect 39908 155524 39914 155536
rect 68922 155524 68928 155536
rect 68980 155524 68986 155576
rect 71866 155524 71872 155576
rect 71924 155564 71930 155576
rect 173066 155564 173072 155576
rect 71924 155536 173072 155564
rect 71924 155524 71930 155536
rect 173066 155524 173072 155536
rect 173124 155524 173130 155576
rect 176286 155524 176292 155576
rect 176344 155564 176350 155576
rect 253014 155564 253020 155576
rect 176344 155536 253020 155564
rect 176344 155524 176350 155536
rect 253014 155524 253020 155536
rect 253072 155524 253078 155576
rect 263594 155524 263600 155576
rect 263652 155564 263658 155576
rect 320174 155564 320180 155576
rect 263652 155536 320180 155564
rect 263652 155524 263658 155536
rect 320174 155524 320180 155536
rect 320232 155524 320238 155576
rect 337654 155524 337660 155576
rect 337712 155564 337718 155576
rect 376294 155564 376300 155576
rect 337712 155536 376300 155564
rect 337712 155524 337718 155536
rect 376294 155524 376300 155536
rect 376352 155524 376358 155576
rect 65150 155456 65156 155508
rect 65208 155496 65214 155508
rect 168374 155496 168380 155508
rect 65208 155468 168380 155496
rect 65208 155456 65214 155468
rect 168374 155456 168380 155468
rect 168432 155456 168438 155508
rect 169386 155456 169392 155508
rect 169444 155496 169450 155508
rect 247954 155496 247960 155508
rect 169444 155468 247960 155496
rect 169444 155456 169450 155468
rect 247954 155456 247960 155468
rect 248012 155456 248018 155508
rect 260282 155456 260288 155508
rect 260340 155496 260346 155508
rect 317506 155496 317512 155508
rect 260340 155468 317512 155496
rect 260340 155456 260346 155468
rect 317506 155456 317512 155468
rect 317564 155456 317570 155508
rect 333422 155456 333428 155508
rect 333480 155496 333486 155508
rect 373074 155496 373080 155508
rect 333480 155468 373080 155496
rect 333480 155456 333486 155468
rect 373074 155456 373080 155468
rect 373132 155456 373138 155508
rect 4522 155388 4528 155440
rect 4580 155428 4586 155440
rect 122006 155428 122012 155440
rect 4580 155400 122012 155428
rect 4580 155388 4586 155400
rect 122006 155388 122012 155400
rect 122064 155388 122070 155440
rect 122282 155388 122288 155440
rect 122340 155428 122346 155440
rect 211982 155428 211988 155440
rect 122340 155400 211988 155428
rect 122340 155388 122346 155400
rect 211982 155388 211988 155400
rect 212040 155388 212046 155440
rect 214098 155388 214104 155440
rect 214156 155428 214162 155440
rect 261386 155428 261392 155440
rect 214156 155400 261392 155428
rect 214156 155388 214162 155400
rect 261386 155388 261392 155400
rect 261444 155388 261450 155440
rect 330110 155388 330116 155440
rect 330168 155428 330174 155440
rect 370590 155428 370596 155440
rect 330168 155400 370596 155428
rect 330168 155388 330174 155400
rect 370590 155388 370596 155400
rect 370648 155388 370654 155440
rect 7926 155320 7932 155372
rect 7984 155360 7990 155372
rect 124582 155360 124588 155372
rect 7984 155332 124588 155360
rect 7984 155320 7990 155332
rect 124582 155320 124588 155332
rect 124640 155320 124646 155372
rect 142522 155320 142528 155372
rect 142580 155360 142586 155372
rect 227806 155360 227812 155372
rect 142580 155332 227812 155360
rect 142580 155320 142586 155332
rect 227806 155320 227812 155332
rect 227864 155320 227870 155372
rect 253566 155320 253572 155372
rect 253624 155360 253630 155372
rect 312078 155360 312084 155372
rect 253624 155332 312084 155360
rect 253624 155320 253630 155332
rect 312078 155320 312084 155332
rect 312136 155320 312142 155372
rect 319990 155320 319996 155372
rect 320048 155360 320054 155372
rect 363046 155360 363052 155372
rect 320048 155332 363052 155360
rect 320048 155320 320054 155332
rect 363046 155320 363052 155332
rect 363104 155320 363110 155372
rect 8754 155252 8760 155304
rect 8812 155292 8818 155304
rect 125594 155292 125600 155304
rect 8812 155264 125600 155292
rect 8812 155252 8818 155264
rect 125594 155252 125600 155264
rect 125652 155252 125658 155304
rect 128998 155252 129004 155304
rect 129056 155292 129062 155304
rect 217042 155292 217048 155304
rect 129056 155264 217048 155292
rect 129056 155252 129062 155264
rect 217042 155252 217048 155264
rect 217100 155252 217106 155304
rect 233326 155252 233332 155304
rect 233384 155292 233390 155304
rect 296806 155292 296812 155304
rect 233384 155264 296812 155292
rect 233384 155252 233390 155264
rect 296806 155252 296812 155264
rect 296864 155252 296870 155304
rect 299750 155252 299756 155304
rect 299808 155292 299814 155304
rect 347774 155292 347780 155304
rect 299808 155264 347780 155292
rect 299808 155252 299814 155264
rect 347774 155252 347780 155264
rect 347832 155252 347838 155304
rect 373810 155252 373816 155304
rect 373868 155292 373874 155304
rect 403526 155292 403532 155304
rect 373868 155264 403532 155292
rect 373868 155252 373874 155264
rect 403526 155252 403532 155264
rect 403584 155252 403590 155304
rect 5350 155184 5356 155236
rect 5408 155224 5414 155236
rect 122926 155224 122932 155236
rect 5408 155196 122932 155224
rect 5408 155184 5414 155196
rect 122926 155184 122932 155196
rect 122984 155184 122990 155236
rect 125686 155184 125692 155236
rect 125744 155224 125750 155236
rect 214466 155224 214472 155236
rect 125744 155196 214472 155224
rect 125744 155184 125750 155196
rect 214466 155184 214472 155196
rect 214524 155184 214530 155236
rect 240042 155184 240048 155236
rect 240100 155224 240106 155236
rect 302326 155224 302332 155236
rect 240100 155196 302332 155224
rect 240100 155184 240106 155196
rect 302326 155184 302332 155196
rect 302384 155184 302390 155236
rect 303154 155184 303160 155236
rect 303212 155224 303218 155236
rect 350074 155224 350080 155236
rect 303212 155196 350080 155224
rect 303212 155184 303218 155196
rect 350074 155184 350080 155196
rect 350132 155184 350138 155236
rect 370406 155184 370412 155236
rect 370464 155224 370470 155236
rect 401686 155224 401692 155236
rect 370464 155196 401692 155224
rect 370464 155184 370470 155196
rect 401686 155184 401692 155196
rect 401744 155184 401750 155236
rect 92014 155116 92020 155168
rect 92072 155156 92078 155168
rect 189074 155156 189080 155168
rect 92072 155128 189080 155156
rect 92072 155116 92078 155128
rect 189074 155116 189080 155128
rect 189132 155116 189138 155168
rect 189166 155116 189172 155168
rect 189224 155156 189230 155168
rect 194042 155156 194048 155168
rect 189224 155128 194048 155156
rect 189224 155116 189230 155128
rect 194042 155116 194048 155128
rect 194100 155116 194106 155168
rect 196342 155116 196348 155168
rect 196400 155156 196406 155168
rect 268470 155156 268476 155168
rect 196400 155128 268476 155156
rect 196400 155116 196406 155128
rect 268470 155116 268476 155128
rect 268528 155116 268534 155168
rect 306558 155116 306564 155168
rect 306616 155156 306622 155168
rect 352466 155156 352472 155168
rect 306616 155128 352472 155156
rect 306616 155116 306622 155128
rect 352466 155116 352472 155128
rect 352524 155116 352530 155168
rect 95418 155048 95424 155100
rect 95476 155088 95482 155100
rect 95476 155060 186452 155088
rect 95476 155048 95482 155060
rect 98730 154980 98736 155032
rect 98788 155020 98794 155032
rect 186314 155020 186320 155032
rect 98788 154992 186320 155020
rect 98788 154980 98794 154992
rect 186314 154980 186320 154992
rect 186372 154980 186378 155032
rect 186424 155020 186452 155060
rect 186774 155048 186780 155100
rect 186832 155088 186838 155100
rect 186832 155060 195974 155088
rect 186832 155048 186838 155060
rect 191466 155020 191472 155032
rect 186424 154992 191472 155020
rect 191466 154980 191472 154992
rect 191524 154980 191530 155032
rect 195946 155020 195974 155060
rect 199654 155048 199660 155100
rect 199712 155088 199718 155100
rect 271046 155088 271052 155100
rect 199712 155060 271052 155088
rect 199712 155048 199718 155060
rect 271046 155048 271052 155060
rect 271104 155048 271110 155100
rect 200114 155020 200120 155032
rect 195946 154992 200120 155020
rect 200114 154980 200120 154992
rect 200172 154980 200178 155032
rect 207106 154980 207112 155032
rect 207164 155020 207170 155032
rect 269206 155020 269212 155032
rect 207164 154992 269212 155020
rect 207164 154980 207170 154992
rect 269206 154980 269212 154992
rect 269264 154980 269270 155032
rect 15470 154912 15476 154964
rect 15528 154952 15534 154964
rect 109034 154952 109040 154964
rect 15528 154924 109040 154952
rect 15528 154912 15534 154924
rect 109034 154912 109040 154924
rect 109092 154912 109098 154964
rect 110506 154912 110512 154964
rect 110564 154952 110570 154964
rect 139302 154952 139308 154964
rect 110564 154924 139308 154952
rect 110564 154912 110570 154924
rect 139302 154912 139308 154924
rect 139360 154912 139366 154964
rect 145926 154912 145932 154964
rect 145984 154952 145990 154964
rect 230014 154952 230020 154964
rect 145984 154924 230020 154952
rect 145984 154912 145990 154924
rect 230014 154912 230020 154924
rect 230072 154912 230078 154964
rect 250162 154912 250168 154964
rect 250220 154952 250226 154964
rect 309502 154952 309508 154964
rect 250220 154924 309508 154952
rect 250220 154912 250226 154924
rect 309502 154912 309508 154924
rect 309560 154912 309566 154964
rect 106366 154844 106372 154896
rect 106424 154884 106430 154896
rect 186590 154884 186596 154896
rect 106424 154856 186596 154884
rect 106424 154844 106430 154856
rect 186590 154844 186596 154856
rect 186648 154844 186654 154896
rect 186682 154844 186688 154896
rect 186740 154884 186746 154896
rect 245930 154884 245936 154896
rect 186740 154856 245936 154884
rect 186740 154844 186746 154856
rect 245930 154844 245936 154856
rect 245988 154844 245994 154896
rect 109126 154776 109132 154828
rect 109184 154816 109190 154828
rect 133046 154816 133052 154828
rect 109184 154788 133052 154816
rect 109184 154776 109190 154788
rect 133046 154776 133052 154788
rect 133104 154776 133110 154828
rect 149238 154776 149244 154828
rect 149296 154816 149302 154828
rect 232498 154816 232504 154828
rect 149296 154788 232504 154816
rect 149296 154776 149302 154788
rect 232498 154776 232504 154788
rect 232556 154776 232562 154828
rect 155954 154708 155960 154760
rect 156012 154748 156018 154760
rect 237650 154748 237656 154760
rect 156012 154720 237656 154748
rect 156012 154708 156018 154720
rect 237650 154708 237656 154720
rect 237708 154708 237714 154760
rect 162670 154640 162676 154692
rect 162728 154680 162734 154692
rect 242894 154680 242900 154692
rect 162728 154652 242900 154680
rect 162728 154640 162734 154652
rect 242894 154640 242900 154652
rect 242952 154640 242958 154692
rect 154482 154572 154488 154624
rect 154540 154612 154546 154624
rect 154540 154584 155080 154612
rect 154540 154572 154546 154584
rect 51626 154504 51632 154556
rect 51684 154544 51690 154556
rect 154942 154544 154948 154556
rect 51684 154516 154948 154544
rect 51684 154504 51690 154516
rect 154942 154504 154948 154516
rect 155000 154504 155006 154556
rect 155052 154544 155080 154584
rect 159358 154572 159364 154624
rect 159416 154612 159422 154624
rect 240226 154612 240232 154624
rect 159416 154584 240232 154612
rect 159416 154572 159422 154584
rect 240226 154572 240232 154584
rect 240284 154572 240290 154624
rect 156414 154544 156420 154556
rect 155052 154516 156420 154544
rect 156414 154504 156420 154516
rect 156472 154504 156478 154556
rect 156598 154504 156604 154556
rect 156656 154544 156662 154556
rect 212718 154544 212724 154556
rect 156656 154516 212724 154544
rect 156656 154504 156662 154516
rect 212718 154504 212724 154516
rect 212776 154504 212782 154556
rect 219342 154504 219348 154556
rect 219400 154544 219406 154556
rect 286226 154544 286232 154556
rect 219400 154516 286232 154544
rect 219400 154504 219406 154516
rect 286226 154504 286232 154516
rect 286284 154504 286290 154556
rect 286318 154504 286324 154556
rect 286376 154544 286382 154556
rect 337194 154544 337200 154556
rect 286376 154516 337200 154544
rect 286376 154504 286382 154516
rect 337194 154504 337200 154516
rect 337252 154504 337258 154556
rect 353662 154504 353668 154556
rect 353720 154544 353726 154556
rect 388622 154544 388628 154556
rect 353720 154516 388628 154544
rect 353720 154504 353726 154516
rect 388622 154504 388628 154516
rect 388680 154504 388686 154556
rect 44910 154436 44916 154488
rect 44968 154476 44974 154488
rect 142522 154476 142528 154488
rect 44968 154448 142528 154476
rect 44968 154436 44974 154448
rect 142522 154436 142528 154448
rect 142580 154436 142586 154488
rect 142614 154436 142620 154488
rect 142672 154476 142678 154488
rect 191006 154476 191012 154488
rect 142672 154448 191012 154476
rect 142672 154436 142678 154448
rect 191006 154436 191012 154448
rect 191064 154436 191070 154488
rect 202414 154476 202420 154488
rect 191116 154448 202420 154476
rect 41598 154368 41604 154420
rect 41656 154408 41662 154420
rect 142798 154408 142804 154420
rect 41656 154380 142804 154408
rect 41656 154368 41662 154380
rect 142798 154368 142804 154380
rect 142856 154368 142862 154420
rect 142890 154368 142896 154420
rect 142948 154408 142954 154420
rect 142948 154380 181208 154408
rect 142948 154368 142954 154380
rect 113818 154300 113824 154352
rect 113876 154340 113882 154352
rect 181070 154340 181076 154352
rect 113876 154312 181076 154340
rect 113876 154300 113882 154312
rect 181070 154300 181076 154312
rect 181128 154300 181134 154352
rect 181180 154340 181208 154380
rect 181438 154368 181444 154420
rect 181496 154408 181502 154420
rect 189534 154408 189540 154420
rect 181496 154380 189540 154408
rect 181496 154368 181502 154380
rect 189534 154368 189540 154380
rect 189592 154368 189598 154420
rect 191116 154340 191144 154448
rect 202414 154436 202420 154448
rect 202472 154436 202478 154488
rect 208946 154436 208952 154488
rect 209004 154476 209010 154488
rect 278130 154476 278136 154488
rect 209004 154448 278136 154476
rect 209004 154436 209010 154448
rect 278130 154436 278136 154448
rect 278188 154436 278194 154488
rect 279970 154436 279976 154488
rect 280028 154476 280034 154488
rect 332134 154476 332140 154488
rect 280028 154448 332140 154476
rect 280028 154436 280034 154448
rect 332134 154436 332140 154448
rect 332192 154436 332198 154488
rect 350258 154436 350264 154488
rect 350316 154476 350322 154488
rect 386046 154476 386052 154488
rect 350316 154448 386052 154476
rect 350316 154436 350322 154448
rect 386046 154436 386052 154448
rect 386104 154436 386110 154488
rect 191190 154368 191196 154420
rect 191248 154408 191254 154420
rect 258258 154408 258264 154420
rect 191248 154380 258264 154408
rect 191248 154368 191254 154380
rect 258258 154368 258264 154380
rect 258316 154368 258322 154420
rect 266170 154368 266176 154420
rect 266228 154408 266234 154420
rect 321830 154408 321836 154420
rect 266228 154380 321836 154408
rect 266228 154368 266234 154380
rect 321830 154368 321836 154380
rect 321888 154368 321894 154420
rect 346854 154368 346860 154420
rect 346912 154408 346918 154420
rect 383654 154408 383660 154420
rect 346912 154380 383660 154408
rect 346912 154368 346918 154380
rect 383654 154368 383660 154380
rect 383712 154368 383718 154420
rect 390646 154368 390652 154420
rect 390704 154408 390710 154420
rect 416866 154408 416872 154420
rect 390704 154380 416872 154408
rect 390704 154368 390710 154380
rect 416866 154368 416872 154380
rect 416924 154368 416930 154420
rect 181180 154312 191144 154340
rect 191374 154300 191380 154352
rect 191432 154340 191438 154352
rect 201770 154340 201776 154352
rect 191432 154312 201776 154340
rect 191432 154300 191438 154312
rect 201770 154300 201776 154312
rect 201828 154300 201834 154352
rect 205542 154300 205548 154352
rect 205600 154340 205606 154352
rect 275554 154340 275560 154352
rect 205600 154312 275560 154340
rect 205600 154300 205606 154312
rect 275554 154300 275560 154312
rect 275612 154300 275618 154352
rect 276198 154300 276204 154352
rect 276256 154340 276262 154352
rect 329834 154340 329840 154352
rect 276256 154312 329840 154340
rect 276256 154300 276262 154312
rect 329834 154300 329840 154312
rect 329892 154300 329898 154352
rect 340138 154300 340144 154352
rect 340196 154340 340202 154352
rect 378318 154340 378324 154352
rect 340196 154312 378324 154340
rect 340196 154300 340202 154312
rect 378318 154300 378324 154312
rect 378376 154300 378382 154352
rect 387610 154300 387616 154352
rect 387668 154340 387674 154352
rect 414290 154340 414296 154352
rect 387668 154312 414296 154340
rect 387668 154300 387674 154312
rect 414290 154300 414296 154312
rect 414348 154300 414354 154352
rect 38470 154232 38476 154284
rect 38528 154272 38534 154284
rect 38528 154244 142752 154272
rect 38528 154232 38534 154244
rect 23934 154164 23940 154216
rect 23992 154204 23998 154216
rect 23992 154176 132816 154204
rect 23992 154164 23998 154176
rect 27246 154096 27252 154148
rect 27304 154136 27310 154148
rect 132586 154136 132592 154148
rect 27304 154108 132592 154136
rect 27304 154096 27310 154108
rect 132586 154096 132592 154108
rect 132644 154096 132650 154148
rect 13814 154028 13820 154080
rect 13872 154068 13878 154080
rect 129182 154068 129188 154080
rect 13872 154040 129188 154068
rect 13872 154028 13878 154040
rect 129182 154028 129188 154040
rect 129240 154028 129246 154080
rect 132788 154068 132816 154176
rect 132862 154164 132868 154216
rect 132920 154204 132926 154216
rect 132920 154176 133092 154204
rect 132920 154164 132926 154176
rect 133064 154136 133092 154176
rect 133138 154164 133144 154216
rect 133196 154204 133202 154216
rect 142614 154204 142620 154216
rect 133196 154176 142620 154204
rect 133196 154164 133202 154176
rect 142614 154164 142620 154176
rect 142672 154164 142678 154216
rect 139486 154136 139492 154148
rect 133064 154108 139492 154136
rect 139486 154096 139492 154108
rect 139544 154096 139550 154148
rect 139578 154096 139584 154148
rect 139636 154136 139642 154148
rect 142338 154136 142344 154148
rect 139636 154108 142344 154136
rect 139636 154096 139642 154108
rect 142338 154096 142344 154108
rect 142396 154096 142402 154148
rect 142724 154136 142752 154244
rect 147674 154232 147680 154284
rect 147732 154272 147738 154284
rect 156598 154272 156604 154284
rect 147732 154244 156604 154272
rect 147732 154232 147738 154244
rect 156598 154232 156604 154244
rect 156656 154232 156662 154284
rect 172790 154232 172796 154284
rect 172848 154272 172854 154284
rect 250530 154272 250536 154284
rect 172848 154244 250536 154272
rect 172848 154232 172854 154244
rect 250530 154232 250536 154244
rect 250588 154232 250594 154284
rect 256050 154232 256056 154284
rect 256108 154272 256114 154284
rect 314102 154272 314108 154284
rect 256108 154244 314108 154272
rect 256108 154232 256114 154244
rect 314102 154232 314108 154244
rect 314160 154232 314166 154284
rect 343542 154232 343548 154284
rect 343600 154272 343606 154284
rect 380894 154272 380900 154284
rect 343600 154244 380900 154272
rect 343600 154232 343606 154244
rect 380894 154232 380900 154244
rect 380952 154232 380958 154284
rect 383930 154232 383936 154284
rect 383988 154272 383994 154284
rect 411714 154272 411720 154284
rect 383988 154244 411720 154272
rect 383988 154232 383994 154244
rect 411714 154232 411720 154244
rect 411772 154232 411778 154284
rect 142798 154164 142804 154216
rect 142856 154204 142862 154216
rect 150434 154204 150440 154216
rect 142856 154176 150440 154204
rect 142856 154164 142862 154176
rect 150434 154164 150440 154176
rect 150492 154164 150498 154216
rect 152550 154164 152556 154216
rect 152608 154204 152614 154216
rect 152608 154176 156644 154204
rect 152608 154164 152614 154176
rect 147490 154136 147496 154148
rect 142724 154108 147496 154136
rect 147490 154096 147496 154108
rect 147548 154096 147554 154148
rect 147582 154096 147588 154148
rect 147640 154136 147646 154148
rect 156322 154136 156328 154148
rect 147640 154108 156328 154136
rect 147640 154096 147646 154108
rect 156322 154096 156328 154108
rect 156380 154096 156386 154148
rect 156616 154136 156644 154176
rect 156782 154164 156788 154216
rect 156840 154204 156846 154216
rect 163222 154204 163228 154216
rect 156840 154176 163228 154204
rect 156840 154164 156846 154176
rect 163222 154164 163228 154176
rect 163280 154164 163286 154216
rect 166074 154164 166080 154216
rect 166132 154204 166138 154216
rect 245654 154204 245660 154216
rect 166132 154176 245660 154204
rect 166132 154164 166138 154176
rect 245654 154164 245660 154176
rect 245712 154164 245718 154216
rect 249702 154164 249708 154216
rect 249760 154204 249766 154216
rect 309226 154204 309232 154216
rect 249760 154176 309232 154204
rect 249760 154164 249766 154176
rect 309226 154164 309232 154176
rect 309284 154164 309290 154216
rect 326706 154164 326712 154216
rect 326764 154204 326770 154216
rect 368014 154204 368020 154216
rect 326764 154176 368020 154204
rect 326764 154164 326770 154176
rect 368014 154164 368020 154176
rect 368072 154164 368078 154216
rect 380802 154164 380808 154216
rect 380860 154204 380866 154216
rect 409230 154204 409236 154216
rect 380860 154176 409236 154204
rect 380860 154164 380866 154176
rect 409230 154164 409236 154176
rect 409288 154164 409294 154216
rect 156616 154108 158208 154136
rect 136910 154068 136916 154080
rect 132788 154040 136916 154068
rect 136910 154028 136916 154040
rect 136968 154028 136974 154080
rect 137370 154028 137376 154080
rect 137428 154068 137434 154080
rect 142890 154068 142896 154080
rect 137428 154040 142896 154068
rect 137428 154028 137434 154040
rect 142890 154028 142896 154040
rect 142948 154028 142954 154080
rect 153194 154068 153200 154080
rect 143000 154040 153200 154068
rect 10410 153960 10416 154012
rect 10468 154000 10474 154012
rect 126606 154000 126612 154012
rect 10468 153972 126612 154000
rect 10468 153960 10474 153972
rect 126606 153960 126612 153972
rect 126664 153960 126670 154012
rect 127618 153960 127624 154012
rect 127676 154000 127682 154012
rect 142430 154000 142436 154012
rect 127676 153972 142436 154000
rect 127676 153960 127682 153972
rect 142430 153960 142436 153972
rect 142488 153960 142494 154012
rect 142522 153960 142528 154012
rect 142580 154000 142586 154012
rect 143000 154000 143028 154040
rect 153194 154028 153200 154040
rect 153252 154028 153258 154080
rect 154942 154028 154948 154080
rect 155000 154068 155006 154080
rect 158070 154068 158076 154080
rect 155000 154040 158076 154068
rect 155000 154028 155006 154040
rect 158070 154028 158076 154040
rect 158128 154028 158134 154080
rect 158180 154068 158208 154108
rect 160186 154096 160192 154148
rect 160244 154136 160250 154148
rect 240962 154136 240968 154148
rect 160244 154108 240968 154136
rect 160244 154096 160250 154108
rect 240962 154096 240968 154108
rect 241020 154096 241026 154148
rect 242618 154096 242624 154148
rect 242676 154136 242682 154148
rect 303798 154136 303804 154148
rect 242676 154108 303804 154136
rect 242676 154096 242682 154108
rect 303798 154096 303804 154108
rect 303856 154096 303862 154148
rect 323302 154096 323308 154148
rect 323360 154136 323366 154148
rect 365714 154136 365720 154148
rect 323360 154108 365720 154136
rect 323360 154096 323366 154108
rect 365714 154096 365720 154108
rect 365772 154096 365778 154148
rect 367094 154096 367100 154148
rect 367152 154136 367158 154148
rect 398834 154136 398840 154148
rect 367152 154108 398840 154136
rect 367152 154096 367158 154108
rect 398834 154096 398840 154108
rect 398892 154096 398898 154148
rect 401594 154096 401600 154148
rect 401652 154136 401658 154148
rect 425330 154136 425336 154148
rect 401652 154108 425336 154136
rect 401652 154096 401658 154108
rect 425330 154096 425336 154108
rect 425388 154096 425394 154148
rect 235166 154068 235172 154080
rect 158180 154040 235172 154068
rect 235166 154028 235172 154040
rect 235224 154028 235230 154080
rect 235902 154028 235908 154080
rect 235960 154068 235966 154080
rect 298738 154068 298744 154080
rect 235960 154040 298744 154068
rect 235960 154028 235966 154040
rect 298738 154028 298744 154040
rect 298796 154028 298802 154080
rect 316586 154028 316592 154080
rect 316644 154068 316650 154080
rect 360378 154068 360384 154080
rect 316644 154040 360384 154068
rect 316644 154028 316650 154040
rect 360378 154028 360384 154040
rect 360436 154028 360442 154080
rect 363690 154028 363696 154080
rect 363748 154068 363754 154080
rect 396350 154068 396356 154080
rect 363748 154040 396356 154068
rect 363748 154028 363754 154040
rect 396350 154028 396356 154040
rect 396408 154028 396414 154080
rect 398190 154028 398196 154080
rect 398248 154068 398254 154080
rect 422662 154068 422668 154080
rect 398248 154040 422668 154068
rect 398248 154028 398254 154040
rect 422662 154028 422668 154040
rect 422720 154028 422726 154080
rect 142580 153972 143028 154000
rect 142580 153960 142586 153972
rect 143074 153960 143080 154012
rect 143132 154000 143138 154012
rect 222930 154000 222936 154012
rect 143132 153972 222936 154000
rect 143132 153960 143138 153972
rect 222930 153960 222936 153972
rect 222988 153960 222994 154012
rect 288434 154000 288440 154012
rect 223040 153972 288440 154000
rect 7098 153892 7104 153944
rect 7156 153932 7162 153944
rect 124214 153932 124220 153944
rect 7156 153904 124220 153932
rect 7156 153892 7162 153904
rect 124214 153892 124220 153904
rect 124272 153892 124278 153944
rect 125502 153892 125508 153944
rect 125560 153932 125566 153944
rect 133138 153932 133144 153944
rect 125560 153904 133144 153932
rect 125560 153892 125566 153904
rect 133138 153892 133144 153904
rect 133196 153892 133202 153944
rect 133230 153892 133236 153944
rect 133288 153932 133294 153944
rect 219710 153932 219716 153944
rect 133288 153904 219716 153932
rect 133288 153892 133294 153904
rect 219710 153892 219716 153904
rect 219768 153892 219774 153944
rect 222378 153892 222384 153944
rect 222436 153932 222442 153944
rect 223040 153932 223068 153972
rect 288434 153960 288440 153972
rect 288492 153960 288498 154012
rect 313274 153960 313280 154012
rect 313332 154000 313338 154012
rect 357802 154000 357808 154012
rect 313332 153972 357808 154000
rect 313332 153960 313338 153972
rect 357802 153960 357808 153972
rect 357860 153960 357866 154012
rect 360470 153960 360476 154012
rect 360528 154000 360534 154012
rect 393774 154000 393780 154012
rect 360528 153972 393780 154000
rect 360528 153960 360534 153972
rect 393774 153960 393780 153972
rect 393832 153960 393838 154012
rect 397362 153960 397368 154012
rect 397420 154000 397426 154012
rect 422294 154000 422300 154012
rect 397420 153972 422300 154000
rect 397420 153960 397426 153972
rect 422294 153960 422300 153972
rect 422352 153960 422358 154012
rect 222436 153904 223068 153932
rect 222436 153892 222442 153904
rect 225782 153892 225788 153944
rect 225840 153932 225846 153944
rect 291194 153932 291200 153944
rect 225840 153904 291200 153932
rect 225840 153892 225846 153904
rect 291194 153892 291200 153904
rect 291252 153892 291258 153944
rect 309870 153892 309876 153944
rect 309928 153932 309934 153944
rect 355226 153932 355232 153944
rect 309928 153904 355232 153932
rect 309928 153892 309934 153904
rect 355226 153892 355232 153904
rect 355284 153892 355290 153944
rect 357342 153892 357348 153944
rect 357400 153932 357406 153944
rect 391198 153932 391204 153944
rect 357400 153904 391204 153932
rect 357400 153892 357406 153904
rect 391198 153892 391204 153904
rect 391256 153892 391262 153944
rect 393958 153892 393964 153944
rect 394016 153932 394022 153944
rect 419534 153932 419540 153944
rect 394016 153904 419540 153932
rect 394016 153892 394022 153904
rect 419534 153892 419540 153904
rect 419592 153892 419598 153944
rect 1210 153824 1216 153876
rect 1268 153864 1274 153876
rect 119522 153864 119528 153876
rect 1268 153836 119528 153864
rect 1268 153824 1274 153836
rect 119522 153824 119528 153836
rect 119580 153824 119586 153876
rect 119614 153824 119620 153876
rect 119672 153864 119678 153876
rect 209774 153864 209780 153876
rect 119672 153836 209780 153864
rect 119672 153824 119678 153836
rect 209774 153824 209780 153836
rect 209832 153824 209838 153876
rect 215662 153824 215668 153876
rect 215720 153864 215726 153876
rect 283282 153864 283288 153876
rect 215720 153836 283288 153864
rect 215720 153824 215726 153836
rect 283282 153824 283288 153836
rect 283340 153824 283346 153876
rect 283374 153824 283380 153876
rect 283432 153864 283438 153876
rect 334618 153864 334624 153876
rect 283432 153836 334624 153864
rect 283432 153824 283438 153836
rect 334618 153824 334624 153836
rect 334676 153824 334682 153876
rect 336826 153824 336832 153876
rect 336884 153864 336890 153876
rect 375742 153864 375748 153876
rect 336884 153836 375748 153864
rect 336884 153824 336890 153836
rect 375742 153824 375748 153836
rect 375800 153824 375806 153876
rect 377214 153824 377220 153876
rect 377272 153864 377278 153876
rect 406562 153864 406568 153876
rect 377272 153836 406568 153864
rect 377272 153824 377278 153836
rect 406562 153824 406568 153836
rect 406620 153824 406626 153876
rect 48314 153756 48320 153808
rect 48372 153796 48378 153808
rect 155494 153796 155500 153808
rect 48372 153768 155500 153796
rect 48372 153756 48378 153768
rect 155494 153756 155500 153768
rect 155552 153756 155558 153808
rect 156414 153756 156420 153808
rect 156472 153796 156478 153808
rect 218054 153796 218060 153808
rect 156472 153768 218060 153796
rect 156472 153756 156478 153768
rect 218054 153756 218060 153768
rect 218112 153756 218118 153808
rect 232590 153756 232596 153808
rect 232648 153796 232654 153808
rect 296162 153796 296168 153808
rect 232648 153768 296168 153796
rect 232648 153756 232654 153768
rect 296162 153756 296168 153768
rect 296220 153756 296226 153808
rect 435174 153756 435180 153808
rect 435232 153796 435238 153808
rect 442902 153796 442908 153808
rect 435232 153768 442908 153796
rect 435232 153756 435238 153768
rect 442902 153756 442908 153768
rect 442960 153756 442966 153808
rect 61746 153688 61752 153740
rect 61804 153728 61810 153740
rect 165798 153728 165804 153740
rect 61804 153700 165804 153728
rect 61804 153688 61810 153700
rect 165798 153688 165804 153700
rect 165856 153688 165862 153740
rect 210142 153728 210148 153740
rect 171106 153700 210148 153728
rect 58342 153620 58348 153672
rect 58400 153660 58406 153672
rect 156506 153660 156512 153672
rect 58400 153632 156512 153660
rect 58400 153620 58406 153632
rect 156506 153620 156512 153632
rect 156564 153620 156570 153672
rect 156598 153620 156604 153672
rect 156656 153660 156662 153672
rect 171106 153660 171134 153700
rect 210142 153688 210148 153700
rect 210200 153688 210206 153740
rect 229094 153688 229100 153740
rect 229152 153728 229158 153740
rect 293586 153728 293592 153740
rect 229152 153700 293592 153728
rect 229152 153688 229158 153700
rect 293586 153688 293592 153700
rect 293644 153688 293650 153740
rect 156656 153632 171134 153660
rect 156656 153620 156662 153632
rect 176654 153620 176660 153672
rect 176712 153660 176718 153672
rect 176712 153632 179552 153660
rect 176712 153620 176718 153632
rect 79410 153552 79416 153604
rect 79468 153592 79474 153604
rect 179414 153592 179420 153604
rect 79468 153564 179420 153592
rect 79468 153552 79474 153564
rect 179414 153552 179420 153564
rect 179472 153552 179478 153604
rect 179524 153592 179552 153632
rect 182910 153620 182916 153672
rect 182968 153660 182974 153672
rect 191190 153660 191196 153672
rect 182968 153632 191196 153660
rect 182968 153620 182974 153632
rect 191190 153620 191196 153632
rect 191248 153620 191254 153672
rect 191282 153620 191288 153672
rect 191340 153660 191346 153672
rect 195974 153660 195980 153672
rect 191340 153632 195980 153660
rect 191340 153620 191346 153632
rect 195974 153620 195980 153632
rect 196032 153620 196038 153672
rect 196066 153620 196072 153672
rect 196124 153660 196130 153672
rect 238386 153660 238392 153672
rect 196124 153632 238392 153660
rect 196124 153620 196130 153632
rect 238386 153620 238392 153632
rect 238444 153620 238450 153672
rect 239214 153620 239220 153672
rect 239272 153660 239278 153672
rect 301314 153660 301320 153672
rect 239272 153632 301320 153660
rect 239272 153620 239278 153632
rect 301314 153620 301320 153632
rect 301372 153620 301378 153672
rect 230658 153592 230664 153604
rect 179524 153564 230664 153592
rect 230658 153552 230664 153564
rect 230716 153552 230722 153604
rect 246022 153552 246028 153604
rect 246080 153592 246086 153604
rect 306374 153592 306380 153604
rect 246080 153564 306380 153592
rect 246080 153552 246086 153564
rect 306374 153552 306380 153564
rect 306432 153552 306438 153604
rect 102134 153484 102140 153536
rect 102192 153524 102198 153536
rect 196618 153524 196624 153536
rect 102192 153496 196624 153524
rect 102192 153484 102198 153496
rect 196618 153484 196624 153496
rect 196676 153484 196682 153536
rect 196710 153484 196716 153536
rect 196768 153524 196774 153536
rect 196768 153496 197400 153524
rect 196768 153484 196774 153496
rect 105446 153416 105452 153468
rect 105504 153456 105510 153468
rect 197262 153456 197268 153468
rect 105504 153428 197268 153456
rect 105504 153416 105510 153428
rect 197262 153416 197268 153428
rect 197320 153416 197326 153468
rect 197372 153456 197400 153496
rect 200482 153484 200488 153536
rect 200540 153524 200546 153536
rect 258902 153524 258908 153536
rect 200540 153496 258908 153524
rect 200540 153484 200546 153496
rect 258902 153484 258908 153496
rect 258960 153484 258966 153536
rect 262766 153484 262772 153536
rect 262824 153524 262830 153536
rect 319254 153524 319260 153536
rect 262824 153496 319260 153524
rect 262824 153484 262830 153496
rect 319254 153484 319260 153496
rect 319312 153484 319318 153536
rect 197372 153428 197492 153456
rect 108850 153348 108856 153400
rect 108908 153388 108914 153400
rect 191374 153388 191380 153400
rect 108908 153360 191380 153388
rect 108908 153348 108914 153360
rect 191374 153348 191380 153360
rect 191432 153348 191438 153400
rect 191742 153348 191748 153400
rect 191800 153388 191806 153400
rect 195882 153388 195888 153400
rect 191800 153360 195888 153388
rect 191800 153348 191806 153360
rect 195882 153348 195888 153360
rect 195940 153348 195946 153400
rect 195974 153348 195980 153400
rect 196032 153388 196038 153400
rect 197354 153388 197360 153400
rect 196032 153360 197360 153388
rect 196032 153348 196038 153360
rect 197354 153348 197360 153360
rect 197412 153348 197418 153400
rect 197464 153388 197492 153428
rect 197630 153416 197636 153468
rect 197688 153456 197694 153468
rect 199194 153456 199200 153468
rect 197688 153428 199200 153456
rect 197688 153416 197694 153428
rect 199194 153416 199200 153428
rect 199252 153416 199258 153468
rect 199286 153416 199292 153468
rect 199344 153456 199350 153468
rect 248598 153456 248604 153468
rect 199344 153428 248604 153456
rect 199344 153416 199350 153428
rect 248598 153416 248604 153428
rect 248656 153416 248662 153468
rect 252646 153416 252652 153468
rect 252704 153456 252710 153468
rect 311526 153456 311532 153468
rect 252704 153428 311532 153456
rect 252704 153416 252710 153428
rect 311526 153416 311532 153428
rect 311584 153416 311590 153468
rect 243446 153388 243452 153400
rect 197464 153360 243452 153388
rect 243446 153348 243452 153360
rect 243504 153348 243510 153400
rect 259454 153348 259460 153400
rect 259512 153388 259518 153400
rect 316770 153388 316776 153400
rect 259512 153360 316776 153388
rect 259512 153348 259518 153360
rect 316770 153348 316776 153360
rect 316828 153348 316834 153400
rect 116394 153280 116400 153332
rect 116452 153320 116458 153332
rect 207566 153320 207572 153332
rect 116452 153292 207572 153320
rect 116452 153280 116458 153292
rect 207566 153280 207572 153292
rect 207624 153280 207630 153332
rect 272886 153280 272892 153332
rect 272944 153320 272950 153332
rect 327074 153320 327080 153332
rect 272944 153292 327080 153320
rect 272944 153280 272950 153292
rect 327074 153280 327080 153292
rect 327132 153280 327138 153332
rect 34790 153212 34796 153264
rect 34848 153252 34854 153264
rect 142338 153252 142344 153264
rect 34848 153224 142344 153252
rect 34848 153212 34854 153224
rect 142338 153212 142344 153224
rect 142396 153212 142402 153264
rect 142430 153212 142436 153264
rect 142488 153252 142494 153264
rect 204990 153252 204996 153264
rect 142488 153224 204996 153252
rect 142488 153212 142494 153224
rect 204990 153212 204996 153224
rect 205048 153212 205054 153264
rect 269482 153212 269488 153264
rect 269540 153252 269546 153264
rect 324406 153252 324412 153264
rect 269540 153224 324412 153252
rect 269540 153212 269546 153224
rect 324406 153212 324412 153224
rect 324464 153212 324470 153264
rect 66714 153144 66720 153196
rect 66772 153184 66778 153196
rect 159358 153184 159364 153196
rect 66772 153156 159364 153184
rect 66772 153144 66778 153156
rect 159358 153144 159364 153156
rect 159416 153144 159422 153196
rect 172514 153144 172520 153196
rect 172572 153184 172578 153196
rect 249242 153184 249248 153196
rect 172572 153156 249248 153184
rect 172572 153144 172578 153156
rect 249242 153144 249248 153156
rect 249300 153144 249306 153196
rect 255314 153144 255320 153196
rect 255372 153184 255378 153196
rect 312814 153184 312820 153196
rect 255372 153156 312820 153184
rect 255372 153144 255378 153156
rect 312814 153144 312820 153156
rect 312872 153144 312878 153196
rect 316954 153144 316960 153196
rect 317012 153184 317018 153196
rect 317966 153184 317972 153196
rect 317012 153156 317972 153184
rect 317012 153144 317018 153156
rect 317966 153144 317972 153156
rect 318024 153144 318030 153196
rect 318610 153144 318616 153196
rect 318668 153184 318674 153196
rect 318668 153156 320588 153184
rect 318668 153144 318674 153156
rect 30190 153076 30196 153128
rect 30248 153116 30254 153128
rect 109586 153116 109592 153128
rect 30248 153088 109592 153116
rect 30248 153076 30254 153088
rect 109586 153076 109592 153088
rect 109644 153076 109650 153128
rect 109862 153076 109868 153128
rect 109920 153116 109926 153128
rect 197906 153116 197912 153128
rect 109920 153088 197912 153116
rect 109920 153076 109926 153088
rect 197906 153076 197912 153088
rect 197964 153076 197970 153128
rect 203702 153076 203708 153128
rect 203760 153116 203766 153128
rect 266906 153116 266912 153128
rect 203760 153088 266912 153116
rect 203760 153076 203766 153088
rect 266906 153076 266912 153088
rect 266964 153076 266970 153128
rect 267090 153076 267096 153128
rect 267148 153116 267154 153128
rect 320450 153116 320456 153128
rect 267148 153088 320456 153116
rect 267148 153076 267154 153088
rect 320450 153076 320456 153088
rect 320508 153076 320514 153128
rect 320560 153116 320588 153156
rect 320634 153144 320640 153196
rect 320692 153184 320698 153196
rect 361022 153184 361028 153196
rect 320692 153156 361028 153184
rect 320692 153144 320698 153156
rect 361022 153144 361028 153156
rect 361080 153144 361086 153196
rect 366266 153144 366272 153196
rect 366324 153184 366330 153196
rect 366324 153156 366864 153184
rect 366324 153144 366330 153156
rect 320560 153088 320772 153116
rect 80054 153008 80060 153060
rect 80112 153048 80118 153060
rect 174814 153048 174820 153060
rect 80112 153020 174820 153048
rect 80112 153008 80118 153020
rect 174814 153008 174820 153020
rect 174872 153008 174878 153060
rect 174906 153008 174912 153060
rect 174964 153048 174970 153060
rect 251818 153048 251824 153060
rect 174964 153020 251824 153048
rect 174964 153008 174970 153020
rect 251818 153008 251824 153020
rect 251876 153008 251882 153060
rect 257706 153008 257712 153060
rect 257764 153048 257770 153060
rect 315390 153048 315396 153060
rect 257764 153020 315396 153048
rect 257764 153008 257770 153020
rect 315390 153008 315396 153020
rect 315448 153008 315454 153060
rect 317414 153008 317420 153060
rect 317472 153048 317478 153060
rect 320634 153048 320640 153060
rect 317472 153020 320640 153048
rect 317472 153008 317478 153020
rect 320634 153008 320640 153020
rect 320692 153008 320698 153060
rect 320744 153048 320772 153088
rect 325050 153076 325056 153128
rect 325108 153116 325114 153128
rect 366726 153116 366732 153128
rect 325108 153088 366732 153116
rect 325108 153076 325114 153088
rect 366726 153076 366732 153088
rect 366784 153076 366790 153128
rect 366836 153116 366864 153156
rect 367186 153144 367192 153196
rect 367244 153184 367250 153196
rect 368658 153184 368664 153196
rect 367244 153156 368664 153184
rect 367244 153144 367250 153156
rect 368658 153144 368664 153156
rect 368716 153144 368722 153196
rect 371326 153144 371332 153196
rect 371384 153184 371390 153196
rect 402054 153184 402060 153196
rect 371384 153156 402060 153184
rect 371384 153144 371390 153156
rect 402054 153144 402060 153156
rect 402112 153144 402118 153196
rect 407850 153184 407856 153196
rect 402946 153156 407856 153184
rect 397914 153116 397920 153128
rect 366836 153088 397920 153116
rect 397914 153076 397920 153088
rect 397972 153076 397978 153128
rect 398098 153076 398104 153128
rect 398156 153116 398162 153128
rect 402946 153116 402974 153156
rect 407850 153144 407856 153156
rect 407908 153144 407914 153196
rect 415302 153144 415308 153196
rect 415360 153184 415366 153196
rect 435450 153184 435456 153196
rect 415360 153156 435456 153184
rect 415360 153144 415366 153156
rect 435450 153144 435456 153156
rect 435508 153144 435514 153196
rect 437750 153144 437756 153196
rect 437808 153184 437814 153196
rect 452838 153184 452844 153196
rect 437808 153156 452844 153184
rect 437808 153144 437814 153156
rect 452838 153144 452844 153156
rect 452896 153144 452902 153196
rect 456794 153144 456800 153196
rect 456852 153184 456858 153196
rect 459186 153184 459192 153196
rect 456852 153156 459192 153184
rect 456852 153144 456858 153156
rect 459186 153144 459192 153156
rect 459244 153144 459250 153196
rect 461854 153144 461860 153196
rect 461912 153184 461918 153196
rect 463050 153184 463056 153196
rect 461912 153156 463056 153184
rect 461912 153144 461918 153156
rect 463050 153144 463056 153156
rect 463108 153144 463114 153196
rect 466454 153144 466460 153196
rect 466512 153184 466518 153196
rect 469490 153184 469496 153196
rect 466512 153156 469496 153184
rect 466512 153144 466518 153156
rect 469490 153144 469496 153156
rect 469548 153144 469554 153196
rect 471238 153144 471244 153196
rect 471296 153184 471302 153196
rect 473538 153184 473544 153196
rect 471296 153156 473544 153184
rect 471296 153144 471302 153156
rect 473538 153144 473544 153156
rect 473596 153144 473602 153196
rect 474826 153144 474832 153196
rect 474884 153184 474890 153196
rect 476574 153184 476580 153196
rect 474884 153156 476580 153184
rect 474884 153144 474890 153156
rect 476574 153144 476580 153156
rect 476632 153144 476638 153196
rect 485682 153144 485688 153196
rect 485740 153184 485746 153196
rect 489362 153184 489368 153196
rect 485740 153156 489368 153184
rect 485740 153144 485746 153156
rect 489362 153144 489368 153156
rect 489420 153144 489426 153196
rect 492398 153144 492404 153196
rect 492456 153184 492462 153196
rect 494514 153184 494520 153196
rect 492456 153156 494520 153184
rect 492456 153144 492462 153156
rect 494514 153144 494520 153156
rect 494572 153144 494578 153196
rect 495250 153144 495256 153196
rect 495308 153184 495314 153196
rect 496446 153184 496452 153196
rect 495308 153156 496452 153184
rect 495308 153144 495314 153156
rect 496446 153144 496452 153156
rect 496504 153144 496510 153196
rect 496630 153144 496636 153196
rect 496688 153184 496694 153196
rect 497734 153184 497740 153196
rect 496688 153156 497740 153184
rect 496688 153144 496694 153156
rect 497734 153144 497740 153156
rect 497792 153144 497798 153196
rect 498286 153144 498292 153196
rect 498344 153184 498350 153196
rect 499022 153184 499028 153196
rect 498344 153156 499028 153184
rect 498344 153144 498350 153156
rect 499022 153144 499028 153156
rect 499080 153144 499086 153196
rect 500954 153144 500960 153196
rect 501012 153184 501018 153196
rect 501598 153184 501604 153196
rect 501012 153156 501604 153184
rect 501012 153144 501018 153156
rect 501598 153144 501604 153156
rect 501656 153144 501662 153196
rect 510430 153144 510436 153196
rect 510488 153184 510494 153196
rect 511994 153184 512000 153196
rect 510488 153156 512000 153184
rect 510488 153144 510494 153156
rect 511994 153144 512000 153156
rect 512052 153144 512058 153196
rect 512546 153144 512552 153196
rect 512604 153184 512610 153196
rect 514846 153184 514852 153196
rect 512604 153156 514852 153184
rect 512604 153144 512610 153156
rect 514846 153144 514852 153156
rect 514904 153144 514910 153196
rect 398156 153088 402974 153116
rect 398156 153076 398162 153088
rect 405826 153076 405832 153128
rect 405884 153116 405890 153128
rect 408494 153116 408500 153128
rect 405884 153088 408500 153116
rect 405884 153076 405890 153088
rect 408494 153076 408500 153088
rect 408552 153076 408558 153128
rect 411622 153076 411628 153128
rect 411680 153116 411686 153128
rect 411680 153088 431954 153116
rect 411680 153076 411686 153088
rect 361666 153048 361672 153060
rect 320744 153020 361672 153048
rect 361666 153008 361672 153020
rect 361724 153008 361730 153060
rect 364518 153008 364524 153060
rect 364576 153048 364582 153060
rect 396902 153048 396908 153060
rect 364576 153020 396908 153048
rect 364576 153008 364582 153020
rect 396902 153008 396908 153020
rect 396960 153008 396966 153060
rect 407022 153008 407028 153060
rect 407080 153048 407086 153060
rect 429194 153048 429200 153060
rect 407080 153020 429200 153048
rect 407080 153008 407086 153020
rect 429194 153008 429200 153020
rect 429252 153008 429258 153060
rect 431926 153048 431954 153088
rect 432690 153076 432696 153128
rect 432748 153116 432754 153128
rect 448974 153116 448980 153128
rect 432748 153088 448980 153116
rect 432748 153076 432754 153088
rect 448974 153076 448980 153088
rect 449032 153076 449038 153128
rect 466546 153076 466552 153128
rect 466604 153116 466610 153128
rect 470134 153116 470140 153128
rect 466604 153088 470140 153116
rect 466604 153076 466610 153088
rect 470134 153076 470140 153088
rect 470192 153076 470198 153128
rect 471698 153076 471704 153128
rect 471756 153116 471762 153128
rect 472710 153116 472716 153128
rect 471756 153088 472716 153116
rect 471756 153076 471762 153088
rect 472710 153076 472716 153088
rect 472768 153076 472774 153128
rect 473354 153076 473360 153128
rect 473412 153116 473418 153128
rect 475286 153116 475292 153128
rect 473412 153088 475292 153116
rect 473412 153076 473418 153088
rect 475286 153076 475292 153088
rect 475344 153076 475350 153128
rect 476114 153076 476120 153128
rect 476172 153116 476178 153128
rect 477862 153116 477868 153128
rect 476172 153088 477868 153116
rect 476172 153076 476178 153088
rect 477862 153076 477868 153088
rect 477920 153076 477926 153128
rect 484302 153076 484308 153128
rect 484360 153116 484366 153128
rect 488166 153116 488172 153128
rect 484360 153088 488172 153116
rect 484360 153076 484366 153088
rect 488166 153076 488172 153088
rect 488224 153076 488230 153128
rect 489914 153076 489920 153128
rect 489972 153116 489978 153128
rect 492766 153116 492772 153128
rect 489972 153088 492772 153116
rect 489972 153076 489978 153088
rect 492766 153076 492772 153088
rect 492824 153076 492830 153128
rect 493226 153076 493232 153128
rect 493284 153116 493290 153128
rect 495434 153116 495440 153128
rect 493284 153088 495440 153116
rect 493284 153076 493290 153088
rect 495434 153076 495440 153088
rect 495492 153076 495498 153128
rect 495802 153076 495808 153128
rect 495860 153116 495866 153128
rect 497090 153116 497096 153128
rect 495860 153088 497096 153116
rect 495860 153076 495866 153088
rect 497090 153076 497096 153088
rect 497148 153076 497154 153128
rect 511258 153076 511264 153128
rect 511316 153116 511322 153128
rect 513466 153116 513472 153128
rect 511316 153088 513472 153116
rect 511316 153076 511322 153088
rect 513466 153076 513472 153088
rect 513524 153076 513530 153128
rect 432874 153048 432880 153060
rect 431926 153020 432880 153048
rect 432874 153008 432880 153020
rect 432932 153008 432938 153060
rect 433518 153008 433524 153060
rect 433576 153048 433582 153060
rect 449894 153048 449900 153060
rect 433576 153020 449900 153048
rect 433576 153008 433582 153020
rect 449894 153008 449900 153020
rect 449952 153008 449958 153060
rect 465074 153008 465080 153060
rect 465132 153048 465138 153060
rect 468846 153048 468852 153060
rect 465132 153020 468852 153048
rect 465132 153008 465138 153020
rect 468846 153008 468852 153020
rect 468904 153008 468910 153060
rect 472250 153008 472256 153060
rect 472308 153048 472314 153060
rect 473998 153048 474004 153060
rect 472308 153020 474004 153048
rect 472308 153008 472314 153020
rect 473998 153008 474004 153020
rect 474056 153008 474062 153060
rect 484854 153008 484860 153060
rect 484912 153048 484918 153060
rect 488718 153048 488724 153060
rect 484912 153020 488724 153048
rect 484912 153008 484918 153020
rect 488718 153008 488724 153020
rect 488776 153008 488782 153060
rect 497458 153008 497464 153060
rect 497516 153048 497522 153060
rect 498286 153048 498292 153060
rect 497516 153020 498292 153048
rect 497516 153008 497522 153020
rect 498286 153008 498292 153020
rect 498344 153008 498350 153060
rect 511718 153008 511724 153060
rect 511776 153048 511782 153060
rect 514294 153048 514300 153060
rect 511776 153020 514300 153048
rect 511776 153008 511782 153020
rect 514294 153008 514300 153020
rect 514352 153008 514358 153060
rect 97074 152940 97080 152992
rect 97132 152980 97138 152992
rect 192754 152980 192760 152992
rect 97132 152952 192760 152980
rect 97132 152940 97138 152952
rect 192754 152940 192760 152952
rect 192812 152940 192818 152992
rect 194962 152940 194968 152992
rect 195020 152980 195026 152992
rect 218422 152980 218428 152992
rect 195020 152952 218428 152980
rect 195020 152940 195026 152952
rect 218422 152940 218428 152952
rect 218480 152940 218486 152992
rect 225138 152940 225144 152992
rect 225196 152980 225202 152992
rect 228726 152980 228732 152992
rect 225196 152952 228732 152980
rect 225196 152940 225202 152952
rect 228726 152940 228732 152952
rect 228784 152940 228790 152992
rect 228818 152940 228824 152992
rect 228876 152980 228882 152992
rect 284570 152980 284576 152992
rect 228876 152952 284576 152980
rect 228876 152940 228882 152952
rect 284570 152940 284576 152952
rect 284628 152940 284634 152992
rect 285490 152940 285496 152992
rect 285548 152980 285554 152992
rect 336734 152980 336740 152992
rect 285548 152952 336740 152980
rect 285548 152940 285554 152952
rect 336734 152940 336740 152952
rect 336792 152940 336798 152992
rect 339494 152940 339500 152992
rect 339552 152980 339558 152992
rect 377030 152980 377036 152992
rect 339552 152952 377036 152980
rect 339552 152940 339558 152952
rect 377030 152940 377036 152952
rect 377088 152940 377094 152992
rect 382182 152940 382188 152992
rect 382240 152980 382246 152992
rect 410426 152980 410432 152992
rect 382240 152952 410432 152980
rect 382240 152940 382246 152952
rect 410426 152940 410432 152952
rect 410484 152940 410490 152992
rect 410886 152940 410892 152992
rect 410944 152980 410950 152992
rect 430942 152980 430948 152992
rect 410944 152952 430948 152980
rect 410944 152940 410950 152952
rect 430942 152940 430948 152952
rect 431000 152940 431006 152992
rect 431034 152940 431040 152992
rect 431092 152980 431098 152992
rect 447686 152980 447692 152992
rect 431092 152952 447692 152980
rect 431092 152940 431098 152952
rect 447686 152940 447692 152952
rect 447744 152940 447750 152992
rect 472342 152940 472348 152992
rect 472400 152980 472406 152992
rect 474734 152980 474740 152992
rect 472400 152952 474740 152980
rect 472400 152940 472406 152952
rect 474734 152940 474740 152952
rect 474792 152940 474798 152992
rect 483198 152940 483204 152992
rect 483256 152980 483262 152992
rect 487522 152980 487528 152992
rect 483256 152952 487528 152980
rect 483256 152940 483262 152952
rect 487522 152940 487528 152952
rect 487580 152940 487586 152992
rect 490742 152940 490748 152992
rect 490800 152980 490806 152992
rect 493226 152980 493232 152992
rect 490800 152952 493232 152980
rect 490800 152940 490806 152952
rect 493226 152940 493232 152952
rect 493284 152940 493290 152992
rect 494054 152940 494060 152992
rect 494112 152980 494118 152992
rect 495802 152980 495808 152992
rect 494112 152952 495808 152980
rect 494112 152940 494118 152952
rect 495802 152940 495808 152952
rect 495860 152940 495866 152992
rect 502886 152940 502892 152992
rect 502944 152980 502950 152992
rect 503346 152980 503352 152992
rect 502944 152952 503352 152980
rect 502944 152940 502950 152952
rect 503346 152940 503352 152952
rect 503404 152940 503410 152992
rect 513190 152940 513196 152992
rect 513248 152980 513254 152992
rect 515950 152980 515956 152992
rect 513248 152952 515956 152980
rect 513248 152940 513254 152952
rect 515950 152940 515956 152952
rect 516008 152940 516014 152992
rect 92474 152872 92480 152924
rect 92532 152912 92538 152924
rect 187694 152912 187700 152924
rect 92532 152884 187700 152912
rect 92532 152872 92538 152884
rect 187694 152872 187700 152884
rect 187752 152872 187758 152924
rect 187878 152872 187884 152924
rect 187936 152912 187942 152924
rect 262214 152912 262220 152924
rect 187936 152884 262220 152912
rect 187936 152872 187942 152884
rect 262214 152872 262220 152884
rect 262272 152872 262278 152924
rect 265342 152872 265348 152924
rect 265400 152912 265406 152924
rect 321186 152912 321192 152924
rect 265400 152884 321192 152912
rect 265400 152872 265406 152884
rect 321186 152872 321192 152884
rect 321244 152872 321250 152924
rect 324222 152872 324228 152924
rect 324280 152912 324286 152924
rect 366082 152912 366088 152924
rect 324280 152884 366088 152912
rect 324280 152872 324286 152884
rect 366082 152872 366088 152884
rect 366140 152872 366146 152924
rect 368750 152872 368756 152924
rect 368808 152912 368814 152924
rect 400214 152912 400220 152924
rect 368808 152884 400220 152912
rect 368808 152872 368814 152884
rect 400214 152872 400220 152884
rect 400272 152872 400278 152924
rect 402422 152872 402428 152924
rect 402480 152912 402486 152924
rect 425882 152912 425888 152924
rect 402480 152884 425888 152912
rect 402480 152872 402486 152884
rect 425882 152872 425888 152884
rect 425940 152872 425946 152924
rect 428458 152872 428464 152924
rect 428516 152912 428522 152924
rect 439498 152912 439504 152924
rect 428516 152884 439504 152912
rect 428516 152872 428522 152884
rect 439498 152872 439504 152884
rect 439556 152872 439562 152924
rect 440234 152872 440240 152924
rect 440292 152912 440298 152924
rect 441522 152912 441528 152924
rect 440292 152884 441528 152912
rect 440292 152872 440298 152884
rect 441522 152872 441528 152884
rect 441580 152872 441586 152924
rect 441982 152872 441988 152924
rect 442040 152912 442046 152924
rect 442718 152912 442724 152924
rect 442040 152884 442724 152912
rect 442040 152872 442046 152884
rect 442718 152872 442724 152884
rect 442776 152872 442782 152924
rect 442994 152872 443000 152924
rect 443052 152912 443058 152924
rect 445754 152912 445760 152924
rect 443052 152884 445760 152912
rect 443052 152872 443058 152884
rect 445754 152872 445760 152884
rect 445812 152872 445818 152924
rect 446950 152872 446956 152924
rect 447008 152912 447014 152924
rect 459830 152912 459836 152924
rect 447008 152884 459836 152912
rect 447008 152872 447014 152884
rect 459830 152872 459836 152884
rect 459888 152872 459894 152924
rect 513834 152872 513840 152924
rect 513892 152912 513898 152924
rect 516134 152912 516140 152924
rect 513892 152884 516140 152912
rect 513892 152872 513898 152884
rect 516134 152872 516140 152884
rect 516192 152872 516198 152924
rect 33134 152804 33140 152856
rect 33192 152844 33198 152856
rect 143994 152844 144000 152856
rect 33192 152816 144000 152844
rect 33192 152804 33198 152816
rect 143994 152804 144000 152816
rect 144052 152804 144058 152856
rect 144822 152804 144828 152856
rect 144880 152844 144886 152856
rect 161934 152844 161940 152856
rect 144880 152816 161940 152844
rect 144880 152804 144886 152816
rect 161934 152804 161940 152816
rect 161992 152804 161998 152856
rect 164418 152804 164424 152856
rect 164476 152844 164482 152856
rect 244274 152844 244280 152856
rect 164476 152816 244280 152844
rect 164476 152804 164482 152816
rect 244274 152804 244280 152816
rect 244332 152804 244338 152856
rect 251910 152804 251916 152856
rect 251968 152844 251974 152856
rect 310882 152844 310888 152856
rect 251968 152816 310888 152844
rect 251968 152804 251974 152816
rect 310882 152804 310888 152816
rect 310940 152804 310946 152856
rect 311986 152804 311992 152856
rect 312044 152844 312050 152856
rect 356054 152844 356060 152856
rect 312044 152816 356060 152844
rect 312044 152804 312050 152816
rect 356054 152804 356060 152816
rect 356112 152804 356118 152856
rect 362034 152804 362040 152856
rect 362092 152844 362098 152856
rect 395062 152844 395068 152856
rect 362092 152816 395068 152844
rect 362092 152804 362098 152816
rect 395062 152804 395068 152816
rect 395120 152804 395126 152856
rect 395154 152804 395160 152856
rect 395212 152844 395218 152856
rect 397546 152844 397552 152856
rect 395212 152816 397552 152844
rect 395212 152804 395218 152816
rect 397546 152804 397552 152816
rect 397604 152804 397610 152856
rect 400122 152804 400128 152856
rect 400180 152844 400186 152856
rect 423950 152844 423956 152856
rect 400180 152816 423956 152844
rect 400180 152804 400186 152816
rect 423950 152804 423956 152816
rect 424008 152804 424014 152856
rect 426250 152804 426256 152856
rect 426308 152844 426314 152856
rect 443822 152844 443828 152856
rect 426308 152816 443828 152844
rect 426308 152804 426314 152816
rect 443822 152804 443828 152816
rect 443880 152804 443886 152856
rect 445662 152804 445668 152856
rect 445720 152844 445726 152856
rect 458542 152844 458548 152856
rect 445720 152816 458548 152844
rect 445720 152804 445726 152816
rect 458542 152804 458548 152816
rect 458600 152804 458606 152856
rect 491570 152804 491576 152856
rect 491628 152844 491634 152856
rect 494054 152844 494060 152856
rect 491628 152816 494060 152844
rect 491628 152804 491634 152816
rect 494054 152804 494060 152816
rect 494112 152804 494118 152856
rect 26418 152736 26424 152788
rect 26476 152776 26482 152788
rect 138842 152776 138848 152788
rect 26476 152748 138848 152776
rect 26476 152736 26482 152748
rect 138842 152736 138848 152748
rect 138900 152736 138906 152788
rect 142338 152736 142344 152788
rect 142396 152776 142402 152788
rect 145282 152776 145288 152788
rect 142396 152748 145288 152776
rect 142396 152736 142402 152748
rect 145282 152736 145288 152748
rect 145340 152736 145346 152788
rect 149054 152736 149060 152788
rect 149112 152776 149118 152788
rect 231302 152776 231308 152788
rect 149112 152748 231308 152776
rect 149112 152736 149118 152748
rect 231302 152736 231308 152748
rect 231360 152736 231366 152788
rect 245102 152736 245108 152788
rect 245160 152776 245166 152788
rect 305730 152776 305736 152788
rect 245160 152748 305736 152776
rect 245160 152736 245166 152748
rect 305730 152736 305736 152748
rect 305788 152736 305794 152788
rect 307662 152736 307668 152788
rect 307720 152776 307726 152788
rect 352006 152776 352012 152788
rect 307720 152748 352012 152776
rect 307720 152736 307726 152748
rect 352006 152736 352012 152748
rect 352064 152736 352070 152788
rect 352742 152736 352748 152788
rect 352800 152776 352806 152788
rect 387978 152776 387984 152788
rect 352800 152748 387984 152776
rect 352800 152736 352806 152748
rect 387978 152736 387984 152748
rect 388036 152736 388042 152788
rect 390370 152736 390376 152788
rect 390428 152776 390434 152788
rect 414934 152776 414940 152788
rect 390428 152748 414940 152776
rect 390428 152736 390434 152748
rect 414934 152736 414940 152748
rect 414992 152736 414998 152788
rect 415854 152736 415860 152788
rect 415912 152776 415918 152788
rect 436094 152776 436100 152788
rect 415912 152748 436100 152776
rect 415912 152736 415918 152748
rect 436094 152736 436100 152748
rect 436152 152736 436158 152788
rect 437290 152736 437296 152788
rect 437348 152776 437354 152788
rect 452194 152776 452200 152788
rect 437348 152748 442028 152776
rect 437348 152736 437354 152748
rect 28902 152668 28908 152720
rect 28960 152708 28966 152720
rect 140774 152708 140780 152720
rect 28960 152680 140780 152708
rect 28960 152668 28966 152680
rect 140774 152668 140780 152680
rect 140832 152668 140838 152720
rect 140866 152668 140872 152720
rect 140924 152708 140930 152720
rect 140924 152680 142384 152708
rect 140924 152668 140930 152680
rect 22186 152600 22192 152652
rect 22244 152640 22250 152652
rect 135622 152640 135628 152652
rect 22244 152612 135628 152640
rect 22244 152600 22250 152612
rect 135622 152600 135628 152612
rect 135680 152600 135686 152652
rect 137094 152600 137100 152652
rect 137152 152640 137158 152652
rect 142246 152640 142252 152652
rect 137152 152612 142252 152640
rect 137152 152600 137158 152612
rect 142246 152600 142252 152612
rect 142304 152600 142310 152652
rect 142356 152640 142384 152680
rect 143258 152668 143264 152720
rect 143316 152708 143322 152720
rect 156782 152708 156788 152720
rect 143316 152680 156788 152708
rect 143316 152668 143322 152680
rect 156782 152668 156788 152680
rect 156840 152668 156846 152720
rect 172422 152668 172428 152720
rect 172480 152708 172486 152720
rect 176102 152708 176108 152720
rect 172480 152680 176108 152708
rect 172480 152668 172486 152680
rect 176102 152668 176108 152680
rect 176160 152668 176166 152720
rect 220722 152668 220728 152720
rect 220780 152708 220786 152720
rect 228818 152708 228824 152720
rect 220780 152680 228824 152708
rect 220780 152668 220786 152680
rect 228818 152668 228824 152680
rect 228876 152668 228882 152720
rect 247678 152668 247684 152720
rect 247736 152708 247742 152720
rect 307754 152708 307760 152720
rect 247736 152680 307760 152708
rect 247736 152668 247742 152680
rect 307754 152668 307760 152680
rect 307812 152668 307818 152720
rect 311802 152668 311808 152720
rect 311860 152708 311866 152720
rect 356514 152708 356520 152720
rect 311860 152680 356520 152708
rect 311860 152668 311866 152680
rect 356514 152668 356520 152680
rect 356572 152668 356578 152720
rect 359550 152668 359556 152720
rect 359608 152708 359614 152720
rect 393314 152708 393320 152720
rect 359608 152680 393320 152708
rect 359608 152668 359614 152680
rect 393314 152668 393320 152680
rect 393372 152668 393378 152720
rect 394878 152668 394884 152720
rect 394936 152708 394942 152720
rect 420086 152708 420092 152720
rect 394936 152680 420092 152708
rect 394936 152668 394942 152680
rect 420086 152668 420092 152680
rect 420144 152668 420150 152720
rect 423398 152668 423404 152720
rect 423456 152708 423462 152720
rect 441890 152708 441896 152720
rect 423456 152680 441896 152708
rect 423456 152668 423462 152680
rect 441890 152668 441896 152680
rect 441948 152668 441954 152720
rect 442000 152708 442028 152748
rect 444346 152748 452200 152776
rect 444346 152708 444374 152748
rect 452194 152736 452200 152748
rect 452252 152736 452258 152788
rect 442000 152680 444374 152708
rect 444466 152668 444472 152720
rect 444524 152708 444530 152720
rect 458174 152708 458180 152720
rect 444524 152680 458180 152708
rect 444524 152668 444530 152680
rect 458174 152668 458180 152680
rect 458232 152668 458238 152720
rect 226334 152640 226340 152652
rect 142356 152612 226340 152640
rect 226334 152600 226340 152612
rect 226392 152600 226398 152652
rect 234522 152600 234528 152652
rect 234580 152640 234586 152652
rect 297450 152640 297456 152652
rect 234580 152612 297456 152640
rect 234580 152600 234586 152612
rect 297450 152600 297456 152612
rect 297508 152600 297514 152652
rect 304810 152600 304816 152652
rect 304868 152640 304874 152652
rect 351362 152640 351368 152652
rect 304868 152612 351368 152640
rect 304868 152600 304874 152612
rect 351362 152600 351368 152612
rect 351420 152600 351426 152652
rect 354490 152600 354496 152652
rect 354548 152640 354554 152652
rect 389266 152640 389272 152652
rect 354548 152612 389272 152640
rect 354548 152600 354554 152612
rect 389266 152600 389272 152612
rect 389324 152600 389330 152652
rect 393130 152600 393136 152652
rect 393188 152640 393194 152652
rect 418798 152640 418804 152652
rect 393188 152612 418804 152640
rect 393188 152600 393194 152612
rect 418798 152600 418804 152612
rect 418856 152600 418862 152652
rect 419258 152600 419264 152652
rect 419316 152640 419322 152652
rect 438854 152640 438860 152652
rect 419316 152612 438860 152640
rect 419316 152600 419322 152612
rect 438854 152600 438860 152612
rect 438912 152600 438918 152652
rect 442810 152600 442816 152652
rect 442868 152640 442874 152652
rect 456794 152640 456800 152652
rect 442868 152612 456800 152640
rect 442868 152600 442874 152612
rect 456794 152600 456800 152612
rect 456852 152600 456858 152652
rect 19702 152532 19708 152584
rect 19760 152572 19766 152584
rect 133874 152572 133880 152584
rect 19760 152544 133880 152572
rect 19760 152532 19766 152544
rect 133874 152532 133880 152544
rect 133932 152532 133938 152584
rect 134058 152532 134064 152584
rect 134116 152572 134122 152584
rect 220998 152572 221004 152584
rect 134116 152544 221004 152572
rect 134116 152532 134122 152544
rect 220998 152532 221004 152544
rect 221056 152532 221062 152584
rect 228266 152532 228272 152584
rect 228324 152572 228330 152584
rect 292942 152572 292948 152584
rect 228324 152544 292948 152572
rect 228324 152532 228330 152544
rect 292942 152532 292948 152544
rect 293000 152532 293006 152584
rect 299382 152532 299388 152584
rect 299440 152572 299446 152584
rect 346854 152572 346860 152584
rect 299440 152544 346860 152572
rect 299440 152532 299446 152544
rect 346854 152532 346860 152544
rect 346912 152532 346918 152584
rect 349062 152532 349068 152584
rect 349120 152572 349126 152584
rect 385034 152572 385040 152584
rect 349120 152544 385040 152572
rect 349120 152532 349126 152544
rect 385034 152532 385040 152544
rect 385092 152532 385098 152584
rect 386414 152532 386420 152584
rect 386472 152572 386478 152584
rect 413646 152572 413652 152584
rect 386472 152544 413652 152572
rect 386472 152532 386478 152544
rect 413646 152532 413652 152544
rect 413704 152532 413710 152584
rect 413922 152532 413928 152584
rect 413980 152572 413986 152584
rect 433518 152572 433524 152584
rect 413980 152544 433524 152572
rect 413980 152532 413986 152544
rect 433518 152532 433524 152544
rect 433576 152532 433582 152584
rect 434622 152532 434628 152584
rect 434680 152572 434686 152584
rect 450262 152572 450268 152584
rect 434680 152544 450268 152572
rect 434680 152532 434686 152544
rect 450262 152532 450268 152544
rect 450320 152532 450326 152584
rect 2866 152464 2872 152516
rect 2924 152504 2930 152516
rect 120810 152504 120816 152516
rect 2924 152476 120816 152504
rect 2924 152464 2930 152476
rect 120810 152464 120816 152476
rect 120868 152464 120874 152516
rect 210786 152504 210792 152516
rect 120920 152476 210792 152504
rect 23290 152396 23296 152448
rect 23348 152436 23354 152448
rect 110966 152436 110972 152448
rect 23348 152408 110972 152436
rect 23348 152396 23354 152408
rect 110966 152396 110972 152408
rect 111024 152396 111030 152448
rect 120626 152396 120632 152448
rect 120684 152436 120690 152448
rect 120920 152436 120948 152476
rect 210786 152464 210792 152476
rect 210844 152464 210850 152516
rect 212442 152464 212448 152516
rect 212500 152504 212506 152516
rect 277486 152504 277492 152516
rect 212500 152476 277492 152504
rect 212500 152464 212506 152476
rect 277486 152464 277492 152476
rect 277544 152464 277550 152516
rect 278774 152464 278780 152516
rect 278832 152504 278838 152516
rect 278832 152476 279556 152504
rect 278832 152464 278838 152476
rect 120684 152408 120948 152436
rect 120684 152396 120690 152408
rect 120994 152396 121000 152448
rect 121052 152436 121058 152448
rect 205634 152436 205640 152448
rect 121052 152408 205640 152436
rect 121052 152396 121058 152408
rect 205634 152396 205640 152408
rect 205692 152396 205698 152448
rect 215294 152396 215300 152448
rect 215352 152436 215358 152448
rect 279418 152436 279424 152448
rect 215352 152408 279424 152436
rect 215352 152396 215358 152408
rect 279418 152396 279424 152408
rect 279476 152396 279482 152448
rect 279528 152436 279556 152476
rect 279602 152464 279608 152516
rect 279660 152504 279666 152516
rect 330846 152504 330852 152516
rect 279660 152476 330852 152504
rect 279660 152464 279666 152476
rect 330846 152464 330852 152476
rect 330904 152464 330910 152516
rect 330938 152464 330944 152516
rect 330996 152504 331002 152516
rect 371234 152504 371240 152516
rect 330996 152476 371240 152504
rect 330996 152464 331002 152476
rect 371234 152464 371240 152476
rect 371292 152464 371298 152516
rect 372982 152464 372988 152516
rect 373040 152504 373046 152516
rect 403342 152504 403348 152516
rect 373040 152476 403348 152504
rect 373040 152464 373046 152476
rect 403342 152464 403348 152476
rect 403400 152464 403406 152516
rect 404906 152464 404912 152516
rect 404964 152504 404970 152516
rect 427814 152504 427820 152516
rect 404964 152476 427820 152504
rect 404964 152464 404970 152476
rect 427814 152464 427820 152476
rect 427872 152464 427878 152516
rect 430206 152464 430212 152516
rect 430264 152504 430270 152516
rect 447134 152504 447140 152516
rect 430264 152476 447140 152504
rect 430264 152464 430270 152476
rect 447134 152464 447140 152476
rect 447192 152464 447198 152516
rect 331490 152436 331496 152448
rect 279528 152408 331496 152436
rect 331490 152396 331496 152408
rect 331548 152396 331554 152448
rect 332594 152396 332600 152448
rect 332652 152436 332658 152448
rect 372614 152436 372620 152448
rect 332652 152408 372620 152436
rect 332652 152396 332658 152408
rect 372614 152396 372620 152408
rect 372672 152396 372678 152448
rect 375466 152396 375472 152448
rect 375524 152436 375530 152448
rect 405274 152436 405280 152448
rect 375524 152408 405280 152436
rect 375524 152396 375530 152408
rect 405274 152396 405280 152408
rect 405332 152396 405338 152448
rect 408586 152396 408592 152448
rect 408644 152436 408650 152448
rect 417418 152436 417424 152448
rect 408644 152408 417424 152436
rect 408644 152396 408650 152408
rect 417418 152396 417424 152408
rect 417476 152396 417482 152448
rect 418430 152396 418436 152448
rect 418488 152436 418494 152448
rect 438026 152436 438032 152448
rect 418488 152408 438032 152436
rect 418488 152396 418494 152408
rect 438026 152396 438032 152408
rect 438084 152396 438090 152448
rect 438578 152396 438584 152448
rect 438636 152436 438642 152448
rect 453482 152436 453488 152448
rect 438636 152408 453488 152436
rect 438636 152396 438642 152408
rect 453482 152396 453488 152408
rect 453540 152396 453546 152448
rect 514478 152396 514484 152448
rect 514536 152436 514542 152448
rect 517422 152436 517428 152448
rect 514536 152408 517428 152436
rect 514536 152396 514542 152408
rect 517422 152396 517428 152408
rect 517480 152396 517486 152448
rect 91094 152328 91100 152380
rect 91152 152368 91158 152380
rect 179966 152368 179972 152380
rect 91152 152340 179972 152368
rect 91152 152328 91158 152340
rect 179966 152328 179972 152340
rect 180024 152328 180030 152380
rect 181254 152328 181260 152380
rect 181312 152368 181318 152380
rect 256970 152368 256976 152380
rect 181312 152340 256976 152368
rect 181312 152328 181318 152340
rect 256970 152328 256976 152340
rect 257028 152328 257034 152380
rect 260926 152328 260932 152380
rect 260984 152368 260990 152380
rect 316034 152368 316040 152380
rect 260984 152340 316040 152368
rect 260984 152328 260990 152340
rect 316034 152328 316040 152340
rect 316092 152328 316098 152380
rect 320266 152328 320272 152380
rect 320324 152368 320330 152380
rect 323118 152368 323124 152380
rect 320324 152340 323124 152368
rect 320324 152328 320330 152340
rect 323118 152328 323124 152340
rect 323176 152328 323182 152380
rect 323210 152328 323216 152380
rect 323268 152368 323274 152380
rect 330478 152368 330484 152380
rect 323268 152340 330484 152368
rect 323268 152328 323274 152340
rect 330478 152328 330484 152340
rect 330536 152328 330542 152380
rect 330570 152328 330576 152380
rect 330628 152368 330634 152380
rect 367370 152368 367376 152380
rect 330628 152340 367376 152368
rect 330628 152328 330634 152340
rect 367370 152328 367376 152340
rect 367428 152328 367434 152380
rect 381354 152328 381360 152380
rect 381412 152368 381418 152380
rect 409874 152368 409880 152380
rect 381412 152340 409880 152368
rect 381412 152328 381418 152340
rect 409874 152328 409880 152340
rect 409932 152328 409938 152380
rect 413830 152328 413836 152380
rect 413888 152368 413894 152380
rect 416222 152368 416228 152380
rect 413888 152340 416228 152368
rect 413888 152328 413894 152340
rect 416222 152328 416228 152340
rect 416280 152328 416286 152380
rect 416590 152328 416596 152380
rect 416648 152368 416654 152380
rect 416648 152340 417556 152368
rect 416648 152328 416654 152340
rect 33594 152260 33600 152312
rect 33652 152300 33658 152312
rect 109678 152300 109684 152312
rect 33652 152272 109684 152300
rect 33652 152260 33658 152272
rect 109678 152260 109684 152272
rect 109736 152260 109742 152312
rect 109770 152260 109776 152312
rect 109828 152300 109834 152312
rect 127894 152300 127900 152312
rect 109828 152272 127900 152300
rect 109828 152260 109834 152272
rect 127894 152260 127900 152272
rect 127952 152260 127958 152312
rect 127986 152260 127992 152312
rect 128044 152300 128050 152312
rect 215846 152300 215852 152312
rect 128044 152272 215852 152300
rect 128044 152260 128050 152272
rect 215846 152260 215852 152272
rect 215904 152260 215910 152312
rect 223850 152260 223856 152312
rect 223908 152300 223914 152312
rect 287790 152300 287796 152312
rect 223908 152272 287796 152300
rect 223908 152260 223914 152272
rect 287790 152260 287796 152272
rect 287848 152260 287854 152312
rect 288342 152260 288348 152312
rect 288400 152300 288406 152312
rect 289906 152300 289912 152312
rect 288400 152272 289912 152300
rect 288400 152260 288406 152272
rect 289906 152260 289912 152272
rect 289964 152260 289970 152312
rect 292206 152260 292212 152312
rect 292264 152300 292270 152312
rect 341702 152300 341708 152312
rect 292264 152272 341708 152300
rect 292264 152260 292270 152272
rect 341702 152260 341708 152272
rect 341760 152260 341766 152312
rect 342438 152260 342444 152312
rect 342496 152300 342502 152312
rect 344278 152300 344284 152312
rect 342496 152272 344284 152300
rect 342496 152260 342502 152272
rect 344278 152260 344284 152272
rect 344336 152260 344342 152312
rect 345198 152260 345204 152312
rect 345256 152300 345262 152312
rect 382274 152300 382280 152312
rect 345256 152272 382280 152300
rect 345256 152260 345262 152272
rect 382274 152260 382280 152272
rect 382332 152260 382338 152312
rect 382366 152260 382372 152312
rect 382424 152300 382430 152312
rect 386690 152300 386696 152312
rect 382424 152272 386696 152300
rect 382424 152260 382430 152272
rect 386690 152260 386696 152272
rect 386748 152260 386754 152312
rect 389174 152260 389180 152312
rect 389232 152300 389238 152312
rect 412634 152300 412640 152312
rect 389232 152272 412640 152300
rect 389232 152260 389238 152272
rect 412634 152260 412640 152272
rect 412692 152260 412698 152312
rect 9490 152192 9496 152244
rect 9548 152232 9554 152244
rect 82814 152232 82820 152244
rect 9548 152204 82820 152232
rect 9548 152192 9554 152204
rect 82814 152192 82820 152204
rect 82872 152192 82878 152244
rect 82906 152192 82912 152244
rect 82964 152232 82970 152244
rect 169754 152232 169760 152244
rect 82964 152204 169760 152232
rect 82964 152192 82970 152204
rect 169754 152192 169760 152204
rect 169812 152192 169818 152244
rect 169864 152204 175964 152232
rect 78858 152124 78864 152176
rect 78916 152164 78922 152176
rect 164510 152164 164516 152176
rect 78916 152136 164516 152164
rect 78916 152124 78922 152136
rect 164510 152124 164516 152136
rect 164568 152124 164574 152176
rect 166994 152124 167000 152176
rect 167052 152164 167058 152176
rect 169864 152164 169892 152204
rect 167052 152136 169892 152164
rect 167052 152124 167058 152136
rect 169938 152124 169944 152176
rect 169996 152164 170002 152176
rect 175936 152164 175964 152204
rect 176102 152192 176108 152244
rect 176160 152232 176166 152244
rect 190178 152232 190184 152244
rect 176160 152204 190184 152232
rect 176160 152192 176166 152204
rect 190178 152192 190184 152204
rect 190236 152192 190242 152244
rect 194502 152192 194508 152244
rect 194560 152232 194566 152244
rect 213270 152232 213276 152244
rect 194560 152204 213276 152232
rect 194560 152192 194566 152204
rect 213270 152192 213276 152204
rect 213328 152192 213334 152244
rect 221734 152192 221740 152244
rect 221792 152232 221798 152244
rect 282914 152232 282920 152244
rect 221792 152204 282920 152232
rect 221792 152192 221798 152204
rect 282914 152192 282920 152204
rect 282972 152192 282978 152244
rect 285766 152192 285772 152244
rect 285824 152232 285830 152244
rect 335906 152232 335912 152244
rect 285824 152204 335912 152232
rect 285824 152192 285830 152204
rect 335906 152192 335912 152204
rect 335964 152192 335970 152244
rect 341058 152232 341064 152244
rect 338224 152204 341064 152232
rect 182450 152164 182456 152176
rect 169996 152136 175872 152164
rect 175936 152136 182456 152164
rect 169996 152124 170002 152136
rect 68922 152056 68928 152108
rect 68980 152096 68986 152108
rect 149146 152096 149152 152108
rect 68980 152068 149152 152096
rect 68980 152056 68986 152068
rect 149146 152056 149152 152068
rect 149204 152056 149210 152108
rect 156874 152056 156880 152108
rect 156932 152096 156938 152108
rect 172514 152096 172520 152108
rect 156932 152068 172520 152096
rect 156932 152056 156938 152068
rect 172514 152056 172520 152068
rect 172572 152056 172578 152108
rect 175844 152096 175872 152136
rect 182450 152124 182456 152136
rect 182508 152124 182514 152176
rect 183462 152124 183468 152176
rect 183520 152164 183526 152176
rect 183520 152136 186314 152164
rect 183520 152124 183526 152136
rect 185026 152096 185032 152108
rect 175844 152068 185032 152096
rect 185026 152056 185032 152068
rect 185084 152056 185090 152108
rect 186286 152096 186314 152136
rect 191650 152124 191656 152176
rect 191708 152164 191714 152176
rect 208394 152164 208400 152176
rect 191708 152136 208400 152164
rect 191708 152124 191714 152136
rect 208394 152124 208400 152136
rect 208452 152124 208458 152176
rect 213638 152124 213644 152176
rect 213696 152164 213702 152176
rect 274266 152164 274272 152176
rect 213696 152136 274272 152164
rect 213696 152124 213702 152136
rect 274266 152124 274272 152136
rect 274324 152124 274330 152176
rect 277946 152124 277952 152176
rect 278004 152164 278010 152176
rect 279602 152164 279608 152176
rect 278004 152136 279608 152164
rect 278004 152124 278010 152136
rect 279602 152124 279608 152136
rect 279660 152124 279666 152176
rect 291378 152124 291384 152176
rect 291436 152164 291442 152176
rect 338224 152164 338252 152204
rect 341058 152192 341064 152204
rect 341116 152192 341122 152244
rect 341150 152192 341156 152244
rect 341208 152232 341214 152244
rect 375374 152232 375380 152244
rect 341208 152204 375380 152232
rect 341208 152192 341214 152204
rect 375374 152192 375380 152204
rect 375432 152192 375438 152244
rect 385494 152192 385500 152244
rect 385552 152232 385558 152244
rect 387334 152232 387340 152244
rect 385552 152204 387340 152232
rect 385552 152192 385558 152204
rect 387334 152192 387340 152204
rect 387392 152192 387398 152244
rect 388346 152192 388352 152244
rect 388404 152232 388410 152244
rect 388404 152204 393314 152232
rect 388404 152192 388410 152204
rect 291436 152136 338252 152164
rect 291436 152124 291442 152136
rect 340138 152124 340144 152176
rect 340196 152164 340202 152176
rect 346394 152164 346400 152176
rect 340196 152136 346400 152164
rect 340196 152124 340202 152136
rect 346394 152124 346400 152136
rect 346452 152124 346458 152176
rect 349798 152124 349804 152176
rect 349856 152164 349862 152176
rect 380250 152164 380256 152176
rect 349856 152136 380256 152164
rect 349856 152124 349862 152136
rect 380250 152124 380256 152136
rect 380308 152124 380314 152176
rect 383746 152124 383752 152176
rect 383804 152164 383810 152176
rect 391934 152164 391940 152176
rect 383804 152136 391940 152164
rect 383804 152124 383810 152136
rect 391934 152124 391940 152136
rect 391992 152124 391998 152176
rect 393286 152164 393314 152204
rect 394602 152192 394608 152244
rect 394660 152232 394666 152244
rect 417326 152232 417332 152244
rect 394660 152204 417332 152232
rect 394660 152192 394666 152204
rect 417326 152192 417332 152204
rect 417384 152192 417390 152244
rect 417528 152232 417556 152340
rect 421742 152328 421748 152380
rect 421800 152368 421806 152380
rect 436278 152368 436284 152380
rect 421800 152340 436284 152368
rect 421800 152328 421806 152340
rect 436278 152328 436284 152340
rect 436336 152328 436342 152380
rect 441246 152368 441252 152380
rect 436572 152340 441252 152368
rect 417602 152260 417608 152312
rect 417660 152300 417666 152312
rect 421466 152300 421472 152312
rect 417660 152272 421472 152300
rect 417660 152260 417666 152272
rect 421466 152260 421472 152272
rect 421524 152260 421530 152312
rect 425146 152260 425152 152312
rect 425204 152300 425210 152312
rect 425204 152272 426664 152300
rect 425204 152260 425210 152272
rect 426526 152232 426532 152244
rect 417528 152204 426532 152232
rect 426526 152192 426532 152204
rect 426584 152192 426590 152244
rect 426636 152232 426664 152272
rect 426710 152260 426716 152312
rect 426768 152300 426774 152312
rect 436572 152300 436600 152340
rect 441246 152328 441252 152340
rect 441304 152328 441310 152380
rect 441706 152328 441712 152380
rect 441764 152368 441770 152380
rect 455414 152368 455420 152380
rect 441764 152340 455420 152368
rect 441764 152328 441770 152340
rect 455414 152328 455420 152340
rect 455472 152328 455478 152380
rect 426768 152272 436600 152300
rect 426768 152260 426774 152272
rect 441522 152260 441528 152312
rect 441580 152300 441586 152312
rect 454770 152300 454776 152312
rect 441580 152272 454776 152300
rect 441580 152260 441586 152272
rect 454770 152260 454776 152272
rect 454828 152260 454834 152312
rect 443178 152232 443184 152244
rect 426636 152204 443184 152232
rect 443178 152192 443184 152204
rect 443236 152192 443242 152244
rect 443638 152192 443644 152244
rect 443696 152232 443702 152244
rect 457346 152232 457352 152244
rect 443696 152204 457352 152232
rect 443696 152192 443702 152204
rect 457346 152192 457352 152204
rect 457404 152192 457410 152244
rect 407206 152164 407212 152176
rect 393286 152136 407212 152164
rect 407206 152124 407212 152136
rect 407264 152124 407270 152176
rect 409322 152124 409328 152176
rect 409380 152164 409386 152176
rect 428366 152164 428372 152176
rect 409380 152136 428372 152164
rect 409380 152124 409386 152136
rect 428366 152124 428372 152136
rect 428424 152124 428430 152176
rect 429286 152124 429292 152176
rect 429344 152164 429350 152176
rect 446398 152164 446404 152176
rect 429344 152136 446404 152164
rect 429344 152124 429350 152136
rect 446398 152124 446404 152136
rect 446456 152124 446462 152176
rect 200482 152096 200488 152108
rect 186286 152068 200488 152096
rect 200482 152056 200488 152068
rect 200540 152056 200546 152108
rect 242802 152056 242808 152108
rect 242860 152096 242866 152108
rect 300854 152096 300860 152108
rect 242860 152068 300860 152096
rect 242860 152056 242866 152068
rect 300854 152056 300860 152068
rect 300912 152056 300918 152108
rect 303982 152056 303988 152108
rect 304040 152096 304046 152108
rect 350718 152096 350724 152108
rect 304040 152068 350724 152096
rect 304040 152056 304046 152068
rect 350718 152056 350724 152068
rect 350776 152056 350782 152108
rect 355318 152056 355324 152108
rect 355376 152096 355382 152108
rect 389910 152096 389916 152108
rect 355376 152068 389916 152096
rect 355376 152056 355382 152068
rect 389910 152056 389916 152068
rect 389968 152056 389974 152108
rect 405642 152056 405648 152108
rect 405700 152096 405706 152108
rect 405700 152068 416820 152096
rect 405700 152056 405706 152068
rect 75086 151988 75092 152040
rect 75144 152028 75150 152040
rect 154206 152028 154212 152040
rect 75144 152000 154212 152028
rect 75144 151988 75150 152000
rect 154206 151988 154212 152000
rect 154264 151988 154270 152040
rect 162486 151988 162492 152040
rect 162544 152028 162550 152040
rect 177390 152028 177396 152040
rect 162544 152000 177396 152028
rect 162544 151988 162550 152000
rect 177390 151988 177396 152000
rect 177448 151988 177454 152040
rect 184658 151988 184664 152040
rect 184716 152028 184722 152040
rect 195330 152028 195336 152040
rect 184716 152000 195336 152028
rect 184716 151988 184722 152000
rect 195330 151988 195336 152000
rect 195388 151988 195394 152040
rect 243354 151988 243360 152040
rect 243412 152028 243418 152040
rect 302602 152028 302608 152040
rect 243412 152000 302608 152028
rect 243412 151988 243418 152000
rect 302602 151988 302608 152000
rect 302660 151988 302666 152040
rect 325694 152028 325700 152040
rect 316006 152000 325700 152028
rect 19794 151920 19800 151972
rect 19852 151960 19858 151972
rect 97902 151960 97908 151972
rect 19852 151932 97908 151960
rect 19852 151920 19858 151932
rect 97902 151920 97908 151932
rect 97960 151920 97966 151972
rect 103790 151920 103796 151972
rect 103848 151960 103854 151972
rect 109862 151960 109868 151972
rect 103848 151932 109868 151960
rect 103848 151920 103854 151932
rect 109862 151920 109868 151932
rect 109920 151920 109926 151972
rect 109954 151920 109960 151972
rect 110012 151960 110018 151972
rect 138290 151960 138296 151972
rect 110012 151932 138296 151960
rect 110012 151920 110018 151932
rect 138290 151920 138296 151932
rect 138348 151920 138354 151972
rect 139302 151920 139308 151972
rect 139360 151960 139366 151972
rect 203058 151960 203064 151972
rect 139360 151932 171134 151960
rect 139360 151920 139366 151932
rect 74810 151852 74816 151904
rect 74868 151892 74874 151904
rect 81342 151892 81348 151904
rect 74868 151864 81348 151892
rect 74868 151852 74874 151864
rect 81342 151852 81348 151864
rect 81400 151852 81406 151904
rect 109034 151852 109040 151904
rect 109092 151892 109098 151904
rect 130470 151892 130476 151904
rect 109092 151864 130476 151892
rect 109092 151852 109098 151864
rect 130470 151852 130476 151864
rect 130528 151852 130534 151904
rect 130654 151852 130660 151904
rect 130712 151892 130718 151904
rect 146570 151892 146576 151904
rect 130712 151864 146576 151892
rect 130712 151852 130718 151864
rect 146570 151852 146576 151864
rect 146628 151852 146634 151904
rect 146662 151852 146668 151904
rect 146720 151892 146726 151904
rect 167086 151892 167092 151904
rect 146720 151864 167092 151892
rect 146720 151852 146726 151864
rect 167086 151852 167092 151864
rect 167144 151852 167150 151904
rect 171106 151892 171134 151932
rect 176626 151932 203064 151960
rect 176626 151892 176654 151932
rect 203058 151920 203064 151932
rect 203116 151920 203122 151972
rect 213086 151920 213092 151972
rect 213144 151960 213150 151972
rect 272426 151960 272432 151972
rect 213144 151932 272432 151960
rect 213144 151920 213150 151932
rect 272426 151920 272432 151932
rect 272484 151920 272490 151972
rect 272518 151920 272524 151972
rect 272576 151960 272582 151972
rect 316006 151960 316034 152000
rect 325694 151988 325700 152000
rect 325752 151988 325758 152040
rect 330478 151988 330484 152040
rect 330536 152028 330542 152040
rect 362310 152028 362316 152040
rect 330536 152000 362316 152028
rect 330536 151988 330542 152000
rect 362310 151988 362316 152000
rect 362368 151988 362374 152040
rect 387886 151988 387892 152040
rect 387944 152028 387950 152040
rect 404630 152028 404636 152040
rect 387944 152000 404636 152028
rect 387944 151988 387950 152000
rect 404630 151988 404636 152000
rect 404688 151988 404694 152040
rect 413002 152028 413008 152040
rect 407776 152000 413008 152028
rect 272576 151932 316034 151960
rect 272576 151920 272582 151932
rect 325878 151920 325884 151972
rect 325936 151960 325942 151972
rect 330570 151960 330576 151972
rect 325936 151932 330576 151960
rect 325936 151920 325942 151932
rect 330570 151920 330576 151932
rect 330628 151920 330634 151972
rect 331766 151920 331772 151972
rect 331824 151960 331830 151972
rect 371878 151960 371884 151972
rect 331824 151932 371884 151960
rect 331824 151920 331830 151932
rect 371878 151920 371884 151932
rect 371936 151920 371942 151972
rect 378778 151920 378784 151972
rect 378836 151960 378842 151972
rect 384114 151960 384120 151972
rect 378836 151932 384120 151960
rect 378836 151920 378842 151932
rect 384114 151920 384120 151932
rect 384172 151920 384178 151972
rect 385862 151920 385868 151972
rect 385920 151960 385926 151972
rect 399478 151960 399484 151972
rect 385920 151932 399484 151960
rect 385920 151920 385926 151932
rect 399478 151920 399484 151932
rect 399536 151920 399542 151972
rect 399570 151920 399576 151972
rect 399628 151960 399634 151972
rect 407776 151960 407804 152000
rect 413002 151988 413008 152000
rect 413060 151988 413066 152040
rect 416792 152028 416820 152068
rect 417418 152056 417424 152108
rect 417476 152096 417482 152108
rect 417476 152068 422294 152096
rect 417476 152056 417482 152068
rect 420914 152028 420920 152040
rect 416792 152000 420920 152028
rect 420914 151988 420920 152000
rect 420972 151988 420978 152040
rect 422266 152028 422294 152068
rect 422570 152056 422576 152108
rect 422628 152096 422634 152108
rect 426710 152096 426716 152108
rect 422628 152068 426716 152096
rect 422628 152056 422634 152068
rect 426710 152056 426716 152068
rect 426768 152056 426774 152108
rect 426802 152056 426808 152108
rect 426860 152096 426866 152108
rect 444466 152096 444472 152108
rect 426860 152068 444472 152096
rect 426860 152056 426866 152068
rect 444466 152056 444472 152068
rect 444524 152056 444530 152108
rect 515766 152056 515772 152108
rect 515824 152096 515830 152108
rect 518894 152096 518900 152108
rect 515824 152068 518900 152096
rect 515824 152056 515830 152068
rect 518894 152056 518900 152068
rect 518952 152056 518958 152108
rect 423306 152028 423312 152040
rect 422266 152000 423312 152028
rect 423306 151988 423312 152000
rect 423364 151988 423370 152040
rect 423582 151988 423588 152040
rect 423640 152028 423646 152040
rect 439314 152028 439320 152040
rect 423640 152000 439320 152028
rect 423640 151988 423646 152000
rect 439314 151988 439320 152000
rect 439372 151988 439378 152040
rect 439406 151988 439412 152040
rect 439464 152028 439470 152040
rect 454218 152028 454224 152040
rect 439464 152000 454224 152028
rect 439464 151988 439470 152000
rect 454218 151988 454224 152000
rect 454276 151988 454282 152040
rect 459554 151988 459560 152040
rect 459612 152028 459618 152040
rect 461762 152028 461768 152040
rect 459612 152000 461768 152028
rect 459612 151988 459618 152000
rect 461762 151988 461768 152000
rect 461820 151988 461826 152040
rect 486510 151988 486516 152040
rect 486568 152028 486574 152040
rect 490006 152028 490012 152040
rect 486568 152000 490012 152028
rect 486568 151988 486574 152000
rect 490006 151988 490012 152000
rect 490064 151988 490070 152040
rect 515950 151988 515956 152040
rect 516008 152028 516014 152040
rect 519446 152028 519452 152040
rect 516008 152000 519452 152028
rect 516008 151988 516014 152000
rect 519446 151988 519452 152000
rect 519504 151988 519510 152040
rect 399628 151932 407804 151960
rect 399628 151920 399634 151932
rect 413738 151920 413744 151972
rect 413796 151960 413802 151972
rect 413796 151932 418292 151960
rect 413796 151920 413802 151932
rect 171106 151864 176654 151892
rect 283006 151852 283012 151904
rect 283064 151892 283070 151904
rect 287146 151892 287152 151904
rect 283064 151864 287152 151892
rect 283064 151852 283070 151864
rect 287146 151852 287152 151864
rect 287204 151852 287210 151904
rect 299934 151852 299940 151904
rect 299992 151892 299998 151904
rect 340138 151892 340144 151904
rect 299992 151864 340144 151892
rect 299992 151852 299998 151864
rect 340138 151852 340144 151864
rect 340196 151852 340202 151904
rect 349430 151852 349436 151904
rect 349488 151892 349494 151904
rect 349488 151864 373994 151892
rect 349488 151852 349494 151864
rect 71406 151784 71412 151836
rect 71464 151824 71470 151836
rect 92474 151824 92480 151836
rect 71464 151796 92480 151824
rect 71464 151784 71470 151796
rect 92474 151784 92480 151796
rect 92532 151784 92538 151836
rect 105814 151784 105820 151836
rect 105872 151824 105878 151836
rect 110322 151824 110328 151836
rect 105872 151796 110328 151824
rect 105872 151784 105878 151796
rect 110322 151784 110328 151796
rect 110380 151784 110386 151836
rect 113910 151784 113916 151836
rect 113968 151824 113974 151836
rect 120994 151824 121000 151836
rect 113968 151796 121000 151824
rect 113968 151784 113974 151796
rect 120994 151784 121000 151796
rect 121052 151784 121058 151836
rect 138014 151784 138020 151836
rect 138072 151824 138078 151836
rect 141418 151824 141424 151836
rect 138072 151796 141424 151824
rect 138072 151784 138078 151796
rect 141418 151784 141424 151796
rect 141476 151784 141482 151836
rect 142246 151784 142252 151836
rect 142304 151824 142310 151836
rect 151814 151824 151820 151836
rect 142304 151796 151820 151824
rect 142304 151784 142310 151796
rect 151814 151784 151820 151796
rect 151872 151784 151878 151836
rect 154298 151784 154304 151836
rect 154356 151824 154362 151836
rect 236454 151824 236460 151836
rect 154356 151796 236460 151824
rect 154356 151784 154362 151796
rect 236454 151784 236460 151796
rect 236512 151784 236518 151836
rect 272610 151784 272616 151836
rect 272668 151824 272674 151836
rect 326338 151824 326344 151836
rect 272668 151796 326344 151824
rect 272668 151784 272674 151796
rect 326338 151784 326344 151796
rect 326396 151784 326402 151836
rect 335998 151784 336004 151836
rect 336056 151824 336062 151836
rect 341150 151824 341156 151836
rect 336056 151796 341156 151824
rect 336056 151784 336062 151796
rect 341150 151784 341156 151796
rect 341208 151784 341214 151836
rect 343818 151784 343824 151836
rect 343876 151824 343882 151836
rect 349798 151824 349804 151836
rect 343876 151796 349804 151824
rect 343876 151784 343882 151796
rect 349798 151784 349804 151796
rect 349856 151784 349862 151836
rect 362954 151784 362960 151836
rect 363012 151824 363018 151836
rect 364334 151824 364340 151836
rect 363012 151796 364340 151824
rect 363012 151784 363018 151796
rect 364334 151784 364340 151796
rect 364392 151784 364398 151836
rect 373966 151824 373994 151864
rect 386322 151852 386328 151904
rect 386380 151892 386386 151904
rect 394694 151892 394700 151904
rect 386380 151864 394700 151892
rect 386380 151852 386386 151864
rect 394694 151852 394700 151864
rect 394752 151852 394758 151904
rect 396258 151852 396264 151904
rect 396316 151892 396322 151904
rect 402974 151892 402980 151904
rect 396316 151864 402980 151892
rect 396316 151852 396322 151864
rect 402974 151852 402980 151864
rect 403032 151852 403038 151904
rect 404262 151852 404268 151904
rect 404320 151892 404326 151904
rect 418154 151892 418160 151904
rect 404320 151864 418160 151892
rect 404320 151852 404326 151864
rect 418154 151852 418160 151864
rect 418212 151852 418218 151904
rect 418264 151892 418292 151932
rect 419626 151920 419632 151972
rect 419684 151960 419690 151972
rect 436738 151960 436744 151972
rect 419684 151932 436744 151960
rect 419684 151920 419690 151932
rect 436738 151920 436744 151932
rect 436796 151920 436802 151972
rect 451550 151960 451556 151972
rect 440712 151932 451556 151960
rect 421374 151892 421380 151904
rect 418264 151864 421380 151892
rect 421374 151852 421380 151864
rect 421432 151852 421438 151904
rect 421466 151852 421472 151904
rect 421524 151892 421530 151904
rect 431586 151892 431592 151904
rect 421524 151864 431592 151892
rect 421524 151852 421530 151864
rect 431586 151852 431592 151864
rect 431644 151852 431650 151904
rect 436278 151852 436284 151904
rect 436336 151892 436342 151904
rect 440602 151892 440608 151904
rect 436336 151864 440608 151892
rect 436336 151852 436342 151864
rect 440602 151852 440608 151864
rect 440660 151852 440666 151904
rect 385402 151824 385408 151836
rect 373966 151796 385408 151824
rect 385402 151784 385408 151796
rect 385460 151784 385466 151836
rect 403894 151784 403900 151836
rect 403952 151824 403958 151836
rect 415670 151824 415676 151836
rect 403952 151796 415676 151824
rect 403952 151784 403958 151796
rect 415670 151784 415676 151796
rect 415728 151784 415734 151836
rect 419718 151784 419724 151836
rect 419776 151824 419782 151836
rect 434162 151824 434168 151836
rect 419776 151796 434168 151824
rect 419776 151784 419782 151796
rect 434162 151784 434168 151796
rect 434220 151784 434226 151836
rect 436186 151784 436192 151836
rect 436244 151824 436250 151836
rect 440712 151824 440740 151932
rect 451550 151920 451556 151932
rect 451608 151920 451614 151972
rect 469214 151920 469220 151972
rect 469272 151960 469278 151972
rect 472066 151960 472072 151972
rect 469272 151932 472072 151960
rect 469272 151920 469278 151932
rect 472066 151920 472072 151932
rect 472124 151920 472130 151972
rect 487338 151920 487344 151972
rect 487396 151960 487402 151972
rect 490650 151960 490656 151972
rect 487396 151932 490656 151960
rect 487396 151920 487402 151932
rect 490650 151920 490656 151932
rect 490708 151920 490714 151972
rect 507762 151920 507768 151972
rect 507820 151960 507826 151972
rect 509234 151960 509240 151972
rect 507820 151932 509240 151960
rect 507820 151920 507826 151932
rect 509234 151920 509240 151932
rect 509292 151920 509298 151972
rect 517422 151920 517428 151972
rect 517480 151960 517486 151972
rect 521562 151960 521568 151972
rect 517480 151932 521568 151960
rect 517480 151920 517486 151932
rect 521562 151920 521568 151932
rect 521620 151920 521626 151972
rect 442902 151852 442908 151904
rect 442960 151892 442966 151904
rect 450906 151892 450912 151904
rect 442960 151864 450912 151892
rect 442960 151852 442966 151864
rect 450906 151852 450912 151864
rect 450964 151852 450970 151904
rect 468018 151852 468024 151904
rect 468076 151892 468082 151904
rect 470778 151892 470784 151904
rect 468076 151864 470784 151892
rect 468076 151852 468082 151864
rect 470778 151852 470784 151864
rect 470836 151852 470842 151904
rect 489086 151852 489092 151904
rect 489144 151892 489150 151904
rect 491938 151892 491944 151904
rect 489144 151864 491944 151892
rect 489144 151852 489150 151864
rect 491938 151852 491944 151864
rect 491996 151852 492002 151904
rect 436244 151796 440740 151824
rect 436244 151784 436250 151796
rect 442718 151784 442724 151836
rect 442776 151824 442782 151836
rect 456058 151824 456064 151836
rect 442776 151796 456064 151824
rect 442776 151784 442782 151796
rect 456058 151784 456064 151796
rect 456116 151784 456122 151836
rect 467834 151784 467840 151836
rect 467892 151824 467898 151836
rect 471422 151824 471428 151836
rect 467892 151796 471428 151824
rect 467892 151784 467898 151796
rect 471422 151784 471428 151796
rect 471480 151784 471486 151836
rect 488442 151784 488448 151836
rect 488500 151824 488506 151836
rect 491294 151824 491300 151836
rect 488500 151796 491300 151824
rect 488500 151784 488506 151796
rect 491294 151784 491300 151796
rect 491352 151784 491358 151836
rect 509050 151784 509056 151836
rect 509108 151824 509114 151836
rect 510890 151824 510896 151836
rect 509108 151796 510896 151824
rect 509108 151784 509114 151796
rect 510890 151784 510896 151796
rect 510948 151784 510954 151836
rect 517054 151784 517060 151836
rect 517112 151824 517118 151836
rect 520274 151824 520280 151836
rect 517112 151796 520280 151824
rect 517112 151784 517118 151796
rect 520274 151784 520280 151796
rect 520332 151784 520338 151836
rect 81710 151716 81716 151768
rect 81768 151756 81774 151768
rect 112898 151756 112904 151768
rect 81768 151728 112904 151756
rect 81768 151716 81774 151728
rect 112898 151716 112904 151728
rect 112956 151716 112962 151768
rect 98914 151648 98920 151700
rect 98972 151688 98978 151700
rect 116026 151688 116032 151700
rect 98972 151660 116032 151688
rect 98972 151648 98978 151660
rect 116026 151648 116032 151660
rect 116084 151648 116090 151700
rect 95510 151580 95516 151632
rect 95568 151620 95574 151632
rect 115290 151620 115296 151632
rect 95568 151592 115296 151620
rect 95568 151580 95574 151592
rect 115290 151580 115296 151592
rect 115348 151580 115354 151632
rect 92014 151512 92020 151564
rect 92072 151552 92078 151564
rect 113082 151552 113088 151564
rect 92072 151524 113088 151552
rect 92072 151512 92078 151524
rect 113082 151512 113088 151524
rect 113140 151512 113146 151564
rect 26694 151444 26700 151496
rect 26752 151484 26758 151496
rect 116946 151484 116952 151496
rect 26752 151456 116952 151484
rect 26752 151444 26758 151456
rect 116946 151444 116952 151456
rect 117004 151444 117010 151496
rect 16390 151376 16396 151428
rect 16448 151416 16454 151428
rect 116762 151416 116768 151428
rect 16448 151388 116768 151416
rect 16448 151376 16454 151388
rect 116762 151376 116768 151388
rect 116820 151376 116826 151428
rect 12986 151308 12992 151360
rect 13044 151348 13050 151360
rect 116670 151348 116676 151360
rect 13044 151320 116676 151348
rect 13044 151308 13050 151320
rect 116670 151308 116676 151320
rect 116728 151308 116734 151360
rect 68002 151240 68008 151292
rect 68060 151280 68066 151292
rect 112714 151280 112720 151292
rect 68060 151252 112720 151280
rect 68060 151240 68066 151252
rect 112714 151240 112720 151252
rect 112772 151240 112778 151292
rect 64506 151172 64512 151224
rect 64564 151212 64570 151224
rect 112622 151212 112628 151224
rect 64564 151184 112628 151212
rect 64564 151172 64570 151184
rect 112622 151172 112628 151184
rect 112680 151172 112686 151224
rect 61102 151104 61108 151156
rect 61160 151144 61166 151156
rect 112530 151144 112536 151156
rect 61160 151116 112536 151144
rect 61160 151104 61166 151116
rect 112530 151104 112536 151116
rect 112588 151104 112594 151156
rect 57698 151036 57704 151088
rect 57756 151076 57762 151088
rect 110966 151076 110972 151088
rect 57756 151048 110972 151076
rect 57756 151036 57762 151048
rect 110966 151036 110972 151048
rect 111024 151036 111030 151088
rect 54202 150968 54208 151020
rect 54260 151008 54266 151020
rect 112438 151008 112444 151020
rect 54260 150980 112444 151008
rect 54260 150968 54266 150980
rect 112438 150968 112444 150980
rect 112496 150968 112502 151020
rect 50798 150900 50804 150952
rect 50856 150940 50862 150952
rect 111702 150940 111708 150952
rect 50856 150912 111708 150940
rect 50856 150900 50862 150912
rect 111702 150900 111708 150912
rect 111760 150900 111766 150952
rect 47302 150832 47308 150884
rect 47360 150872 47366 150884
rect 111610 150872 111616 150884
rect 47360 150844 111616 150872
rect 47360 150832 47366 150844
rect 111610 150832 111616 150844
rect 111668 150832 111674 150884
rect 43898 150764 43904 150816
rect 43956 150804 43962 150816
rect 111518 150804 111524 150816
rect 43956 150776 111524 150804
rect 43956 150764 43962 150776
rect 111518 150764 111524 150776
rect 111576 150764 111582 150816
rect 40494 150696 40500 150748
rect 40552 150736 40558 150748
rect 111426 150736 111432 150748
rect 40552 150708 111432 150736
rect 40552 150696 40558 150708
rect 111426 150696 111432 150708
rect 111484 150696 111490 150748
rect 36998 150628 37004 150680
rect 37056 150668 37062 150680
rect 111242 150668 111248 150680
rect 37056 150640 111248 150668
rect 37056 150628 37062 150640
rect 111242 150628 111248 150640
rect 111300 150628 111306 150680
rect 88610 150560 88616 150612
rect 88668 150600 88674 150612
rect 112990 150600 112996 150612
rect 88668 150572 112996 150600
rect 88668 150560 88674 150572
rect 112990 150560 112996 150572
rect 113048 150560 113054 150612
rect 85206 150492 85212 150544
rect 85264 150532 85270 150544
rect 115198 150532 115204 150544
rect 85264 150504 115204 150532
rect 85264 150492 85270 150504
rect 115198 150492 115204 150504
rect 115256 150492 115262 150544
rect 285674 150492 285680 150544
rect 285732 150532 285738 150544
rect 286502 150532 286508 150544
rect 285732 150504 286508 150532
rect 285732 150492 285738 150504
rect 286502 150492 286508 150504
rect 286560 150492 286566 150544
rect 342254 150492 342260 150544
rect 342312 150532 342318 150544
rect 342990 150532 342996 150544
rect 342312 150504 342996 150532
rect 342312 150492 342318 150504
rect 342990 150492 342996 150504
rect 343048 150492 343054 150544
rect 102318 150424 102324 150476
rect 102376 150464 102382 150476
rect 116118 150464 116124 150476
rect 102376 150436 116124 150464
rect 102376 150424 102382 150436
rect 116118 150424 116124 150436
rect 116176 150424 116182 150476
rect 78306 150288 78312 150340
rect 78364 150328 78370 150340
rect 112806 150328 112812 150340
rect 78364 150300 112812 150328
rect 78364 150288 78370 150300
rect 112806 150288 112812 150300
rect 112864 150288 112870 150340
rect 109586 150220 109592 150272
rect 109644 150260 109650 150272
rect 117130 150260 117136 150272
rect 109644 150232 117136 150260
rect 109644 150220 109650 150232
rect 117130 150220 117136 150232
rect 117188 150220 117194 150272
rect 97902 150152 97908 150204
rect 97960 150192 97966 150204
rect 116854 150192 116860 150204
rect 97960 150164 116860 150192
rect 97960 150152 97966 150164
rect 116854 150152 116860 150164
rect 116912 150152 116918 150204
rect 81342 150084 81348 150136
rect 81400 150124 81406 150136
rect 81400 150096 84194 150124
rect 81400 150084 81406 150096
rect 84166 150056 84194 150096
rect 92474 150084 92480 150136
rect 92532 150124 92538 150136
rect 117222 150124 117228 150136
rect 92532 150096 117228 150124
rect 92532 150084 92538 150096
rect 117222 150084 117228 150096
rect 117280 150084 117286 150136
rect 116486 150056 116492 150068
rect 84166 150028 116492 150056
rect 116486 150016 116492 150028
rect 116544 150016 116550 150068
rect 111150 148316 111156 148368
rect 111208 148356 111214 148368
rect 117038 148356 117044 148368
rect 111208 148328 117044 148356
rect 111208 148316 111214 148328
rect 117038 148316 117044 148328
rect 117096 148316 117102 148368
rect 113082 140700 113088 140752
rect 113140 140740 113146 140752
rect 116118 140740 116124 140752
rect 113140 140712 116124 140740
rect 113140 140700 113146 140712
rect 116118 140700 116124 140712
rect 116176 140700 116182 140752
rect 112990 137912 112996 137964
rect 113048 137952 113054 137964
rect 116118 137952 116124 137964
rect 113048 137924 116124 137952
rect 113048 137912 113054 137924
rect 116118 137912 116124 137924
rect 116176 137912 116182 137964
rect 112898 133832 112904 133884
rect 112956 133872 112962 133884
rect 116026 133872 116032 133884
rect 112956 133844 116032 133872
rect 112956 133832 112962 133844
rect 116026 133832 116032 133844
rect 116084 133832 116090 133884
rect 114186 132608 114192 132660
rect 114244 132648 114250 132660
rect 115198 132648 115204 132660
rect 114244 132620 115204 132648
rect 114244 132608 114250 132620
rect 115198 132608 115204 132620
rect 115256 132608 115262 132660
rect 112806 132404 112812 132456
rect 112864 132444 112870 132456
rect 116118 132444 116124 132456
rect 112864 132416 116124 132444
rect 112864 132404 112870 132416
rect 116118 132404 116124 132416
rect 116176 132404 116182 132456
rect 112714 126896 112720 126948
rect 112772 126936 112778 126948
rect 116118 126936 116124 126948
rect 112772 126908 116124 126936
rect 112772 126896 112778 126908
rect 116118 126896 116124 126908
rect 116176 126896 116182 126948
rect 112622 124108 112628 124160
rect 112680 124148 112686 124160
rect 116118 124148 116124 124160
rect 112680 124120 116124 124148
rect 112680 124108 112686 124120
rect 116118 124108 116124 124120
rect 116176 124108 116182 124160
rect 112530 122748 112536 122800
rect 112588 122788 112594 122800
rect 115934 122788 115940 122800
rect 112588 122760 115940 122788
rect 112588 122748 112594 122760
rect 115934 122748 115940 122760
rect 115992 122748 115998 122800
rect 111702 121388 111708 121440
rect 111760 121428 111766 121440
rect 116118 121428 116124 121440
rect 111760 121400 116124 121428
rect 111760 121388 111766 121400
rect 116118 121388 116124 121400
rect 116176 121388 116182 121440
rect 112438 118600 112444 118652
rect 112496 118640 112502 118652
rect 116118 118640 116124 118652
rect 112496 118612 116124 118640
rect 112496 118600 112502 118612
rect 116118 118600 116124 118612
rect 116176 118600 116182 118652
rect 111610 117240 111616 117292
rect 111668 117280 111674 117292
rect 116118 117280 116124 117292
rect 111668 117252 116124 117280
rect 111668 117240 111674 117252
rect 116118 117240 116124 117252
rect 116176 117240 116182 117292
rect 111518 114452 111524 114504
rect 111576 114492 111582 114504
rect 116118 114492 116124 114504
rect 111576 114464 116124 114492
rect 111576 114452 111582 114464
rect 116118 114452 116124 114464
rect 116176 114452 116182 114504
rect 111426 113092 111432 113144
rect 111484 113132 111490 113144
rect 115934 113132 115940 113144
rect 111484 113104 115940 113132
rect 111484 113092 111490 113104
rect 115934 113092 115940 113104
rect 115992 113092 115998 113144
rect 111334 111732 111340 111784
rect 111392 111772 111398 111784
rect 116118 111772 116124 111784
rect 111392 111744 116124 111772
rect 111392 111732 111398 111744
rect 116118 111732 116124 111744
rect 116176 111732 116182 111784
rect 111150 108944 111156 108996
rect 111208 108984 111214 108996
rect 116118 108984 116124 108996
rect 111208 108956 116124 108984
rect 111208 108944 111214 108956
rect 116118 108944 116124 108956
rect 116176 108944 116182 108996
rect 111242 92420 111248 92472
rect 111300 92460 111306 92472
rect 116118 92460 116124 92472
rect 111300 92432 116124 92460
rect 111300 92420 111306 92432
rect 116118 92420 116124 92432
rect 116176 92420 116182 92472
rect 111058 89632 111064 89684
rect 111116 89672 111122 89684
rect 116118 89672 116124 89684
rect 111116 89644 116124 89672
rect 111116 89632 111122 89644
rect 116118 89632 116124 89644
rect 116176 89632 116182 89684
rect 113818 88272 113824 88324
rect 113876 88312 113882 88324
rect 116026 88312 116032 88324
rect 113876 88284 116032 88312
rect 113876 88272 113882 88284
rect 116026 88272 116032 88284
rect 116084 88272 116090 88324
rect 113910 83920 113916 83972
rect 113968 83960 113974 83972
rect 116578 83960 116584 83972
rect 113968 83932 116584 83960
rect 113968 83920 113974 83932
rect 116578 83920 116584 83932
rect 116636 83920 116642 83972
rect 114002 82764 114008 82816
rect 114060 82804 114066 82816
rect 116210 82804 116216 82816
rect 114060 82776 116216 82804
rect 114060 82764 114066 82776
rect 116210 82764 116216 82776
rect 116268 82764 116274 82816
rect 114094 79976 114100 80028
rect 114152 80016 114158 80028
rect 115934 80016 115940 80028
rect 114152 79988 115940 80016
rect 114152 79976 114158 79988
rect 115934 79976 115940 79988
rect 115992 79976 115998 80028
rect 114186 78616 114192 78668
rect 114244 78656 114250 78668
rect 116118 78656 116124 78668
rect 114244 78628 116124 78656
rect 114244 78616 114250 78628
rect 116118 78616 116124 78628
rect 116176 78616 116182 78668
rect 114186 71748 114192 71800
rect 114244 71788 114250 71800
rect 116578 71788 116584 71800
rect 114244 71760 116584 71788
rect 114244 71748 114250 71760
rect 116578 71748 116584 71760
rect 116636 71748 116642 71800
rect 114094 69028 114100 69080
rect 114152 69068 114158 69080
rect 116302 69068 116308 69080
rect 114152 69040 116308 69068
rect 114152 69028 114158 69040
rect 116302 69028 116308 69040
rect 116360 69028 116366 69080
rect 114002 67600 114008 67652
rect 114060 67640 114066 67652
rect 116118 67640 116124 67652
rect 114060 67612 116124 67640
rect 114060 67600 114066 67612
rect 116118 67600 116124 67612
rect 116176 67600 116182 67652
rect 113910 66240 113916 66292
rect 113968 66280 113974 66292
rect 116578 66280 116584 66292
rect 113968 66252 116584 66280
rect 113968 66240 113974 66252
rect 116578 66240 116584 66252
rect 116636 66240 116642 66292
rect 113358 64676 113364 64728
rect 113416 64716 113422 64728
rect 116578 64716 116584 64728
rect 113416 64688 116584 64716
rect 113416 64676 113422 64688
rect 116578 64676 116584 64688
rect 116636 64676 116642 64728
rect 113818 63520 113824 63572
rect 113876 63560 113882 63572
rect 116210 63560 116216 63572
rect 113876 63532 116216 63560
rect 113876 63520 113882 63532
rect 116210 63520 116216 63532
rect 116268 63520 116274 63572
rect 112438 62092 112444 62144
rect 112496 62132 112502 62144
rect 116118 62132 116124 62144
rect 112496 62104 116124 62132
rect 112496 62092 112502 62104
rect 116118 62092 116124 62104
rect 116176 62092 116182 62144
rect 112530 42780 112536 42832
rect 112588 42820 112594 42832
rect 116118 42820 116124 42832
rect 112588 42792 116124 42820
rect 112588 42780 112594 42792
rect 116118 42780 116124 42792
rect 116176 42780 116182 42832
rect 116394 7624 116400 7676
rect 116452 7624 116458 7676
rect 116302 7420 116308 7472
rect 116360 7460 116366 7472
rect 116412 7460 116440 7624
rect 116360 7432 116440 7460
rect 116360 7420 116366 7432
rect 111702 2796 111708 2848
rect 111760 2836 111766 2848
rect 111760 2808 143672 2836
rect 111760 2796 111766 2808
rect 143644 2508 143672 2808
rect 425808 2808 443684 2836
rect 425808 2508 425836 2808
rect 443656 2508 443684 2808
rect 143626 2456 143632 2508
rect 143684 2456 143690 2508
rect 425790 2456 425796 2508
rect 425848 2456 425854 2508
rect 443638 2456 443644 2508
rect 443696 2456 443702 2508
rect 92446 1924 99972 1952
rect 42058 1844 42064 1896
rect 42116 1884 42122 1896
rect 44726 1884 44732 1896
rect 42116 1856 44732 1884
rect 42116 1844 42122 1856
rect 44726 1844 44732 1856
rect 44784 1844 44790 1896
rect 58986 1844 58992 1896
rect 59044 1884 59050 1896
rect 66990 1884 66996 1896
rect 59044 1856 66996 1884
rect 59044 1844 59050 1856
rect 66990 1844 66996 1856
rect 67048 1844 67054 1896
rect 90358 1844 90364 1896
rect 90416 1884 90422 1896
rect 92446 1884 92474 1924
rect 99944 1896 99972 1924
rect 102106 1924 109816 1952
rect 90416 1856 92474 1884
rect 90416 1844 90422 1856
rect 92566 1844 92572 1896
rect 92624 1884 92630 1896
rect 95326 1884 95332 1896
rect 92624 1856 95332 1884
rect 92624 1844 92630 1856
rect 95326 1844 95332 1856
rect 95384 1844 95390 1896
rect 99926 1844 99932 1896
rect 99984 1844 99990 1896
rect 100018 1844 100024 1896
rect 100076 1884 100082 1896
rect 102106 1884 102134 1924
rect 109788 1896 109816 1924
rect 100076 1856 102134 1884
rect 100076 1844 100082 1856
rect 102686 1844 102692 1896
rect 102744 1884 102750 1896
rect 102744 1856 105860 1884
rect 102744 1844 102750 1856
rect 59170 1776 59176 1828
rect 59228 1816 59234 1828
rect 63034 1816 63040 1828
rect 59228 1788 63040 1816
rect 59228 1776 59234 1788
rect 63034 1776 63040 1788
rect 63092 1776 63098 1828
rect 89346 1776 89352 1828
rect 89404 1816 89410 1828
rect 105832 1816 105860 1856
rect 105906 1844 105912 1896
rect 105964 1884 105970 1896
rect 109126 1884 109132 1896
rect 105964 1856 109132 1884
rect 105964 1844 105970 1856
rect 109126 1844 109132 1856
rect 109184 1844 109190 1896
rect 109678 1884 109684 1896
rect 109236 1856 109684 1884
rect 109236 1816 109264 1856
rect 109678 1844 109684 1856
rect 109736 1844 109742 1896
rect 109770 1844 109776 1896
rect 109828 1844 109834 1896
rect 109862 1844 109868 1896
rect 109920 1884 109926 1896
rect 109920 1856 118694 1884
rect 109920 1844 109926 1856
rect 89404 1788 104204 1816
rect 105832 1788 109264 1816
rect 89404 1776 89410 1788
rect 59354 1708 59360 1760
rect 59412 1748 59418 1760
rect 76558 1748 76564 1760
rect 59412 1720 76564 1748
rect 59412 1708 59418 1720
rect 76558 1708 76564 1720
rect 76616 1708 76622 1760
rect 86034 1708 86040 1760
rect 86092 1748 86098 1760
rect 104176 1748 104204 1788
rect 109310 1776 109316 1828
rect 109368 1816 109374 1828
rect 112438 1816 112444 1828
rect 109368 1788 112444 1816
rect 109368 1776 109374 1788
rect 112438 1776 112444 1788
rect 112496 1776 112502 1828
rect 109954 1748 109960 1760
rect 86092 1720 104112 1748
rect 104176 1720 109960 1748
rect 86092 1708 86098 1720
rect 82630 1640 82636 1692
rect 82688 1680 82694 1692
rect 103974 1680 103980 1692
rect 82688 1652 103980 1680
rect 82688 1640 82694 1652
rect 103974 1640 103980 1652
rect 104032 1640 104038 1692
rect 104084 1680 104112 1720
rect 109954 1708 109960 1720
rect 110012 1708 110018 1760
rect 110046 1708 110052 1760
rect 110104 1748 110110 1760
rect 116578 1748 116584 1760
rect 110104 1720 116584 1748
rect 110104 1708 110110 1720
rect 116578 1708 116584 1720
rect 116636 1708 116642 1760
rect 104084 1652 109172 1680
rect 69290 1572 69296 1624
rect 69348 1612 69354 1624
rect 101766 1612 101772 1624
rect 69348 1584 101772 1612
rect 69348 1572 69354 1584
rect 101766 1572 101772 1584
rect 101824 1572 101830 1624
rect 105906 1612 105912 1624
rect 103900 1584 105912 1612
rect 79318 1504 79324 1556
rect 79376 1544 79382 1556
rect 103900 1544 103928 1584
rect 105906 1572 105912 1584
rect 105964 1572 105970 1624
rect 105998 1572 106004 1624
rect 106056 1612 106062 1624
rect 109034 1612 109040 1624
rect 106056 1584 109040 1612
rect 106056 1572 106062 1584
rect 109034 1572 109040 1584
rect 109092 1572 109098 1624
rect 109144 1612 109172 1652
rect 109218 1640 109224 1692
rect 109276 1680 109282 1692
rect 110598 1680 110604 1692
rect 109276 1652 110604 1680
rect 109276 1640 109282 1652
rect 110598 1640 110604 1652
rect 110656 1640 110662 1692
rect 110138 1612 110144 1624
rect 109144 1584 110144 1612
rect 110138 1572 110144 1584
rect 110196 1572 110202 1624
rect 79376 1516 103928 1544
rect 79376 1504 79382 1516
rect 103974 1504 103980 1556
rect 104032 1544 104038 1556
rect 110230 1544 110236 1556
rect 104032 1516 110236 1544
rect 104032 1504 104038 1516
rect 110230 1504 110236 1516
rect 110288 1504 110294 1556
rect 46014 1436 46020 1488
rect 46072 1476 46078 1488
rect 64598 1476 64604 1488
rect 46072 1448 64604 1476
rect 46072 1436 46078 1448
rect 64598 1436 64604 1448
rect 64656 1436 64662 1488
rect 72694 1436 72700 1488
rect 72752 1476 72758 1488
rect 109586 1476 109592 1488
rect 72752 1448 109592 1476
rect 72752 1436 72758 1448
rect 109586 1436 109592 1448
rect 109644 1436 109650 1488
rect 118666 1476 118694 1856
rect 193582 1476 193588 1488
rect 118666 1448 193588 1476
rect 193582 1436 193588 1448
rect 193640 1436 193646 1488
rect 32674 1368 32680 1420
rect 32732 1408 32738 1420
rect 109126 1408 109132 1420
rect 32732 1380 109132 1408
rect 32732 1368 32738 1380
rect 109126 1368 109132 1380
rect 109184 1368 109190 1420
rect 109218 1368 109224 1420
rect 109276 1408 109282 1420
rect 110046 1408 110052 1420
rect 109276 1380 110052 1408
rect 109276 1368 109282 1380
rect 110046 1368 110052 1380
rect 110104 1368 110110 1420
rect 116394 1408 116400 1420
rect 110156 1380 116400 1408
rect 2682 1300 2688 1352
rect 2740 1340 2746 1352
rect 2740 1312 109356 1340
rect 2740 1300 2746 1312
rect 35986 1232 35992 1284
rect 36044 1272 36050 1284
rect 109328 1272 109356 1312
rect 109402 1300 109408 1352
rect 109460 1340 109466 1352
rect 110156 1340 110184 1380
rect 116394 1368 116400 1380
rect 116452 1368 116458 1420
rect 294782 1368 294788 1420
rect 294840 1408 294846 1420
rect 343634 1408 343640 1420
rect 294840 1380 343640 1408
rect 294840 1368 294846 1380
rect 343634 1368 343640 1380
rect 343692 1368 343698 1420
rect 491294 1368 491300 1420
rect 491352 1408 491358 1420
rect 493594 1408 493600 1420
rect 491352 1380 493600 1408
rect 491352 1368 491358 1380
rect 493594 1368 493600 1380
rect 493652 1368 493658 1420
rect 109460 1312 110184 1340
rect 109460 1300 109466 1312
rect 116302 1272 116308 1284
rect 36044 1244 109264 1272
rect 109328 1244 116308 1272
rect 36044 1232 36050 1244
rect 39298 1164 39304 1216
rect 39356 1204 39362 1216
rect 109034 1204 109040 1216
rect 39356 1176 109040 1204
rect 39356 1164 39362 1176
rect 109034 1164 109040 1176
rect 109092 1164 109098 1216
rect 109236 1204 109264 1244
rect 116302 1232 116308 1244
rect 116360 1232 116366 1284
rect 116486 1204 116492 1216
rect 109236 1176 116492 1204
rect 116486 1164 116492 1176
rect 116544 1164 116550 1216
rect 49326 1096 49332 1148
rect 49384 1136 49390 1148
rect 117038 1136 117044 1148
rect 49384 1108 117044 1136
rect 49384 1096 49390 1108
rect 117038 1096 117044 1108
rect 117096 1096 117102 1148
rect 52638 1028 52644 1080
rect 52696 1068 52702 1080
rect 52696 1040 109172 1068
rect 52696 1028 52702 1040
rect 65978 960 65984 1012
rect 66036 1000 66042 1012
rect 101398 1000 101404 1012
rect 66036 972 101404 1000
rect 66036 960 66042 972
rect 101398 960 101404 972
rect 101456 960 101462 1012
rect 109144 1000 109172 1040
rect 116854 1000 116860 1012
rect 101508 972 106274 1000
rect 109144 972 116860 1000
rect 76006 892 76012 944
rect 76064 932 76070 944
rect 101508 932 101536 972
rect 76064 904 101536 932
rect 106246 932 106274 972
rect 116854 960 116860 972
rect 116912 960 116918 1012
rect 112530 932 112536 944
rect 106246 904 112536 932
rect 76064 892 76070 904
rect 112530 892 112536 904
rect 112588 892 112594 944
rect 89714 824 89720 876
rect 89772 864 89778 876
rect 89772 836 93854 864
rect 89772 824 89778 836
rect 93826 796 93854 836
rect 95970 824 95976 876
rect 96028 864 96034 876
rect 100846 864 100852 876
rect 96028 836 100852 864
rect 96028 824 96034 836
rect 100846 824 100852 836
rect 100904 824 100910 876
rect 101398 824 101404 876
rect 101456 864 101462 876
rect 116670 864 116676 876
rect 101456 836 116676 864
rect 101456 824 101462 836
rect 116670 824 116676 836
rect 116728 824 116734 876
rect 102778 796 102784 808
rect 93826 768 102784 796
rect 102778 756 102784 768
rect 102836 756 102842 808
rect 109034 756 109040 808
rect 109092 796 109098 808
rect 117222 796 117228 808
rect 109092 768 117228 796
rect 109092 756 109098 768
rect 117222 756 117228 768
rect 117280 756 117286 808
<< via1 >>
rect 63408 160012 63460 160064
rect 144920 160080 144972 160132
rect 141884 160012 141936 160064
rect 154488 160012 154540 160064
rect 156788 160012 156840 160064
rect 191748 160012 191800 160064
rect 197176 160012 197228 160064
rect 207112 160012 207164 160064
rect 211436 160012 211488 160064
rect 280344 160012 280396 160064
rect 281264 160012 281316 160064
rect 330668 160080 330720 160132
rect 327448 160012 327500 160064
rect 333980 160012 334032 160064
rect 334256 160012 334308 160064
rect 336096 160080 336148 160132
rect 335084 160012 335136 160064
rect 338488 160012 338540 160064
rect 339500 160012 339552 160064
rect 374460 160012 374512 160064
rect 378876 160012 378928 160064
rect 398104 160012 398156 160064
rect 455420 160012 455472 160064
rect 466644 160012 466696 160064
rect 468024 160012 468076 160064
rect 476028 160012 476080 160064
rect 25596 159944 25648 159996
rect 109960 159944 110012 159996
rect 117228 159944 117280 159996
rect 191656 159944 191708 159996
rect 198004 159944 198056 159996
rect 269764 159944 269816 159996
rect 271236 159944 271288 159996
rect 272524 159944 272576 159996
rect 275376 159944 275428 159996
rect 328828 159944 328880 159996
rect 329196 159944 329248 159996
rect 370044 159944 370096 159996
rect 372160 159944 372212 159996
rect 396264 159944 396316 159996
rect 403256 159944 403308 159996
rect 416596 159944 416648 159996
rect 467196 159944 467248 159996
rect 473360 159944 473412 159996
rect 76932 159876 76984 159928
rect 162492 159876 162544 159928
rect 166908 159876 166960 159928
rect 186412 159876 186464 159928
rect 191288 159876 191340 159928
rect 264888 159876 264940 159928
rect 268660 159876 268712 159928
rect 323676 159876 323728 159928
rect 328368 159876 328420 159928
rect 369216 159876 369268 159928
rect 373632 159876 373684 159928
rect 379428 159876 379480 159928
rect 379704 159876 379756 159928
rect 405832 159876 405884 159928
rect 409972 159876 410024 159928
rect 417608 159876 417660 159928
rect 480628 159876 480680 159928
rect 485872 159876 485924 159928
rect 70124 159808 70176 159860
rect 156880 159808 156932 159860
rect 166264 159808 166316 159860
rect 172428 159808 172480 159860
rect 56692 159740 56744 159792
rect 137284 159740 137336 159792
rect 137376 159740 137428 159792
rect 139584 159740 139636 159792
rect 139860 159740 139912 159792
rect 144828 159740 144880 159792
rect 144920 159740 144972 159792
rect 146484 159740 146536 159792
rect 146668 159740 146720 159792
rect 153292 159740 153344 159792
rect 153476 159740 153528 159792
rect 180708 159808 180760 159860
rect 184572 159808 184624 159860
rect 259644 159808 259696 159860
rect 261944 159808 261996 159860
rect 318984 159808 319036 159860
rect 320824 159808 320876 159860
rect 356060 159808 356112 159860
rect 177856 159740 177908 159792
rect 254308 159740 254360 159792
rect 255228 159740 255280 159792
rect 313372 159740 313424 159792
rect 314108 159740 314160 159792
rect 355968 159740 356020 159792
rect 18880 159672 18932 159724
rect 109132 159672 109184 159724
rect 113088 159672 113140 159724
rect 126428 159672 126480 159724
rect 126520 159672 126572 159724
rect 156328 159672 156380 159724
rect 49976 159604 50028 159656
rect 143264 159604 143316 159656
rect 143356 159604 143408 159656
rect 156420 159604 156472 159656
rect 43260 159536 43312 159588
rect 137100 159536 137152 159588
rect 137284 159536 137336 159588
rect 139860 159536 139912 159588
rect 139952 159536 140004 159588
rect 164148 159672 164200 159724
rect 167736 159672 167788 159724
rect 246672 159672 246724 159724
rect 250996 159672 251048 159724
rect 310612 159672 310664 159724
rect 315764 159672 315816 159724
rect 359740 159808 359792 159860
rect 376300 159808 376352 159860
rect 405924 159808 405976 159860
rect 449532 159808 449584 159860
rect 459560 159808 459612 159860
rect 461308 159808 461360 159860
rect 468024 159808 468076 159860
rect 478972 159808 479024 159860
rect 484584 159808 484636 159860
rect 357808 159740 357860 159792
rect 365352 159740 365404 159792
rect 365444 159740 365496 159792
rect 395160 159740 395212 159792
rect 396540 159740 396592 159792
rect 413744 159740 413796 159792
rect 420920 159740 420972 159792
rect 440424 159740 440476 159792
rect 453764 159740 453816 159792
rect 464988 159740 465040 159792
rect 471428 159740 471480 159792
rect 478420 159740 478472 159792
rect 369584 159672 369636 159724
rect 400680 159672 400732 159724
rect 407488 159672 407540 159724
rect 429568 159672 429620 159724
rect 450360 159672 450412 159724
rect 462228 159672 462280 159724
rect 468852 159672 468904 159724
rect 474832 159672 474884 159724
rect 156788 159604 156840 159656
rect 160100 159604 160152 159656
rect 161020 159604 161072 159656
rect 241428 159604 241480 159656
rect 244280 159604 244332 159656
rect 297824 159604 297876 159656
rect 157616 159536 157668 159588
rect 238944 159536 238996 159588
rect 241796 159536 241848 159588
rect 303068 159604 303120 159656
rect 309048 159604 309100 159656
rect 354864 159604 354916 159656
rect 356152 159604 356204 159656
rect 359648 159604 359700 159656
rect 362868 159604 362920 159656
rect 395252 159604 395304 159656
rect 399024 159604 399076 159656
rect 408592 159604 408644 159656
rect 410800 159604 410852 159656
rect 432144 159604 432196 159656
rect 451188 159604 451240 159656
rect 461860 159604 461912 159656
rect 476120 159604 476172 159656
rect 482284 159604 482336 159656
rect 487436 159604 487488 159656
rect 302332 159536 302384 159588
rect 347136 159536 347188 159588
rect 347780 159536 347832 159588
rect 36544 159468 36596 159520
rect 126336 159468 126388 159520
rect 126428 159468 126480 159520
rect 127624 159468 127676 159520
rect 129924 159468 129976 159520
rect 141884 159468 141936 159520
rect 144184 159468 144236 159520
rect 225144 159468 225196 159520
rect 231676 159468 231728 159520
rect 295524 159468 295576 159520
rect 295616 159468 295668 159520
rect 335912 159468 335964 159520
rect 336096 159468 336148 159520
rect 339132 159468 339184 159520
rect 339316 159468 339368 159520
rect 349804 159468 349856 159520
rect 351920 159536 351972 159588
rect 385500 159536 385552 159588
rect 389824 159536 389876 159588
rect 413836 159536 413888 159588
rect 414204 159536 414256 159588
rect 434812 159536 434864 159588
rect 452016 159536 452068 159588
rect 463608 159536 463660 159588
rect 470508 159536 470560 159588
rect 472256 159536 472308 159588
rect 479064 159536 479116 159588
rect 479800 159536 479852 159588
rect 484768 159536 484820 159588
rect 359464 159468 359516 159520
rect 32312 159400 32364 159452
rect 6276 159332 6328 159384
rect 122748 159332 122800 159384
rect 123116 159400 123168 159452
rect 147404 159400 147456 159452
rect 150900 159400 150952 159452
rect 233792 159400 233844 159452
rect 234988 159400 235040 159452
rect 298008 159400 298060 159452
rect 301504 159400 301556 159452
rect 348792 159400 348844 159452
rect 348976 159400 349028 159452
rect 353852 159400 353904 159452
rect 355968 159400 356020 159452
rect 357992 159400 358044 159452
rect 358636 159400 358688 159452
rect 392400 159468 392452 159520
rect 424324 159468 424376 159520
rect 442448 159468 442500 159520
rect 446128 159468 446180 159520
rect 456800 159468 456852 159520
rect 458732 159468 458784 159520
rect 465080 159468 465132 159520
rect 469680 159468 469732 159520
rect 477408 159468 477460 159520
rect 478144 159468 478196 159520
rect 483664 159468 483716 159520
rect 518348 159468 518400 159520
rect 522672 159468 522724 159520
rect 359648 159400 359700 159452
rect 390744 159400 390796 159452
rect 400772 159400 400824 159452
rect 424508 159400 424560 159452
rect 427636 159400 427688 159452
rect 445024 159400 445076 159452
rect 447876 159400 447928 159452
rect 460112 159400 460164 159452
rect 462136 159400 462188 159452
rect 467840 159400 467892 159452
rect 477316 159400 477368 159452
rect 483296 159400 483348 159452
rect 126888 159332 126940 159384
rect 126980 159332 127032 159384
rect 130660 159332 130712 159384
rect 133144 159332 133196 159384
rect 137376 159332 137428 159384
rect 137468 159332 137520 159384
rect 223580 159332 223632 159384
rect 224960 159332 225012 159384
rect 290280 159332 290332 159384
rect 294788 159332 294840 159384
rect 343456 159332 343508 159384
rect 346032 159332 346084 159384
rect 73528 159264 73580 159316
rect 80060 159264 80112 159316
rect 83648 159264 83700 159316
rect 167000 159264 167052 159316
rect 170220 159264 170272 159316
rect 199292 159264 199344 159316
rect 201408 159264 201460 159316
rect 213092 159264 213144 159316
rect 214012 159264 214064 159316
rect 282000 159264 282052 159316
rect 282092 159264 282144 159316
rect 327448 159264 327500 159316
rect 327540 159264 327592 159316
rect 330576 159264 330628 159316
rect 330668 159264 330720 159316
rect 333336 159264 333388 159316
rect 333520 159264 333572 159316
rect 339040 159264 339092 159316
rect 339132 159264 339184 159316
rect 374092 159264 374144 159316
rect 80244 159196 80296 159248
rect 91100 159196 91152 159248
rect 100484 159196 100536 159248
rect 184664 159196 184716 159248
rect 187056 159196 187108 159248
rect 214104 159196 214156 159248
rect 218244 159196 218296 159248
rect 285128 159196 285180 159248
rect 287980 159196 288032 159248
rect 86960 159128 87012 159180
rect 169944 159128 169996 159180
rect 171140 159128 171192 159180
rect 172520 159128 172572 159180
rect 173624 159128 173676 159180
rect 197360 159128 197412 159180
rect 203892 159128 203944 159180
rect 213644 159128 213696 159180
rect 220728 159128 220780 159180
rect 283012 159128 283064 159180
rect 284668 159128 284720 159180
rect 285772 159128 285824 159180
rect 93676 159060 93728 159112
rect 166264 159060 166316 159112
rect 107200 158992 107252 159044
rect 183468 159060 183520 159112
rect 193772 159060 193824 159112
rect 218060 159060 218112 159112
rect 224132 159060 224184 159112
rect 288348 159128 288400 159180
rect 288900 159128 288952 159180
rect 333520 159128 333572 159180
rect 335912 159196 335964 159248
rect 342444 159196 342496 159248
rect 342720 159196 342772 159248
rect 343824 159196 343876 159248
rect 347136 159196 347188 159248
rect 349344 159196 349396 159248
rect 349804 159196 349856 159248
rect 374736 159332 374788 159384
rect 385868 159332 385920 159384
rect 388996 159332 389048 159384
rect 403900 159332 403952 159384
rect 417516 159332 417568 159384
rect 437664 159332 437716 159384
rect 448704 159332 448756 159384
rect 461124 159332 461176 159384
rect 463792 159332 463844 159384
rect 471704 159332 471756 159384
rect 518716 159332 518768 159384
rect 523500 159332 523552 159384
rect 378048 159264 378100 159316
rect 388352 159264 388404 159316
rect 404084 159264 404136 159316
rect 426992 159264 427044 159316
rect 454592 159264 454644 159316
rect 465448 159264 465500 159316
rect 465540 159264 465592 159316
rect 472256 159264 472308 159316
rect 338396 159128 338448 159180
rect 341892 159128 341944 159180
rect 373632 159128 373684 159180
rect 382740 159196 382792 159248
rect 385592 159196 385644 159248
rect 399576 159196 399628 159248
rect 457904 159196 457956 159248
rect 468116 159196 468168 159248
rect 377588 159128 377640 159180
rect 392308 159128 392360 159180
rect 404268 159128 404320 159180
rect 457076 159128 457128 159180
rect 467932 159128 467984 159180
rect 297824 159060 297876 159112
rect 305184 159060 305236 159112
rect 307392 159060 307444 159112
rect 174360 158992 174412 159044
rect 176660 158992 176712 159044
rect 183744 158992 183796 159044
rect 200488 158992 200540 159044
rect 200580 158992 200632 159044
rect 224960 158992 225012 159044
rect 230848 158992 230900 159044
rect 294788 158992 294840 159044
rect 298100 158992 298152 159044
rect 299940 158992 299992 159044
rect 308220 158992 308272 159044
rect 348976 158992 349028 159044
rect 351092 159060 351144 159112
rect 382372 159060 382424 159112
rect 395712 159060 395764 159112
rect 405648 159060 405700 159112
rect 412548 159060 412600 159112
rect 413928 159060 413980 159112
rect 459652 159060 459704 159112
rect 466460 159060 466512 159112
rect 353208 158992 353260 159044
rect 356060 158992 356112 159044
rect 96252 158924 96304 158976
rect 121644 158924 121696 158976
rect 124036 158924 124088 158976
rect 194508 158924 194560 158976
rect 194692 158924 194744 158976
rect 203708 158924 203760 158976
rect 208124 158924 208176 158976
rect 212448 158924 212500 158976
rect 102968 158788 103020 158840
rect 125508 158856 125560 158908
rect 127348 158856 127400 158908
rect 127992 158856 128044 158908
rect 130752 158856 130804 158908
rect 194968 158856 195020 158908
rect 90364 158720 90416 158772
rect 92480 158720 92532 158772
rect 92848 158720 92900 158772
rect 113824 158788 113876 158840
rect 109684 158720 109736 158772
rect 133144 158788 133196 158840
rect 133236 158788 133288 158840
rect 158720 158788 158772 158840
rect 163504 158788 163556 158840
rect 196072 158788 196124 158840
rect 207296 158788 207348 158840
rect 231032 158924 231084 158976
rect 237564 158924 237616 158976
rect 300032 158924 300084 158976
rect 217324 158856 217376 158908
rect 220728 158856 220780 158908
rect 248512 158856 248564 158908
rect 314936 158924 314988 158976
rect 358728 158924 358780 158976
rect 359464 158992 359516 159044
rect 378784 158992 378836 159044
rect 383108 158992 383160 159044
rect 411444 158992 411496 159044
rect 462964 158992 463016 159044
rect 469220 158992 469272 159044
rect 473912 158992 473964 159044
rect 480260 158992 480312 159044
rect 363512 158924 363564 158976
rect 305644 158856 305696 158908
rect 307668 158856 307720 158908
rect 308220 158856 308272 158908
rect 310704 158856 310756 158908
rect 311992 158856 312044 158908
rect 312452 158856 312504 158908
rect 313464 158856 313516 158908
rect 319168 158856 319220 158908
rect 322848 158856 322900 158908
rect 364800 158924 364852 158976
rect 365352 158924 365404 158976
rect 371884 158924 371936 158976
rect 374552 158924 374604 158976
rect 386328 158924 386380 158976
rect 391480 158924 391532 158976
rect 394608 158924 394660 158976
rect 409144 158924 409196 158976
rect 410892 158924 410944 158976
rect 420092 158924 420144 158976
rect 423588 158924 423640 158976
rect 460480 158924 460532 158976
rect 466552 158924 466604 158976
rect 475568 158924 475620 158976
rect 481732 158924 481784 158976
rect 214840 158788 214892 158840
rect 221740 158788 221792 158840
rect 238392 158788 238444 158840
rect 242808 158788 242860 158840
rect 261116 158788 261168 158840
rect 316960 158788 317012 158840
rect 322480 158788 322532 158840
rect 118976 158720 119028 158772
rect 119620 158720 119672 158772
rect 119804 158720 119856 158772
rect 147404 158720 147456 158772
rect 147496 158720 147548 158772
rect 149060 158720 149112 158772
rect 153292 158720 153344 158772
rect 174360 158720 174412 158772
rect 174452 158720 174504 158772
rect 174912 158720 174964 158772
rect 180340 158720 180392 158772
rect 204904 158720 204956 158772
rect 210608 158720 210660 158772
rect 215300 158720 215352 158772
rect 221556 158720 221608 158772
rect 223856 158720 223908 158772
rect 240876 158720 240928 158772
rect 243360 158720 243412 158772
rect 254400 158720 254452 158772
rect 255320 158720 255372 158772
rect 258540 158720 258592 158772
rect 260932 158720 260984 158772
rect 264428 158720 264480 158772
rect 267096 158720 267148 158772
rect 267832 158720 267884 158772
rect 320272 158720 320324 158772
rect 321652 158720 321704 158772
rect 361120 158788 361172 158840
rect 361212 158788 361264 158840
rect 330576 158720 330628 158772
rect 367192 158720 367244 158772
rect 81072 158652 81124 158704
rect 180800 158652 180852 158704
rect 180892 158652 180944 158704
rect 181904 158652 181956 158704
rect 181996 158652 182048 158704
rect 257528 158652 257580 158704
rect 371884 158788 371936 158840
rect 374828 158788 374880 158840
rect 384764 158856 384816 158908
rect 389180 158856 389232 158908
rect 405740 158856 405792 158908
rect 409328 158856 409380 158908
rect 416688 158856 416740 158908
rect 419632 158856 419684 158908
rect 452844 158856 452896 158908
rect 464252 158856 464304 158908
rect 466368 158856 466420 158908
rect 472348 158856 472400 158908
rect 474740 158856 474792 158908
rect 480996 158856 481048 158908
rect 508688 158856 508740 158908
rect 510068 158856 510120 158908
rect 367928 158720 367980 158772
rect 374736 158720 374788 158772
rect 383660 158788 383712 158840
rect 387892 158788 387944 158840
rect 388076 158788 388128 158840
rect 390376 158788 390428 158840
rect 456248 158788 456300 158840
rect 466828 158788 466880 158840
rect 476396 158788 476448 158840
rect 482376 158788 482428 158840
rect 506388 158788 506440 158840
rect 507584 158788 507636 158840
rect 413376 158720 413428 158772
rect 419724 158720 419776 158772
rect 464620 158720 464672 158772
rect 471244 158720 471296 158772
rect 473084 158720 473136 158772
rect 479708 158720 479760 158772
rect 481456 158720 481508 158772
rect 486148 158720 486200 158772
rect 504088 158720 504140 158772
rect 505008 158720 505060 158772
rect 506204 158720 506256 158772
rect 506756 158720 506808 158772
rect 507492 158720 507544 158772
rect 508412 158720 508464 158772
rect 509976 158720 510028 158772
rect 511724 158720 511776 158772
rect 515128 158720 515180 158772
rect 518532 158720 518584 158772
rect 374552 158652 374604 158704
rect 74356 158584 74408 158636
rect 175188 158584 175240 158636
rect 175280 158584 175332 158636
rect 252560 158584 252612 158636
rect 71044 158516 71096 158568
rect 172704 158516 172756 158568
rect 178684 158516 178736 158568
rect 255412 158516 255464 158568
rect 361120 158516 361172 158568
rect 362960 158516 363012 158568
rect 67640 158448 67692 158500
rect 170220 158448 170272 158500
rect 171968 158448 172020 158500
rect 249800 158448 249852 158500
rect 60924 158380 60976 158432
rect 165068 158380 165120 158432
rect 165252 158380 165304 158432
rect 244648 158380 244700 158432
rect 64236 158312 64288 158364
rect 167552 158312 167604 158364
rect 168564 158312 168616 158364
rect 247224 158312 247276 158364
rect 54208 158244 54260 158296
rect 160284 158244 160336 158296
rect 161848 158244 161900 158296
rect 242072 158244 242124 158296
rect 50804 158176 50856 158228
rect 157340 158176 157392 158228
rect 158444 158176 158496 158228
rect 239680 158176 239732 158228
rect 256884 158176 256936 158228
rect 314752 158176 314804 158228
rect 47492 158108 47544 158160
rect 154764 158108 154816 158160
rect 155132 158108 155184 158160
rect 237380 158108 237432 158160
rect 246764 158108 246816 158160
rect 306932 158108 306984 158160
rect 37372 158040 37424 158092
rect 147128 158040 147180 158092
rect 148416 158040 148468 158092
rect 231860 158040 231912 158092
rect 243452 158040 243504 158092
rect 304356 158040 304408 158092
rect 388 157972 440 158024
rect 118884 157972 118936 158024
rect 122748 157972 122800 158024
rect 123392 157972 123444 158024
rect 131580 157972 131632 158024
rect 218980 157972 219032 158024
rect 236736 157972 236788 158024
rect 299572 157972 299624 158024
rect 77760 157904 77812 157956
rect 84476 157836 84528 157888
rect 175924 157836 175976 157888
rect 176200 157904 176252 157956
rect 182824 157904 182876 157956
rect 185400 157904 185452 157956
rect 260196 157904 260248 157956
rect 178040 157836 178092 157888
rect 181536 157836 181588 157888
rect 188160 157836 188212 157888
rect 188804 157836 188856 157888
rect 262680 157836 262732 157888
rect 87788 157768 87840 157820
rect 181628 157768 181680 157820
rect 181812 157768 181864 157820
rect 190644 157768 190696 157820
rect 195520 157768 195572 157820
rect 267740 157768 267792 157820
rect 91192 157700 91244 157752
rect 181260 157700 181312 157752
rect 181904 157700 181956 157752
rect 94596 157632 94648 157684
rect 181536 157632 181588 157684
rect 181720 157632 181772 157684
rect 185584 157632 185636 157684
rect 190460 157700 190512 157752
rect 264060 157700 264112 157752
rect 236092 157632 236144 157684
rect 97908 157564 97960 157616
rect 193220 157564 193272 157616
rect 197360 157564 197412 157616
rect 251272 157564 251324 157616
rect 111340 157496 111392 157548
rect 203432 157496 203484 157548
rect 204904 157496 204956 157548
rect 256332 157496 256384 157548
rect 114744 157428 114796 157480
rect 206192 157428 206244 157480
rect 141700 157360 141752 157412
rect 226708 157360 226760 157412
rect 49148 157292 49200 157344
rect 156052 157292 156104 157344
rect 156328 157292 156380 157344
rect 212540 157292 212592 157344
rect 213184 157292 213236 157344
rect 281632 157292 281684 157344
rect 45744 157224 45796 157276
rect 153476 157224 153528 157276
rect 192116 157224 192168 157276
rect 265164 157224 265216 157276
rect 39028 157156 39080 157208
rect 148232 157156 148284 157208
rect 160100 157156 160152 157208
rect 164056 157156 164108 157208
rect 164148 157156 164200 157208
rect 171600 157156 171652 157208
rect 177028 157156 177080 157208
rect 254032 157156 254084 157208
rect 290556 157156 290608 157208
rect 339960 157156 340012 157208
rect 42432 157088 42484 157140
rect 150900 157088 150952 157140
rect 151728 157088 151780 157140
rect 234620 157088 234672 157140
rect 287152 157088 287204 157140
rect 338120 157088 338172 157140
rect 35716 157020 35768 157072
rect 24768 156952 24820 157004
rect 137560 156952 137612 157004
rect 145012 157020 145064 157072
rect 229284 157020 229336 157072
rect 231032 157020 231084 157072
rect 276848 157020 276900 157072
rect 280436 157020 280488 157072
rect 332692 157020 332744 157072
rect 146024 156952 146076 157004
rect 150072 156952 150124 157004
rect 233240 156952 233292 157004
rect 283840 156952 283892 157004
rect 335452 156952 335504 157004
rect 18052 156884 18104 156936
rect 132500 156884 132552 156936
rect 138296 156884 138348 156936
rect 224132 156884 224184 156936
rect 273720 156884 273772 156936
rect 327540 156884 327592 156936
rect 21364 156816 21416 156868
rect 135260 156816 135312 156868
rect 135812 156816 135864 156868
rect 222200 156816 222252 156868
rect 224960 156816 225012 156868
rect 271972 156816 272024 156868
rect 277124 156816 277176 156868
rect 330024 156816 330076 156868
rect 11244 156748 11296 156800
rect 127164 156748 127216 156800
rect 139124 156748 139176 156800
rect 225052 156748 225104 156800
rect 226616 156748 226668 156800
rect 291568 156748 291620 156800
rect 297272 156748 297324 156800
rect 345572 156748 345624 156800
rect 14648 156680 14700 156732
rect 129832 156680 129884 156732
rect 134892 156680 134944 156732
rect 221372 156680 221424 156732
rect 230020 156680 230072 156732
rect 294052 156680 294104 156732
rect 300676 156680 300728 156732
rect 348056 156680 348108 156732
rect 2044 156612 2096 156664
rect 120172 156612 120224 156664
rect 128176 156612 128228 156664
rect 216680 156612 216732 156664
rect 223212 156612 223264 156664
rect 288992 156612 289044 156664
rect 293868 156612 293920 156664
rect 342260 156612 342312 156664
rect 52460 156544 52512 156596
rect 158628 156544 158680 156596
rect 158720 156544 158772 156596
rect 219992 156544 220044 156596
rect 59268 156476 59320 156528
rect 163780 156476 163832 156528
rect 164056 156476 164108 156528
rect 69296 156408 69348 156460
rect 164148 156408 164200 156460
rect 164332 156476 164384 156528
rect 225512 156476 225564 156528
rect 227996 156408 228048 156460
rect 82820 156340 82872 156392
rect 181812 156340 181864 156392
rect 198832 156340 198884 156392
rect 200948 156340 201000 156392
rect 209780 156340 209832 156392
rect 278872 156340 278924 156392
rect 101312 156272 101364 156324
rect 196164 156272 196216 156324
rect 200764 156272 200816 156324
rect 211344 156272 211396 156324
rect 212540 156272 212592 156324
rect 215392 156272 215444 156324
rect 216496 156272 216548 156324
rect 283472 156272 283524 156324
rect 99564 156204 99616 156256
rect 194692 156204 194744 156256
rect 108028 156136 108080 156188
rect 200672 156136 200724 156188
rect 118148 156068 118200 156120
rect 203064 156204 203116 156256
rect 208768 156136 208820 156188
rect 200948 156068 201000 156120
rect 219900 156204 219952 156256
rect 285680 156204 285732 156256
rect 218060 156136 218112 156188
rect 266544 156136 266596 156188
rect 121460 156000 121512 156052
rect 200764 156000 200816 156052
rect 202236 156000 202288 156052
rect 214288 156000 214340 156052
rect 124864 155932 124916 155984
rect 213920 155932 213972 155984
rect 273536 156068 273588 156120
rect 214564 156000 214616 156052
rect 273260 156000 273312 156052
rect 270500 155932 270552 155984
rect 89536 155864 89588 155916
rect 186964 155864 187016 155916
rect 192944 155864 192996 155916
rect 265900 155864 265952 155916
rect 293040 155864 293092 155916
rect 342352 155864 342404 155916
rect 53380 155796 53432 155848
rect 66720 155796 66772 155848
rect 66812 155796 66864 155848
rect 82912 155796 82964 155848
rect 88708 155796 88760 155848
rect 186412 155796 186464 155848
rect 189632 155796 189684 155848
rect 263692 155796 263744 155848
rect 296444 155796 296496 155848
rect 345112 155796 345164 155848
rect 12164 155728 12216 155780
rect 109776 155728 109828 155780
rect 112260 155728 112312 155780
rect 204352 155728 204404 155780
rect 206468 155728 206520 155780
rect 276112 155728 276164 155780
rect 289728 155728 289780 155780
rect 339592 155728 339644 155780
rect 60096 155660 60148 155712
rect 78864 155660 78916 155712
rect 81900 155660 81952 155712
rect 181168 155660 181220 155712
rect 186228 155660 186280 155712
rect 260840 155660 260892 155712
rect 267004 155660 267056 155712
rect 322112 155660 322164 155712
rect 340972 155660 341024 155712
rect 378692 155660 378744 155712
rect 46572 155592 46624 155644
rect 75092 155592 75144 155644
rect 75184 155592 75236 155644
rect 176016 155592 176068 155644
rect 179512 155592 179564 155644
rect 255596 155592 255648 155644
rect 270316 155592 270368 155644
rect 324964 155592 325016 155644
rect 344376 155592 344428 155644
rect 381452 155592 381504 155644
rect 39856 155524 39908 155576
rect 68928 155524 68980 155576
rect 71872 155524 71924 155576
rect 173072 155524 173124 155576
rect 176292 155524 176344 155576
rect 253020 155524 253072 155576
rect 263600 155524 263652 155576
rect 320180 155524 320232 155576
rect 337660 155524 337712 155576
rect 376300 155524 376352 155576
rect 65156 155456 65208 155508
rect 168380 155456 168432 155508
rect 169392 155456 169444 155508
rect 247960 155456 248012 155508
rect 260288 155456 260340 155508
rect 317512 155456 317564 155508
rect 333428 155456 333480 155508
rect 373080 155456 373132 155508
rect 4528 155388 4580 155440
rect 122012 155388 122064 155440
rect 122288 155388 122340 155440
rect 211988 155388 212040 155440
rect 214104 155388 214156 155440
rect 261392 155388 261444 155440
rect 330116 155388 330168 155440
rect 370596 155388 370648 155440
rect 7932 155320 7984 155372
rect 124588 155320 124640 155372
rect 142528 155320 142580 155372
rect 227812 155320 227864 155372
rect 253572 155320 253624 155372
rect 312084 155320 312136 155372
rect 319996 155320 320048 155372
rect 363052 155320 363104 155372
rect 8760 155252 8812 155304
rect 125600 155252 125652 155304
rect 129004 155252 129056 155304
rect 217048 155252 217100 155304
rect 233332 155252 233384 155304
rect 296812 155252 296864 155304
rect 299756 155252 299808 155304
rect 347780 155252 347832 155304
rect 373816 155252 373868 155304
rect 403532 155252 403584 155304
rect 5356 155184 5408 155236
rect 122932 155184 122984 155236
rect 125692 155184 125744 155236
rect 214472 155184 214524 155236
rect 240048 155184 240100 155236
rect 302332 155184 302384 155236
rect 303160 155184 303212 155236
rect 350080 155184 350132 155236
rect 370412 155184 370464 155236
rect 401692 155184 401744 155236
rect 92020 155116 92072 155168
rect 189080 155116 189132 155168
rect 189172 155116 189224 155168
rect 194048 155116 194100 155168
rect 196348 155116 196400 155168
rect 268476 155116 268528 155168
rect 306564 155116 306616 155168
rect 352472 155116 352524 155168
rect 95424 155048 95476 155100
rect 98736 154980 98788 155032
rect 186320 154980 186372 155032
rect 186780 155048 186832 155100
rect 191472 154980 191524 155032
rect 199660 155048 199712 155100
rect 271052 155048 271104 155100
rect 200120 154980 200172 155032
rect 207112 154980 207164 155032
rect 269212 154980 269264 155032
rect 15476 154912 15528 154964
rect 109040 154912 109092 154964
rect 110512 154912 110564 154964
rect 139308 154912 139360 154964
rect 145932 154912 145984 154964
rect 230020 154912 230072 154964
rect 250168 154912 250220 154964
rect 309508 154912 309560 154964
rect 106372 154844 106424 154896
rect 186596 154844 186648 154896
rect 186688 154844 186740 154896
rect 245936 154844 245988 154896
rect 109132 154776 109184 154828
rect 133052 154776 133104 154828
rect 149244 154776 149296 154828
rect 232504 154776 232556 154828
rect 155960 154708 156012 154760
rect 237656 154708 237708 154760
rect 162676 154640 162728 154692
rect 242900 154640 242952 154692
rect 154488 154572 154540 154624
rect 51632 154504 51684 154556
rect 154948 154504 155000 154556
rect 159364 154572 159416 154624
rect 240232 154572 240284 154624
rect 156420 154504 156472 154556
rect 156604 154504 156656 154556
rect 212724 154504 212776 154556
rect 219348 154504 219400 154556
rect 286232 154504 286284 154556
rect 286324 154504 286376 154556
rect 337200 154504 337252 154556
rect 353668 154504 353720 154556
rect 388628 154504 388680 154556
rect 44916 154436 44968 154488
rect 142528 154436 142580 154488
rect 142620 154436 142672 154488
rect 191012 154436 191064 154488
rect 41604 154368 41656 154420
rect 142804 154368 142856 154420
rect 142896 154368 142948 154420
rect 113824 154300 113876 154352
rect 181076 154300 181128 154352
rect 181444 154368 181496 154420
rect 189540 154368 189592 154420
rect 202420 154436 202472 154488
rect 208952 154436 209004 154488
rect 278136 154436 278188 154488
rect 279976 154436 280028 154488
rect 332140 154436 332192 154488
rect 350264 154436 350316 154488
rect 386052 154436 386104 154488
rect 191196 154368 191248 154420
rect 258264 154368 258316 154420
rect 266176 154368 266228 154420
rect 321836 154368 321888 154420
rect 346860 154368 346912 154420
rect 383660 154368 383712 154420
rect 390652 154368 390704 154420
rect 416872 154368 416924 154420
rect 191380 154300 191432 154352
rect 201776 154300 201828 154352
rect 205548 154300 205600 154352
rect 275560 154300 275612 154352
rect 276204 154300 276256 154352
rect 329840 154300 329892 154352
rect 340144 154300 340196 154352
rect 378324 154300 378376 154352
rect 387616 154300 387668 154352
rect 414296 154300 414348 154352
rect 38476 154232 38528 154284
rect 23940 154164 23992 154216
rect 27252 154096 27304 154148
rect 132592 154096 132644 154148
rect 13820 154028 13872 154080
rect 129188 154028 129240 154080
rect 132868 154164 132920 154216
rect 133144 154164 133196 154216
rect 142620 154164 142672 154216
rect 139492 154096 139544 154148
rect 139584 154096 139636 154148
rect 142344 154096 142396 154148
rect 147680 154232 147732 154284
rect 156604 154232 156656 154284
rect 172796 154232 172848 154284
rect 250536 154232 250588 154284
rect 256056 154232 256108 154284
rect 314108 154232 314160 154284
rect 343548 154232 343600 154284
rect 380900 154232 380952 154284
rect 383936 154232 383988 154284
rect 411720 154232 411772 154284
rect 142804 154164 142856 154216
rect 150440 154164 150492 154216
rect 152556 154164 152608 154216
rect 147496 154096 147548 154148
rect 147588 154096 147640 154148
rect 156328 154096 156380 154148
rect 156788 154164 156840 154216
rect 163228 154164 163280 154216
rect 166080 154164 166132 154216
rect 245660 154164 245712 154216
rect 249708 154164 249760 154216
rect 309232 154164 309284 154216
rect 326712 154164 326764 154216
rect 368020 154164 368072 154216
rect 380808 154164 380860 154216
rect 409236 154164 409288 154216
rect 136916 154028 136968 154080
rect 137376 154028 137428 154080
rect 142896 154028 142948 154080
rect 10416 153960 10468 154012
rect 126612 153960 126664 154012
rect 127624 153960 127676 154012
rect 142436 153960 142488 154012
rect 142528 153960 142580 154012
rect 153200 154028 153252 154080
rect 154948 154028 155000 154080
rect 158076 154028 158128 154080
rect 160192 154096 160244 154148
rect 240968 154096 241020 154148
rect 242624 154096 242676 154148
rect 303804 154096 303856 154148
rect 323308 154096 323360 154148
rect 365720 154096 365772 154148
rect 367100 154096 367152 154148
rect 398840 154096 398892 154148
rect 401600 154096 401652 154148
rect 425336 154096 425388 154148
rect 235172 154028 235224 154080
rect 235908 154028 235960 154080
rect 298744 154028 298796 154080
rect 316592 154028 316644 154080
rect 360384 154028 360436 154080
rect 363696 154028 363748 154080
rect 396356 154028 396408 154080
rect 398196 154028 398248 154080
rect 422668 154028 422720 154080
rect 143080 153960 143132 154012
rect 222936 153960 222988 154012
rect 7104 153892 7156 153944
rect 124220 153892 124272 153944
rect 125508 153892 125560 153944
rect 133144 153892 133196 153944
rect 133236 153892 133288 153944
rect 219716 153892 219768 153944
rect 222384 153892 222436 153944
rect 288440 153960 288492 154012
rect 313280 153960 313332 154012
rect 357808 153960 357860 154012
rect 360476 153960 360528 154012
rect 393780 153960 393832 154012
rect 397368 153960 397420 154012
rect 422300 153960 422352 154012
rect 225788 153892 225840 153944
rect 291200 153892 291252 153944
rect 309876 153892 309928 153944
rect 355232 153892 355284 153944
rect 357348 153892 357400 153944
rect 391204 153892 391256 153944
rect 393964 153892 394016 153944
rect 419540 153892 419592 153944
rect 1216 153824 1268 153876
rect 119528 153824 119580 153876
rect 119620 153824 119672 153876
rect 209780 153824 209832 153876
rect 215668 153824 215720 153876
rect 283288 153824 283340 153876
rect 283380 153824 283432 153876
rect 334624 153824 334676 153876
rect 336832 153824 336884 153876
rect 375748 153824 375800 153876
rect 377220 153824 377272 153876
rect 406568 153824 406620 153876
rect 48320 153756 48372 153808
rect 155500 153756 155552 153808
rect 156420 153756 156472 153808
rect 218060 153756 218112 153808
rect 232596 153756 232648 153808
rect 296168 153756 296220 153808
rect 435180 153756 435232 153808
rect 442908 153756 442960 153808
rect 61752 153688 61804 153740
rect 165804 153688 165856 153740
rect 58348 153620 58400 153672
rect 156512 153620 156564 153672
rect 156604 153620 156656 153672
rect 210148 153688 210200 153740
rect 229100 153688 229152 153740
rect 293592 153688 293644 153740
rect 176660 153620 176712 153672
rect 79416 153552 79468 153604
rect 179420 153552 179472 153604
rect 182916 153620 182968 153672
rect 191196 153620 191248 153672
rect 191288 153620 191340 153672
rect 195980 153620 196032 153672
rect 196072 153620 196124 153672
rect 238392 153620 238444 153672
rect 239220 153620 239272 153672
rect 301320 153620 301372 153672
rect 230664 153552 230716 153604
rect 246028 153552 246080 153604
rect 306380 153552 306432 153604
rect 102140 153484 102192 153536
rect 196624 153484 196676 153536
rect 196716 153484 196768 153536
rect 105452 153416 105504 153468
rect 197268 153416 197320 153468
rect 200488 153484 200540 153536
rect 258908 153484 258960 153536
rect 262772 153484 262824 153536
rect 319260 153484 319312 153536
rect 108856 153348 108908 153400
rect 191380 153348 191432 153400
rect 191748 153348 191800 153400
rect 195888 153348 195940 153400
rect 195980 153348 196032 153400
rect 197360 153348 197412 153400
rect 197636 153416 197688 153468
rect 199200 153416 199252 153468
rect 199292 153416 199344 153468
rect 248604 153416 248656 153468
rect 252652 153416 252704 153468
rect 311532 153416 311584 153468
rect 243452 153348 243504 153400
rect 259460 153348 259512 153400
rect 316776 153348 316828 153400
rect 116400 153280 116452 153332
rect 207572 153280 207624 153332
rect 272892 153280 272944 153332
rect 327080 153280 327132 153332
rect 34796 153212 34848 153264
rect 142344 153212 142396 153264
rect 142436 153212 142488 153264
rect 204996 153212 205048 153264
rect 269488 153212 269540 153264
rect 324412 153212 324464 153264
rect 66720 153144 66772 153196
rect 159364 153144 159416 153196
rect 172520 153144 172572 153196
rect 249248 153144 249300 153196
rect 255320 153144 255372 153196
rect 312820 153144 312872 153196
rect 316960 153144 317012 153196
rect 317972 153144 318024 153196
rect 318616 153144 318668 153196
rect 30196 153076 30248 153128
rect 109592 153076 109644 153128
rect 109868 153076 109920 153128
rect 197912 153076 197964 153128
rect 203708 153076 203760 153128
rect 266912 153076 266964 153128
rect 267096 153076 267148 153128
rect 320456 153076 320508 153128
rect 320640 153144 320692 153196
rect 361028 153144 361080 153196
rect 366272 153144 366324 153196
rect 80060 153008 80112 153060
rect 174820 153008 174872 153060
rect 174912 153008 174964 153060
rect 251824 153008 251876 153060
rect 257712 153008 257764 153060
rect 315396 153008 315448 153060
rect 317420 153008 317472 153060
rect 320640 153008 320692 153060
rect 325056 153076 325108 153128
rect 366732 153076 366784 153128
rect 367192 153144 367244 153196
rect 368664 153144 368716 153196
rect 371332 153144 371384 153196
rect 402060 153144 402112 153196
rect 397920 153076 397972 153128
rect 398104 153076 398156 153128
rect 407856 153144 407908 153196
rect 415308 153144 415360 153196
rect 435456 153144 435508 153196
rect 437756 153144 437808 153196
rect 452844 153144 452896 153196
rect 456800 153144 456852 153196
rect 459192 153144 459244 153196
rect 461860 153144 461912 153196
rect 463056 153144 463108 153196
rect 466460 153144 466512 153196
rect 469496 153144 469548 153196
rect 471244 153144 471296 153196
rect 473544 153144 473596 153196
rect 474832 153144 474884 153196
rect 476580 153144 476632 153196
rect 485688 153144 485740 153196
rect 489368 153144 489420 153196
rect 492404 153144 492456 153196
rect 494520 153144 494572 153196
rect 495256 153144 495308 153196
rect 496452 153144 496504 153196
rect 496636 153144 496688 153196
rect 497740 153144 497792 153196
rect 498292 153144 498344 153196
rect 499028 153144 499080 153196
rect 500960 153144 501012 153196
rect 501604 153144 501656 153196
rect 510436 153144 510488 153196
rect 512000 153144 512052 153196
rect 512552 153144 512604 153196
rect 514852 153144 514904 153196
rect 405832 153076 405884 153128
rect 408500 153076 408552 153128
rect 411628 153076 411680 153128
rect 361672 153008 361724 153060
rect 364524 153008 364576 153060
rect 396908 153008 396960 153060
rect 407028 153008 407080 153060
rect 429200 153008 429252 153060
rect 432696 153076 432748 153128
rect 448980 153076 449032 153128
rect 466552 153076 466604 153128
rect 470140 153076 470192 153128
rect 471704 153076 471756 153128
rect 472716 153076 472768 153128
rect 473360 153076 473412 153128
rect 475292 153076 475344 153128
rect 476120 153076 476172 153128
rect 477868 153076 477920 153128
rect 484308 153076 484360 153128
rect 488172 153076 488224 153128
rect 489920 153076 489972 153128
rect 492772 153076 492824 153128
rect 493232 153076 493284 153128
rect 495440 153076 495492 153128
rect 495808 153076 495860 153128
rect 497096 153076 497148 153128
rect 511264 153076 511316 153128
rect 513472 153076 513524 153128
rect 432880 153008 432932 153060
rect 433524 153008 433576 153060
rect 449900 153008 449952 153060
rect 465080 153008 465132 153060
rect 468852 153008 468904 153060
rect 472256 153008 472308 153060
rect 474004 153008 474056 153060
rect 484860 153008 484912 153060
rect 488724 153008 488776 153060
rect 497464 153008 497516 153060
rect 498292 153008 498344 153060
rect 511724 153008 511776 153060
rect 514300 153008 514352 153060
rect 97080 152940 97132 152992
rect 192760 152940 192812 152992
rect 194968 152940 195020 152992
rect 218428 152940 218480 152992
rect 225144 152940 225196 152992
rect 228732 152940 228784 152992
rect 228824 152940 228876 152992
rect 284576 152940 284628 152992
rect 285496 152940 285548 152992
rect 336740 152940 336792 152992
rect 339500 152940 339552 152992
rect 377036 152940 377088 152992
rect 382188 152940 382240 152992
rect 410432 152940 410484 152992
rect 410892 152940 410944 152992
rect 430948 152940 431000 152992
rect 431040 152940 431092 152992
rect 447692 152940 447744 152992
rect 472348 152940 472400 152992
rect 474740 152940 474792 152992
rect 483204 152940 483256 152992
rect 487528 152940 487580 152992
rect 490748 152940 490800 152992
rect 493232 152940 493284 152992
rect 494060 152940 494112 152992
rect 495808 152940 495860 152992
rect 502892 152940 502944 152992
rect 503352 152940 503404 152992
rect 513196 152940 513248 152992
rect 515956 152940 516008 152992
rect 92480 152872 92532 152924
rect 187700 152872 187752 152924
rect 187884 152872 187936 152924
rect 262220 152872 262272 152924
rect 265348 152872 265400 152924
rect 321192 152872 321244 152924
rect 324228 152872 324280 152924
rect 366088 152872 366140 152924
rect 368756 152872 368808 152924
rect 400220 152872 400272 152924
rect 402428 152872 402480 152924
rect 425888 152872 425940 152924
rect 428464 152872 428516 152924
rect 439504 152872 439556 152924
rect 440240 152872 440292 152924
rect 441528 152872 441580 152924
rect 441988 152872 442040 152924
rect 442724 152872 442776 152924
rect 443000 152872 443052 152924
rect 445760 152872 445812 152924
rect 446956 152872 447008 152924
rect 459836 152872 459888 152924
rect 513840 152872 513892 152924
rect 516140 152872 516192 152924
rect 33140 152804 33192 152856
rect 144000 152804 144052 152856
rect 144828 152804 144880 152856
rect 161940 152804 161992 152856
rect 164424 152804 164476 152856
rect 244280 152804 244332 152856
rect 251916 152804 251968 152856
rect 310888 152804 310940 152856
rect 311992 152804 312044 152856
rect 356060 152804 356112 152856
rect 362040 152804 362092 152856
rect 395068 152804 395120 152856
rect 395160 152804 395212 152856
rect 397552 152804 397604 152856
rect 400128 152804 400180 152856
rect 423956 152804 424008 152856
rect 426256 152804 426308 152856
rect 443828 152804 443880 152856
rect 445668 152804 445720 152856
rect 458548 152804 458600 152856
rect 491576 152804 491628 152856
rect 494060 152804 494112 152856
rect 26424 152736 26476 152788
rect 138848 152736 138900 152788
rect 142344 152736 142396 152788
rect 145288 152736 145340 152788
rect 149060 152736 149112 152788
rect 231308 152736 231360 152788
rect 245108 152736 245160 152788
rect 305736 152736 305788 152788
rect 307668 152736 307720 152788
rect 352012 152736 352064 152788
rect 352748 152736 352800 152788
rect 387984 152736 388036 152788
rect 390376 152736 390428 152788
rect 414940 152736 414992 152788
rect 415860 152736 415912 152788
rect 436100 152736 436152 152788
rect 437296 152736 437348 152788
rect 28908 152668 28960 152720
rect 140780 152668 140832 152720
rect 140872 152668 140924 152720
rect 22192 152600 22244 152652
rect 135628 152600 135680 152652
rect 137100 152600 137152 152652
rect 142252 152600 142304 152652
rect 143264 152668 143316 152720
rect 156788 152668 156840 152720
rect 172428 152668 172480 152720
rect 176108 152668 176160 152720
rect 220728 152668 220780 152720
rect 228824 152668 228876 152720
rect 247684 152668 247736 152720
rect 307760 152668 307812 152720
rect 311808 152668 311860 152720
rect 356520 152668 356572 152720
rect 359556 152668 359608 152720
rect 393320 152668 393372 152720
rect 394884 152668 394936 152720
rect 420092 152668 420144 152720
rect 423404 152668 423456 152720
rect 441896 152668 441948 152720
rect 452200 152736 452252 152788
rect 444472 152668 444524 152720
rect 458180 152668 458232 152720
rect 226340 152600 226392 152652
rect 234528 152600 234580 152652
rect 297456 152600 297508 152652
rect 304816 152600 304868 152652
rect 351368 152600 351420 152652
rect 354496 152600 354548 152652
rect 389272 152600 389324 152652
rect 393136 152600 393188 152652
rect 418804 152600 418856 152652
rect 419264 152600 419316 152652
rect 438860 152600 438912 152652
rect 442816 152600 442868 152652
rect 456800 152600 456852 152652
rect 19708 152532 19760 152584
rect 133880 152532 133932 152584
rect 134064 152532 134116 152584
rect 221004 152532 221056 152584
rect 228272 152532 228324 152584
rect 292948 152532 293000 152584
rect 299388 152532 299440 152584
rect 346860 152532 346912 152584
rect 349068 152532 349120 152584
rect 385040 152532 385092 152584
rect 386420 152532 386472 152584
rect 413652 152532 413704 152584
rect 413928 152532 413980 152584
rect 433524 152532 433576 152584
rect 434628 152532 434680 152584
rect 450268 152532 450320 152584
rect 2872 152464 2924 152516
rect 120816 152464 120868 152516
rect 23296 152396 23348 152448
rect 110972 152396 111024 152448
rect 120632 152396 120684 152448
rect 210792 152464 210844 152516
rect 212448 152464 212500 152516
rect 277492 152464 277544 152516
rect 278780 152464 278832 152516
rect 121000 152396 121052 152448
rect 205640 152396 205692 152448
rect 215300 152396 215352 152448
rect 279424 152396 279476 152448
rect 279608 152464 279660 152516
rect 330852 152464 330904 152516
rect 330944 152464 330996 152516
rect 371240 152464 371292 152516
rect 372988 152464 373040 152516
rect 403348 152464 403400 152516
rect 404912 152464 404964 152516
rect 427820 152464 427872 152516
rect 430212 152464 430264 152516
rect 447140 152464 447192 152516
rect 331496 152396 331548 152448
rect 332600 152396 332652 152448
rect 372620 152396 372672 152448
rect 375472 152396 375524 152448
rect 405280 152396 405332 152448
rect 408592 152396 408644 152448
rect 417424 152396 417476 152448
rect 418436 152396 418488 152448
rect 438032 152396 438084 152448
rect 438584 152396 438636 152448
rect 453488 152396 453540 152448
rect 514484 152396 514536 152448
rect 517428 152396 517480 152448
rect 91100 152328 91152 152380
rect 179972 152328 180024 152380
rect 181260 152328 181312 152380
rect 256976 152328 257028 152380
rect 260932 152328 260984 152380
rect 316040 152328 316092 152380
rect 320272 152328 320324 152380
rect 323124 152328 323176 152380
rect 323216 152328 323268 152380
rect 330484 152328 330536 152380
rect 330576 152328 330628 152380
rect 367376 152328 367428 152380
rect 381360 152328 381412 152380
rect 409880 152328 409932 152380
rect 413836 152328 413888 152380
rect 416228 152328 416280 152380
rect 416596 152328 416648 152380
rect 33600 152260 33652 152312
rect 109684 152260 109736 152312
rect 109776 152260 109828 152312
rect 127900 152260 127952 152312
rect 127992 152260 128044 152312
rect 215852 152260 215904 152312
rect 223856 152260 223908 152312
rect 287796 152260 287848 152312
rect 288348 152260 288400 152312
rect 289912 152260 289964 152312
rect 292212 152260 292264 152312
rect 341708 152260 341760 152312
rect 342444 152260 342496 152312
rect 344284 152260 344336 152312
rect 345204 152260 345256 152312
rect 382280 152260 382332 152312
rect 382372 152260 382424 152312
rect 386696 152260 386748 152312
rect 389180 152260 389232 152312
rect 412640 152260 412692 152312
rect 9496 152192 9548 152244
rect 82820 152192 82872 152244
rect 82912 152192 82964 152244
rect 169760 152192 169812 152244
rect 78864 152124 78916 152176
rect 164516 152124 164568 152176
rect 167000 152124 167052 152176
rect 169944 152124 169996 152176
rect 176108 152192 176160 152244
rect 190184 152192 190236 152244
rect 194508 152192 194560 152244
rect 213276 152192 213328 152244
rect 221740 152192 221792 152244
rect 282920 152192 282972 152244
rect 285772 152192 285824 152244
rect 335912 152192 335964 152244
rect 68928 152056 68980 152108
rect 149152 152056 149204 152108
rect 156880 152056 156932 152108
rect 172520 152056 172572 152108
rect 182456 152124 182508 152176
rect 183468 152124 183520 152176
rect 185032 152056 185084 152108
rect 191656 152124 191708 152176
rect 208400 152124 208452 152176
rect 213644 152124 213696 152176
rect 274272 152124 274324 152176
rect 277952 152124 278004 152176
rect 279608 152124 279660 152176
rect 291384 152124 291436 152176
rect 341064 152192 341116 152244
rect 341156 152192 341208 152244
rect 375380 152192 375432 152244
rect 385500 152192 385552 152244
rect 387340 152192 387392 152244
rect 388352 152192 388404 152244
rect 340144 152124 340196 152176
rect 346400 152124 346452 152176
rect 349804 152124 349856 152176
rect 380256 152124 380308 152176
rect 383752 152124 383804 152176
rect 391940 152124 391992 152176
rect 394608 152192 394660 152244
rect 417332 152192 417384 152244
rect 421748 152328 421800 152380
rect 436284 152328 436336 152380
rect 417608 152260 417660 152312
rect 421472 152260 421524 152312
rect 425152 152260 425204 152312
rect 426532 152192 426584 152244
rect 426716 152260 426768 152312
rect 441252 152328 441304 152380
rect 441712 152328 441764 152380
rect 455420 152328 455472 152380
rect 441528 152260 441580 152312
rect 454776 152260 454828 152312
rect 443184 152192 443236 152244
rect 443644 152192 443696 152244
rect 457352 152192 457404 152244
rect 407212 152124 407264 152176
rect 409328 152124 409380 152176
rect 428372 152124 428424 152176
rect 429292 152124 429344 152176
rect 446404 152124 446456 152176
rect 200488 152056 200540 152108
rect 242808 152056 242860 152108
rect 300860 152056 300912 152108
rect 303988 152056 304040 152108
rect 350724 152056 350776 152108
rect 355324 152056 355376 152108
rect 389916 152056 389968 152108
rect 405648 152056 405700 152108
rect 75092 151988 75144 152040
rect 154212 151988 154264 152040
rect 162492 151988 162544 152040
rect 177396 151988 177448 152040
rect 184664 151988 184716 152040
rect 195336 151988 195388 152040
rect 243360 151988 243412 152040
rect 302608 151988 302660 152040
rect 19800 151920 19852 151972
rect 97908 151920 97960 151972
rect 103796 151920 103848 151972
rect 109868 151920 109920 151972
rect 109960 151920 110012 151972
rect 138296 151920 138348 151972
rect 139308 151920 139360 151972
rect 74816 151852 74868 151904
rect 81348 151852 81400 151904
rect 109040 151852 109092 151904
rect 130476 151852 130528 151904
rect 130660 151852 130712 151904
rect 146576 151852 146628 151904
rect 146668 151852 146720 151904
rect 167092 151852 167144 151904
rect 203064 151920 203116 151972
rect 213092 151920 213144 151972
rect 272432 151920 272484 151972
rect 272524 151920 272576 151972
rect 325700 151988 325752 152040
rect 330484 151988 330536 152040
rect 362316 151988 362368 152040
rect 387892 151988 387944 152040
rect 404636 151988 404688 152040
rect 325884 151920 325936 151972
rect 330576 151920 330628 151972
rect 331772 151920 331824 151972
rect 371884 151920 371936 151972
rect 378784 151920 378836 151972
rect 384120 151920 384172 151972
rect 385868 151920 385920 151972
rect 399484 151920 399536 151972
rect 399576 151920 399628 151972
rect 413008 151988 413060 152040
rect 417424 152056 417476 152108
rect 420920 151988 420972 152040
rect 422576 152056 422628 152108
rect 426716 152056 426768 152108
rect 426808 152056 426860 152108
rect 444472 152056 444524 152108
rect 515772 152056 515824 152108
rect 518900 152056 518952 152108
rect 423312 151988 423364 152040
rect 423588 151988 423640 152040
rect 439320 151988 439372 152040
rect 439412 151988 439464 152040
rect 454224 151988 454276 152040
rect 459560 151988 459612 152040
rect 461768 151988 461820 152040
rect 486516 151988 486568 152040
rect 490012 151988 490064 152040
rect 515956 151988 516008 152040
rect 519452 151988 519504 152040
rect 413744 151920 413796 151972
rect 283012 151852 283064 151904
rect 287152 151852 287204 151904
rect 299940 151852 299992 151904
rect 340144 151852 340196 151904
rect 349436 151852 349488 151904
rect 71412 151784 71464 151836
rect 92480 151784 92532 151836
rect 105820 151784 105872 151836
rect 110328 151784 110380 151836
rect 113916 151784 113968 151836
rect 121000 151784 121052 151836
rect 138020 151784 138072 151836
rect 141424 151784 141476 151836
rect 142252 151784 142304 151836
rect 151820 151784 151872 151836
rect 154304 151784 154356 151836
rect 236460 151784 236512 151836
rect 272616 151784 272668 151836
rect 326344 151784 326396 151836
rect 336004 151784 336056 151836
rect 341156 151784 341208 151836
rect 343824 151784 343876 151836
rect 349804 151784 349856 151836
rect 362960 151784 363012 151836
rect 364340 151784 364392 151836
rect 386328 151852 386380 151904
rect 394700 151852 394752 151904
rect 396264 151852 396316 151904
rect 402980 151852 403032 151904
rect 404268 151852 404320 151904
rect 418160 151852 418212 151904
rect 419632 151920 419684 151972
rect 436744 151920 436796 151972
rect 421380 151852 421432 151904
rect 421472 151852 421524 151904
rect 431592 151852 431644 151904
rect 436284 151852 436336 151904
rect 440608 151852 440660 151904
rect 385408 151784 385460 151836
rect 403900 151784 403952 151836
rect 415676 151784 415728 151836
rect 419724 151784 419776 151836
rect 434168 151784 434220 151836
rect 436192 151784 436244 151836
rect 451556 151920 451608 151972
rect 469220 151920 469272 151972
rect 472072 151920 472124 151972
rect 487344 151920 487396 151972
rect 490656 151920 490708 151972
rect 507768 151920 507820 151972
rect 509240 151920 509292 151972
rect 517428 151920 517480 151972
rect 521568 151920 521620 151972
rect 442908 151852 442960 151904
rect 450912 151852 450964 151904
rect 468024 151852 468076 151904
rect 470784 151852 470836 151904
rect 489092 151852 489144 151904
rect 491944 151852 491996 151904
rect 442724 151784 442776 151836
rect 456064 151784 456116 151836
rect 467840 151784 467892 151836
rect 471428 151784 471480 151836
rect 488448 151784 488500 151836
rect 491300 151784 491352 151836
rect 509056 151784 509108 151836
rect 510896 151784 510948 151836
rect 517060 151784 517112 151836
rect 520280 151784 520332 151836
rect 81716 151716 81768 151768
rect 112904 151716 112956 151768
rect 98920 151648 98972 151700
rect 116032 151648 116084 151700
rect 95516 151580 95568 151632
rect 115296 151580 115348 151632
rect 92020 151512 92072 151564
rect 113088 151512 113140 151564
rect 26700 151444 26752 151496
rect 116952 151444 117004 151496
rect 16396 151376 16448 151428
rect 116768 151376 116820 151428
rect 12992 151308 13044 151360
rect 116676 151308 116728 151360
rect 68008 151240 68060 151292
rect 112720 151240 112772 151292
rect 64512 151172 64564 151224
rect 112628 151172 112680 151224
rect 61108 151104 61160 151156
rect 112536 151104 112588 151156
rect 57704 151036 57756 151088
rect 110972 151036 111024 151088
rect 54208 150968 54260 151020
rect 112444 150968 112496 151020
rect 50804 150900 50856 150952
rect 111708 150900 111760 150952
rect 47308 150832 47360 150884
rect 111616 150832 111668 150884
rect 43904 150764 43956 150816
rect 111524 150764 111576 150816
rect 40500 150696 40552 150748
rect 111432 150696 111484 150748
rect 37004 150628 37056 150680
rect 111248 150628 111300 150680
rect 88616 150560 88668 150612
rect 112996 150560 113048 150612
rect 85212 150492 85264 150544
rect 115204 150492 115256 150544
rect 285680 150492 285732 150544
rect 286508 150492 286560 150544
rect 342260 150492 342312 150544
rect 342996 150492 343048 150544
rect 102324 150424 102376 150476
rect 116124 150424 116176 150476
rect 78312 150288 78364 150340
rect 112812 150288 112864 150340
rect 109592 150220 109644 150272
rect 117136 150220 117188 150272
rect 97908 150152 97960 150204
rect 116860 150152 116912 150204
rect 81348 150084 81400 150136
rect 92480 150084 92532 150136
rect 117228 150084 117280 150136
rect 116492 150016 116544 150068
rect 111156 148316 111208 148368
rect 117044 148316 117096 148368
rect 113088 140700 113140 140752
rect 116124 140700 116176 140752
rect 112996 137912 113048 137964
rect 116124 137912 116176 137964
rect 112904 133832 112956 133884
rect 116032 133832 116084 133884
rect 114192 132608 114244 132660
rect 115204 132608 115256 132660
rect 112812 132404 112864 132456
rect 116124 132404 116176 132456
rect 112720 126896 112772 126948
rect 116124 126896 116176 126948
rect 112628 124108 112680 124160
rect 116124 124108 116176 124160
rect 112536 122748 112588 122800
rect 115940 122748 115992 122800
rect 111708 121388 111760 121440
rect 116124 121388 116176 121440
rect 112444 118600 112496 118652
rect 116124 118600 116176 118652
rect 111616 117240 111668 117292
rect 116124 117240 116176 117292
rect 111524 114452 111576 114504
rect 116124 114452 116176 114504
rect 111432 113092 111484 113144
rect 115940 113092 115992 113144
rect 111340 111732 111392 111784
rect 116124 111732 116176 111784
rect 111156 108944 111208 108996
rect 116124 108944 116176 108996
rect 111248 92420 111300 92472
rect 116124 92420 116176 92472
rect 111064 89632 111116 89684
rect 116124 89632 116176 89684
rect 113824 88272 113876 88324
rect 116032 88272 116084 88324
rect 113916 83920 113968 83972
rect 116584 83920 116636 83972
rect 114008 82764 114060 82816
rect 116216 82764 116268 82816
rect 114100 79976 114152 80028
rect 115940 79976 115992 80028
rect 114192 78616 114244 78668
rect 116124 78616 116176 78668
rect 114192 71748 114244 71800
rect 116584 71748 116636 71800
rect 114100 69028 114152 69080
rect 116308 69028 116360 69080
rect 114008 67600 114060 67652
rect 116124 67600 116176 67652
rect 113916 66240 113968 66292
rect 116584 66240 116636 66292
rect 113364 64676 113416 64728
rect 116584 64676 116636 64728
rect 113824 63520 113876 63572
rect 116216 63520 116268 63572
rect 112444 62092 112496 62144
rect 116124 62092 116176 62144
rect 112536 42780 112588 42832
rect 116124 42780 116176 42832
rect 116400 7624 116452 7676
rect 116308 7420 116360 7472
rect 111708 2796 111760 2848
rect 143632 2456 143684 2508
rect 425796 2456 425848 2508
rect 443644 2456 443696 2508
rect 42064 1844 42116 1896
rect 44732 1844 44784 1896
rect 58992 1844 59044 1896
rect 66996 1844 67048 1896
rect 90364 1844 90416 1896
rect 92572 1844 92624 1896
rect 95332 1844 95384 1896
rect 99932 1844 99984 1896
rect 100024 1844 100076 1896
rect 102692 1844 102744 1896
rect 59176 1776 59228 1828
rect 63040 1776 63092 1828
rect 89352 1776 89404 1828
rect 105912 1844 105964 1896
rect 109132 1844 109184 1896
rect 109684 1844 109736 1896
rect 109776 1844 109828 1896
rect 109868 1844 109920 1896
rect 59360 1708 59412 1760
rect 76564 1708 76616 1760
rect 86040 1708 86092 1760
rect 109316 1776 109368 1828
rect 112444 1776 112496 1828
rect 82636 1640 82688 1692
rect 103980 1640 104032 1692
rect 109960 1708 110012 1760
rect 110052 1708 110104 1760
rect 116584 1708 116636 1760
rect 69296 1572 69348 1624
rect 101772 1572 101824 1624
rect 79324 1504 79376 1556
rect 105912 1572 105964 1624
rect 106004 1572 106056 1624
rect 109040 1572 109092 1624
rect 109224 1640 109276 1692
rect 110604 1640 110656 1692
rect 110144 1572 110196 1624
rect 103980 1504 104032 1556
rect 110236 1504 110288 1556
rect 46020 1436 46072 1488
rect 64604 1436 64656 1488
rect 72700 1436 72752 1488
rect 109592 1436 109644 1488
rect 193588 1436 193640 1488
rect 32680 1368 32732 1420
rect 109132 1368 109184 1420
rect 109224 1368 109276 1420
rect 110052 1368 110104 1420
rect 2688 1300 2740 1352
rect 35992 1232 36044 1284
rect 109408 1300 109460 1352
rect 116400 1368 116452 1420
rect 294788 1368 294840 1420
rect 343640 1368 343692 1420
rect 491300 1368 491352 1420
rect 493600 1368 493652 1420
rect 39304 1164 39356 1216
rect 109040 1164 109092 1216
rect 116308 1232 116360 1284
rect 116492 1164 116544 1216
rect 49332 1096 49384 1148
rect 117044 1096 117096 1148
rect 52644 1028 52696 1080
rect 65984 960 66036 1012
rect 101404 960 101456 1012
rect 76012 892 76064 944
rect 116860 960 116912 1012
rect 112536 892 112588 944
rect 89720 824 89772 876
rect 95976 824 96028 876
rect 100852 824 100904 876
rect 101404 824 101456 876
rect 116676 824 116728 876
rect 102784 756 102836 808
rect 109040 756 109092 808
rect 117228 756 117280 808
<< metal2 >>
rect 386 163200 442 164400
rect 1214 163200 1270 164400
rect 2042 163200 2098 164400
rect 2870 163200 2926 164400
rect 3698 163200 3754 164400
rect 3804 163254 4016 163282
rect 400 158030 428 163200
rect 388 158024 440 158030
rect 388 157966 440 157972
rect 1228 153882 1256 163200
rect 2056 156670 2084 163200
rect 2044 156664 2096 156670
rect 2044 156606 2096 156612
rect 1216 153876 1268 153882
rect 1216 153818 1268 153824
rect 2884 152522 2912 163200
rect 3712 163146 3740 163200
rect 3804 163146 3832 163254
rect 3712 163118 3832 163146
rect 3988 153785 4016 163254
rect 4526 163200 4582 164400
rect 5354 163200 5410 164400
rect 6274 163200 6330 164400
rect 7102 163200 7158 164400
rect 7930 163200 7986 164400
rect 8758 163200 8814 164400
rect 9586 163200 9642 164400
rect 10414 163200 10470 164400
rect 11242 163200 11298 164400
rect 12162 163200 12218 164400
rect 12990 163200 13046 164400
rect 13818 163200 13874 164400
rect 14646 163200 14702 164400
rect 15474 163200 15530 164400
rect 16302 163200 16358 164400
rect 17130 163200 17186 164400
rect 18050 163200 18106 164400
rect 18878 163200 18934 164400
rect 19706 163200 19762 164400
rect 20534 163200 20590 164400
rect 21362 163200 21418 164400
rect 22190 163200 22246 164400
rect 23018 163200 23074 164400
rect 23938 163200 23994 164400
rect 24766 163200 24822 164400
rect 25594 163200 25650 164400
rect 26422 163200 26478 164400
rect 27250 163200 27306 164400
rect 28078 163200 28134 164400
rect 28906 163200 28962 164400
rect 29826 163200 29882 164400
rect 30654 163200 30710 164400
rect 31482 163200 31538 164400
rect 32310 163200 32366 164400
rect 33138 163200 33194 164400
rect 33966 163200 34022 164400
rect 34794 163200 34850 164400
rect 35714 163200 35770 164400
rect 36542 163200 36598 164400
rect 37370 163200 37426 164400
rect 38198 163200 38254 164400
rect 38304 163254 38516 163282
rect 4540 155446 4568 163200
rect 4528 155440 4580 155446
rect 4528 155382 4580 155388
rect 5368 155242 5396 163200
rect 6288 159390 6316 163200
rect 6276 159384 6328 159390
rect 6276 159326 6328 159332
rect 5356 155236 5408 155242
rect 5356 155178 5408 155184
rect 7116 153950 7144 163200
rect 7944 155378 7972 163200
rect 7932 155372 7984 155378
rect 7932 155314 7984 155320
rect 8772 155310 8800 163200
rect 8760 155304 8812 155310
rect 8760 155246 8812 155252
rect 7104 153944 7156 153950
rect 7104 153886 7156 153892
rect 3974 153776 4030 153785
rect 3974 153711 4030 153720
rect 2872 152516 2924 152522
rect 2872 152458 2924 152464
rect 9600 152425 9628 163200
rect 10428 154018 10456 163200
rect 11256 156806 11284 163200
rect 11244 156800 11296 156806
rect 11244 156742 11296 156748
rect 12176 155786 12204 163200
rect 12164 155780 12216 155786
rect 12164 155722 12216 155728
rect 10416 154012 10468 154018
rect 10416 153954 10468 153960
rect 13004 152561 13032 163200
rect 13832 154086 13860 163200
rect 14660 156738 14688 163200
rect 14648 156732 14700 156738
rect 14648 156674 14700 156680
rect 15488 154970 15516 163200
rect 16316 159361 16344 163200
rect 16302 159352 16358 159361
rect 16302 159287 16358 159296
rect 15476 154964 15528 154970
rect 15476 154906 15528 154912
rect 13820 154080 13872 154086
rect 17144 154057 17172 163200
rect 18064 156942 18092 163200
rect 18892 159730 18920 163200
rect 18880 159724 18932 159730
rect 18880 159666 18932 159672
rect 18052 156936 18104 156942
rect 18052 156878 18104 156884
rect 13820 154022 13872 154028
rect 17130 154048 17186 154057
rect 17130 153983 17186 153992
rect 19720 152590 19748 163200
rect 20548 153921 20576 163200
rect 21376 156874 21404 163200
rect 21364 156868 21416 156874
rect 21364 156810 21416 156816
rect 20534 153912 20590 153921
rect 20534 153847 20590 153856
rect 22204 152658 22232 163200
rect 23032 159497 23060 163200
rect 23018 159488 23074 159497
rect 23018 159423 23074 159432
rect 23952 154222 23980 163200
rect 24780 157010 24808 163200
rect 25608 160002 25636 163200
rect 25596 159996 25648 160002
rect 25596 159938 25648 159944
rect 24768 157004 24820 157010
rect 24768 156946 24820 156952
rect 23940 154216 23992 154222
rect 23940 154158 23992 154164
rect 26436 152794 26464 163200
rect 27264 154154 27292 163200
rect 28092 156641 28120 163200
rect 28078 156632 28134 156641
rect 28078 156567 28134 156576
rect 27252 154148 27304 154154
rect 27252 154090 27304 154096
rect 26424 152788 26476 152794
rect 26424 152730 26476 152736
rect 28920 152726 28948 163200
rect 29840 159633 29868 163200
rect 29826 159624 29882 159633
rect 29826 159559 29882 159568
rect 30668 154193 30696 163200
rect 31496 156777 31524 163200
rect 32324 159458 32352 163200
rect 32312 159452 32364 159458
rect 32312 159394 32364 159400
rect 31482 156768 31538 156777
rect 31482 156703 31538 156712
rect 30654 154184 30710 154193
rect 30654 154119 30710 154128
rect 30196 153128 30248 153134
rect 30196 153070 30248 153076
rect 28908 152720 28960 152726
rect 28908 152662 28960 152668
rect 22192 152652 22244 152658
rect 22192 152594 22244 152600
rect 19708 152584 19760 152590
rect 12990 152552 13046 152561
rect 19708 152526 19760 152532
rect 12990 152487 13046 152496
rect 23296 152448 23348 152454
rect 9586 152416 9642 152425
rect 23296 152390 23348 152396
rect 9586 152351 9642 152360
rect 9496 152244 9548 152250
rect 9496 152186 9548 152192
rect 6090 150648 6146 150657
rect 6090 150583 6146 150592
rect 2686 150512 2742 150521
rect 2686 150447 2742 150456
rect 2700 149940 2728 150447
rect 6104 149940 6132 150583
rect 9508 149940 9536 152186
rect 19800 151972 19852 151978
rect 19800 151914 19852 151920
rect 16396 151428 16448 151434
rect 16396 151370 16448 151376
rect 12992 151360 13044 151366
rect 12992 151302 13044 151308
rect 13004 149940 13032 151302
rect 16408 149940 16436 151370
rect 19812 149940 19840 151914
rect 23308 149940 23336 152390
rect 26700 151496 26752 151502
rect 26700 151438 26752 151444
rect 26712 149940 26740 151438
rect 30208 149940 30236 153070
rect 33152 152862 33180 163200
rect 33980 158001 34008 163200
rect 33966 157992 34022 158001
rect 33966 157927 34022 157936
rect 34808 153270 34836 163200
rect 35728 157078 35756 163200
rect 36556 159526 36584 163200
rect 36544 159520 36596 159526
rect 36544 159462 36596 159468
rect 37384 158098 37412 163200
rect 38212 163146 38240 163200
rect 38304 163146 38332 163254
rect 38212 163118 38332 163146
rect 37372 158092 37424 158098
rect 37372 158034 37424 158040
rect 35716 157072 35768 157078
rect 35716 157014 35768 157020
rect 38488 154290 38516 163254
rect 39026 163200 39082 164400
rect 39854 163200 39910 164400
rect 40682 163200 40738 164400
rect 41602 163200 41658 164400
rect 42430 163200 42486 164400
rect 43258 163200 43314 164400
rect 44086 163200 44142 164400
rect 44914 163200 44970 164400
rect 45742 163200 45798 164400
rect 46570 163200 46626 164400
rect 47490 163200 47546 164400
rect 48318 163200 48374 164400
rect 49146 163200 49202 164400
rect 49974 163200 50030 164400
rect 50802 163200 50858 164400
rect 51630 163200 51686 164400
rect 52458 163200 52514 164400
rect 53378 163200 53434 164400
rect 54206 163200 54262 164400
rect 55034 163200 55090 164400
rect 55862 163200 55918 164400
rect 56690 163200 56746 164400
rect 57518 163200 57574 164400
rect 58346 163200 58402 164400
rect 59266 163200 59322 164400
rect 60094 163200 60150 164400
rect 60922 163200 60978 164400
rect 61750 163200 61806 164400
rect 62578 163200 62634 164400
rect 63406 163200 63462 164400
rect 64234 163200 64290 164400
rect 65154 163200 65210 164400
rect 65982 163200 66038 164400
rect 66810 163200 66866 164400
rect 67638 163200 67694 164400
rect 68466 163200 68522 164400
rect 69294 163200 69350 164400
rect 70122 163200 70178 164400
rect 71042 163200 71098 164400
rect 71870 163200 71926 164400
rect 72698 163200 72754 164400
rect 73526 163200 73582 164400
rect 74354 163200 74410 164400
rect 75182 163200 75238 164400
rect 76010 163200 76066 164400
rect 76930 163200 76986 164400
rect 77758 163200 77814 164400
rect 78586 163200 78642 164400
rect 79414 163200 79470 164400
rect 80242 163200 80298 164400
rect 81070 163200 81126 164400
rect 81898 163200 81954 164400
rect 82818 163200 82874 164400
rect 83646 163200 83702 164400
rect 84474 163200 84530 164400
rect 85302 163200 85358 164400
rect 86130 163200 86186 164400
rect 86958 163200 87014 164400
rect 87786 163200 87842 164400
rect 88706 163200 88762 164400
rect 89534 163200 89590 164400
rect 90362 163200 90418 164400
rect 91190 163200 91246 164400
rect 92018 163200 92074 164400
rect 92846 163200 92902 164400
rect 93674 163200 93730 164400
rect 94594 163200 94650 164400
rect 95422 163200 95478 164400
rect 96250 163200 96306 164400
rect 97078 163200 97134 164400
rect 97906 163200 97962 164400
rect 98734 163200 98790 164400
rect 99562 163200 99618 164400
rect 100482 163200 100538 164400
rect 101310 163200 101366 164400
rect 102138 163200 102194 164400
rect 102966 163200 103022 164400
rect 103794 163200 103850 164400
rect 104622 163200 104678 164400
rect 105450 163200 105506 164400
rect 106370 163200 106426 164400
rect 107198 163200 107254 164400
rect 108026 163200 108082 164400
rect 108854 163200 108910 164400
rect 109682 163200 109738 164400
rect 110510 163200 110566 164400
rect 111338 163200 111394 164400
rect 112258 163200 112314 164400
rect 113086 163200 113142 164400
rect 113914 163200 113970 164400
rect 114742 163200 114798 164400
rect 115570 163200 115626 164400
rect 116398 163200 116454 164400
rect 117226 163200 117282 164400
rect 118146 163200 118202 164400
rect 118974 163200 119030 164400
rect 119802 163200 119858 164400
rect 120630 163200 120686 164400
rect 121458 163200 121514 164400
rect 122286 163200 122342 164400
rect 123114 163200 123170 164400
rect 124034 163200 124090 164400
rect 124862 163200 124918 164400
rect 125690 163200 125746 164400
rect 126518 163200 126574 164400
rect 127346 163200 127402 164400
rect 128174 163200 128230 164400
rect 129002 163200 129058 164400
rect 129922 163200 129978 164400
rect 130750 163200 130806 164400
rect 131578 163200 131634 164400
rect 132406 163200 132462 164400
rect 133234 163200 133290 164400
rect 134062 163200 134118 164400
rect 134890 163200 134946 164400
rect 135810 163200 135866 164400
rect 136638 163200 136694 164400
rect 136744 163254 137416 163282
rect 39040 157214 39068 163200
rect 39028 157208 39080 157214
rect 39028 157150 39080 157156
rect 39868 155582 39896 163200
rect 40696 158137 40724 163200
rect 40682 158128 40738 158137
rect 40682 158063 40738 158072
rect 39856 155576 39908 155582
rect 39856 155518 39908 155524
rect 41616 154426 41644 163200
rect 42444 157146 42472 163200
rect 43272 159594 43300 163200
rect 43260 159588 43312 159594
rect 43260 159530 43312 159536
rect 44100 158273 44128 163200
rect 44086 158264 44142 158273
rect 44086 158199 44142 158208
rect 42432 157140 42484 157146
rect 42432 157082 42484 157088
rect 44928 154494 44956 163200
rect 45756 157282 45784 163200
rect 45744 157276 45796 157282
rect 45744 157218 45796 157224
rect 46584 155650 46612 163200
rect 47504 158166 47532 163200
rect 47492 158160 47544 158166
rect 47492 158102 47544 158108
rect 46572 155644 46624 155650
rect 46572 155586 46624 155592
rect 44916 154488 44968 154494
rect 44916 154430 44968 154436
rect 41604 154420 41656 154426
rect 41604 154362 41656 154368
rect 38476 154284 38528 154290
rect 38476 154226 38528 154232
rect 48332 153814 48360 163200
rect 49160 157350 49188 163200
rect 49988 159662 50016 163200
rect 49976 159656 50028 159662
rect 49976 159598 50028 159604
rect 50816 158234 50844 163200
rect 50804 158228 50856 158234
rect 50804 158170 50856 158176
rect 49148 157344 49200 157350
rect 49148 157286 49200 157292
rect 51644 154562 51672 163200
rect 52472 156602 52500 163200
rect 52460 156596 52512 156602
rect 52460 156538 52512 156544
rect 53392 155854 53420 163200
rect 54220 158302 54248 163200
rect 54208 158296 54260 158302
rect 54208 158238 54260 158244
rect 53380 155848 53432 155854
rect 53380 155790 53432 155796
rect 51632 154556 51684 154562
rect 51632 154498 51684 154504
rect 55048 154329 55076 163200
rect 55876 156913 55904 163200
rect 56704 159798 56732 163200
rect 56692 159792 56744 159798
rect 56692 159734 56744 159740
rect 57532 158409 57560 163200
rect 57518 158400 57574 158409
rect 57518 158335 57574 158344
rect 55862 156904 55918 156913
rect 55862 156839 55918 156848
rect 55034 154320 55090 154329
rect 55034 154255 55090 154264
rect 48320 153808 48372 153814
rect 48320 153750 48372 153756
rect 58360 153678 58388 163200
rect 59280 156534 59308 163200
rect 59268 156528 59320 156534
rect 59268 156470 59320 156476
rect 60108 155718 60136 163200
rect 60936 158438 60964 163200
rect 60924 158432 60976 158438
rect 60924 158374 60976 158380
rect 60096 155712 60148 155718
rect 60096 155654 60148 155660
rect 61764 153746 61792 163200
rect 62592 155553 62620 163200
rect 63420 160070 63448 163200
rect 63408 160064 63460 160070
rect 63408 160006 63460 160012
rect 64248 158370 64276 163200
rect 64236 158364 64288 158370
rect 64236 158306 64288 158312
rect 62578 155544 62634 155553
rect 65168 155514 65196 163200
rect 62578 155479 62634 155488
rect 65156 155508 65208 155514
rect 65156 155450 65208 155456
rect 65996 155281 66024 163200
rect 66824 155854 66852 163200
rect 67652 158506 67680 163200
rect 67640 158500 67692 158506
rect 67640 158442 67692 158448
rect 66720 155848 66772 155854
rect 66720 155790 66772 155796
rect 66812 155848 66864 155854
rect 66812 155790 66864 155796
rect 65982 155272 66038 155281
rect 65982 155207 66038 155216
rect 61752 153740 61804 153746
rect 61752 153682 61804 153688
rect 58348 153672 58400 153678
rect 58348 153614 58400 153620
rect 34796 153264 34848 153270
rect 34796 153206 34848 153212
rect 66732 153202 66760 155790
rect 68480 155417 68508 163200
rect 69308 156466 69336 163200
rect 70136 159866 70164 163200
rect 70124 159860 70176 159866
rect 70124 159802 70176 159808
rect 71056 158574 71084 163200
rect 71044 158568 71096 158574
rect 71044 158510 71096 158516
rect 69296 156460 69348 156466
rect 69296 156402 69348 156408
rect 71884 155582 71912 163200
rect 72712 157049 72740 163200
rect 73540 159322 73568 163200
rect 73528 159316 73580 159322
rect 73528 159258 73580 159264
rect 74368 158642 74396 163200
rect 74356 158636 74408 158642
rect 74356 158578 74408 158584
rect 72698 157040 72754 157049
rect 72698 156975 72754 156984
rect 75196 155650 75224 163200
rect 76024 155825 76052 163200
rect 76944 159934 76972 163200
rect 76932 159928 76984 159934
rect 76932 159870 76984 159876
rect 77772 157962 77800 163200
rect 77760 157956 77812 157962
rect 77760 157898 77812 157904
rect 76010 155816 76066 155825
rect 76010 155751 76066 155760
rect 78600 155689 78628 163200
rect 78864 155712 78916 155718
rect 78586 155680 78642 155689
rect 75092 155644 75144 155650
rect 75092 155586 75144 155592
rect 75184 155644 75236 155650
rect 78864 155654 78916 155660
rect 78586 155615 78642 155624
rect 75184 155586 75236 155592
rect 68928 155576 68980 155582
rect 68928 155518 68980 155524
rect 71872 155576 71924 155582
rect 71872 155518 71924 155524
rect 68466 155408 68522 155417
rect 68466 155343 68522 155352
rect 66720 153196 66772 153202
rect 66720 153138 66772 153144
rect 33140 152856 33192 152862
rect 33140 152798 33192 152804
rect 33600 152312 33652 152318
rect 33600 152254 33652 152260
rect 33612 149940 33640 152254
rect 68940 152114 68968 155518
rect 68928 152108 68980 152114
rect 68928 152050 68980 152056
rect 75104 152046 75132 155586
rect 78876 152182 78904 155654
rect 79428 153610 79456 163200
rect 80060 159316 80112 159322
rect 80060 159258 80112 159264
rect 79416 153604 79468 153610
rect 79416 153546 79468 153552
rect 80072 153066 80100 159258
rect 80256 159254 80284 163200
rect 80244 159248 80296 159254
rect 80244 159190 80296 159196
rect 81084 158710 81112 163200
rect 81072 158704 81124 158710
rect 81072 158646 81124 158652
rect 81912 155718 81940 163200
rect 82832 156398 82860 163200
rect 83660 159322 83688 163200
rect 83648 159316 83700 159322
rect 83648 159258 83700 159264
rect 84488 157894 84516 163200
rect 84476 157888 84528 157894
rect 84476 157830 84528 157836
rect 82820 156392 82872 156398
rect 82820 156334 82872 156340
rect 85316 155961 85344 163200
rect 85302 155952 85358 155961
rect 85302 155887 85358 155896
rect 82912 155848 82964 155854
rect 82912 155790 82964 155796
rect 81900 155712 81952 155718
rect 81900 155654 81952 155660
rect 80060 153060 80112 153066
rect 80060 153002 80112 153008
rect 82924 152250 82952 155790
rect 86144 154465 86172 163200
rect 86972 159186 87000 163200
rect 86960 159180 87012 159186
rect 86960 159122 87012 159128
rect 87800 157826 87828 163200
rect 87788 157820 87840 157826
rect 87788 157762 87840 157768
rect 88720 155854 88748 163200
rect 89548 155922 89576 163200
rect 90376 158778 90404 163200
rect 91100 159248 91152 159254
rect 91100 159190 91152 159196
rect 90364 158772 90416 158778
rect 90364 158714 90416 158720
rect 89536 155916 89588 155922
rect 89536 155858 89588 155864
rect 88708 155848 88760 155854
rect 88708 155790 88760 155796
rect 86130 154456 86186 154465
rect 86130 154391 86186 154400
rect 91112 152386 91140 159190
rect 91204 157758 91232 163200
rect 91192 157752 91244 157758
rect 91192 157694 91244 157700
rect 92032 155174 92060 163200
rect 92860 158778 92888 163200
rect 93688 159118 93716 163200
rect 93676 159112 93728 159118
rect 93676 159054 93728 159060
rect 92480 158772 92532 158778
rect 92480 158714 92532 158720
rect 92848 158772 92900 158778
rect 92848 158714 92900 158720
rect 92020 155168 92072 155174
rect 92020 155110 92072 155116
rect 92492 152930 92520 158714
rect 94608 157690 94636 163200
rect 94596 157684 94648 157690
rect 94596 157626 94648 157632
rect 95436 155106 95464 163200
rect 96264 158982 96292 163200
rect 96252 158976 96304 158982
rect 96252 158918 96304 158924
rect 95424 155100 95476 155106
rect 95424 155042 95476 155048
rect 97092 152998 97120 163200
rect 97920 157622 97948 163200
rect 97908 157616 97960 157622
rect 97908 157558 97960 157564
rect 98748 155038 98776 163200
rect 99576 156262 99604 163200
rect 100496 159254 100524 163200
rect 100484 159248 100536 159254
rect 100484 159190 100536 159196
rect 101324 156330 101352 163200
rect 101312 156324 101364 156330
rect 101312 156266 101364 156272
rect 99564 156256 99616 156262
rect 99564 156198 99616 156204
rect 98736 155032 98788 155038
rect 98736 154974 98788 154980
rect 102152 153542 102180 163200
rect 102980 158846 103008 163200
rect 102968 158840 103020 158846
rect 102968 158782 103020 158788
rect 102140 153536 102192 153542
rect 102140 153478 102192 153484
rect 97080 152992 97132 152998
rect 97080 152934 97132 152940
rect 92480 152924 92532 152930
rect 92480 152866 92532 152872
rect 91100 152380 91152 152386
rect 91100 152322 91152 152328
rect 82820 152244 82872 152250
rect 82820 152186 82872 152192
rect 82912 152244 82964 152250
rect 82912 152186 82964 152192
rect 78864 152176 78916 152182
rect 78864 152118 78916 152124
rect 75092 152040 75144 152046
rect 75092 151982 75144 151988
rect 74816 151904 74868 151910
rect 74816 151846 74868 151852
rect 81348 151904 81400 151910
rect 81348 151846 81400 151852
rect 71412 151836 71464 151842
rect 71412 151778 71464 151784
rect 68008 151292 68060 151298
rect 68008 151234 68060 151240
rect 64512 151224 64564 151230
rect 64512 151166 64564 151172
rect 61108 151156 61160 151162
rect 61108 151098 61160 151104
rect 57704 151088 57756 151094
rect 57704 151030 57756 151036
rect 54208 151020 54260 151026
rect 54208 150962 54260 150968
rect 50804 150952 50856 150958
rect 50804 150894 50856 150900
rect 47308 150884 47360 150890
rect 47308 150826 47360 150832
rect 43904 150816 43956 150822
rect 43904 150758 43956 150764
rect 40500 150748 40552 150754
rect 40500 150690 40552 150696
rect 37004 150680 37056 150686
rect 37004 150622 37056 150628
rect 37016 149940 37044 150622
rect 40512 149940 40540 150690
rect 43916 149940 43944 150758
rect 47320 149940 47348 150826
rect 50816 149940 50844 150894
rect 54220 149940 54248 150962
rect 57716 149940 57744 151030
rect 61120 149940 61148 151098
rect 64524 149940 64552 151166
rect 68020 149940 68048 151234
rect 71424 149940 71452 151778
rect 74828 149940 74856 151846
rect 78312 150340 78364 150346
rect 78312 150282 78364 150288
rect 78324 149940 78352 150282
rect 81360 150142 81388 151846
rect 81716 151768 81768 151774
rect 81716 151710 81768 151716
rect 81348 150136 81400 150142
rect 81348 150078 81400 150084
rect 81728 149940 81756 151710
rect 82832 149705 82860 152186
rect 103808 151978 103836 163200
rect 104636 158545 104664 163200
rect 104622 158536 104678 158545
rect 104622 158471 104678 158480
rect 105464 153474 105492 163200
rect 106384 154902 106412 163200
rect 107212 159050 107240 163200
rect 107200 159044 107252 159050
rect 107200 158986 107252 158992
rect 108040 156194 108068 163200
rect 108028 156188 108080 156194
rect 108028 156130 108080 156136
rect 106372 154896 106424 154902
rect 106372 154838 106424 154844
rect 105452 153468 105504 153474
rect 105452 153410 105504 153416
rect 108868 153406 108896 163200
rect 109132 159724 109184 159730
rect 109132 159666 109184 159672
rect 109040 154964 109092 154970
rect 109040 154906 109092 154912
rect 108856 153400 108908 153406
rect 108856 153342 108908 153348
rect 97908 151972 97960 151978
rect 97908 151914 97960 151920
rect 103796 151972 103848 151978
rect 103796 151914 103848 151920
rect 92480 151836 92532 151842
rect 92480 151778 92532 151784
rect 92020 151564 92072 151570
rect 92020 151506 92072 151512
rect 88616 150612 88668 150618
rect 88616 150554 88668 150560
rect 85212 150544 85264 150550
rect 85212 150486 85264 150492
rect 85224 149940 85252 150486
rect 88628 149940 88656 150554
rect 92032 149940 92060 151506
rect 92492 150142 92520 151778
rect 95516 151632 95568 151638
rect 95516 151574 95568 151580
rect 92480 150136 92532 150142
rect 92480 150078 92532 150084
rect 95528 149940 95556 151574
rect 97920 150210 97948 151914
rect 109052 151910 109080 154906
rect 109144 154834 109172 159666
rect 109696 158778 109724 163200
rect 109960 159996 110012 160002
rect 109960 159938 110012 159944
rect 109684 158772 109736 158778
rect 109684 158714 109736 158720
rect 109776 155780 109828 155786
rect 109776 155722 109828 155728
rect 109132 154828 109184 154834
rect 109132 154770 109184 154776
rect 109592 153128 109644 153134
rect 109592 153070 109644 153076
rect 109040 151904 109092 151910
rect 109040 151846 109092 151852
rect 105820 151836 105872 151842
rect 105740 151786 105820 151814
rect 98920 151700 98972 151706
rect 98920 151642 98972 151648
rect 97908 150204 97960 150210
rect 97908 150146 97960 150152
rect 98932 149940 98960 151642
rect 102324 150476 102376 150482
rect 102324 150418 102376 150424
rect 102336 149940 102364 150418
rect 105740 149954 105768 151786
rect 105820 151778 105872 151784
rect 109604 150278 109632 153070
rect 109788 152318 109816 155722
rect 109868 153128 109920 153134
rect 109868 153070 109920 153076
rect 109684 152312 109736 152318
rect 109684 152254 109736 152260
rect 109776 152312 109828 152318
rect 109776 152254 109828 152260
rect 109592 150272 109644 150278
rect 109592 150214 109644 150220
rect 105740 149926 105846 149954
rect 82818 149696 82874 149705
rect 82818 149631 82874 149640
rect 109250 149382 109632 149410
rect 109604 148073 109632 149382
rect 109590 148064 109646 148073
rect 109590 147999 109646 148008
rect 109696 132494 109724 152254
rect 109880 151978 109908 153070
rect 109972 151978 110000 159938
rect 110524 154970 110552 163200
rect 111352 157554 111380 163200
rect 111340 157548 111392 157554
rect 111340 157490 111392 157496
rect 112272 155786 112300 163200
rect 113100 159730 113128 163200
rect 113088 159724 113140 159730
rect 113088 159666 113140 159672
rect 113824 158840 113876 158846
rect 113824 158782 113876 158788
rect 112260 155780 112312 155786
rect 112260 155722 112312 155728
rect 110512 154964 110564 154970
rect 110512 154906 110564 154912
rect 113836 154358 113864 158782
rect 113824 154352 113876 154358
rect 113824 154294 113876 154300
rect 110972 152448 111024 152454
rect 110972 152390 111024 152396
rect 109868 151972 109920 151978
rect 109868 151914 109920 151920
rect 109960 151972 110012 151978
rect 109960 151914 110012 151920
rect 110328 151836 110380 151842
rect 110984 151814 111012 152390
rect 113928 151842 113956 163200
rect 114756 157486 114784 163200
rect 114744 157480 114796 157486
rect 114744 157422 114796 157428
rect 115584 157185 115612 163200
rect 115570 157176 115626 157185
rect 115570 157111 115626 157120
rect 116412 153338 116440 163200
rect 117240 160002 117268 163200
rect 117228 159996 117280 160002
rect 117228 159938 117280 159944
rect 118160 156126 118188 163200
rect 118988 158778 119016 163200
rect 119816 158778 119844 163200
rect 118976 158772 119028 158778
rect 118976 158714 119028 158720
rect 119620 158772 119672 158778
rect 119620 158714 119672 158720
rect 119804 158772 119856 158778
rect 119804 158714 119856 158720
rect 118884 158024 118936 158030
rect 118884 157966 118936 157972
rect 118148 156120 118200 156126
rect 118148 156062 118200 156068
rect 116400 153332 116452 153338
rect 116400 153274 116452 153280
rect 113916 151836 113968 151842
rect 110984 151786 111196 151814
rect 110328 151778 110380 151784
rect 110340 146441 110368 151778
rect 110972 151088 111024 151094
rect 110972 151030 111024 151036
rect 110984 147393 111012 151030
rect 111062 150512 111118 150521
rect 111062 150447 111118 150456
rect 110970 147384 111026 147393
rect 110970 147319 111026 147328
rect 110326 146432 110382 146441
rect 110326 146367 110382 146376
rect 109696 132466 110368 132494
rect 110340 106321 110368 132466
rect 110326 106312 110382 106321
rect 110326 106247 110382 106256
rect 111076 89690 111104 150447
rect 111168 148374 111196 151786
rect 113916 151778 113968 151784
rect 112904 151768 112956 151774
rect 112904 151710 112956 151716
rect 112720 151292 112772 151298
rect 112720 151234 112772 151240
rect 112628 151224 112680 151230
rect 112628 151166 112680 151172
rect 112536 151156 112588 151162
rect 112536 151098 112588 151104
rect 112444 151020 112496 151026
rect 112444 150962 112496 150968
rect 111708 150952 111760 150958
rect 111708 150894 111760 150900
rect 111616 150884 111668 150890
rect 111616 150826 111668 150832
rect 111524 150816 111576 150822
rect 111524 150758 111576 150764
rect 111432 150748 111484 150754
rect 111432 150690 111484 150696
rect 111248 150680 111300 150686
rect 111248 150622 111300 150628
rect 111338 150648 111394 150657
rect 111156 148368 111208 148374
rect 111156 148310 111208 148316
rect 111260 148186 111288 150622
rect 111338 150583 111394 150592
rect 111168 148158 111288 148186
rect 111168 109002 111196 148158
rect 111352 148050 111380 150583
rect 111260 148022 111380 148050
rect 111156 108996 111208 109002
rect 111156 108938 111208 108944
rect 111260 92478 111288 148022
rect 111444 147914 111472 150690
rect 111352 147886 111472 147914
rect 111352 111790 111380 147886
rect 111536 147778 111564 150758
rect 111444 147750 111564 147778
rect 111444 113150 111472 147750
rect 111628 147642 111656 150826
rect 111536 147614 111656 147642
rect 111536 114510 111564 147614
rect 111720 147506 111748 150894
rect 111628 147478 111748 147506
rect 111628 117298 111656 147478
rect 111706 147384 111762 147393
rect 111706 147319 111762 147328
rect 111720 121446 111748 147319
rect 111708 121440 111760 121446
rect 111708 121382 111760 121388
rect 112456 118658 112484 150962
rect 112548 122806 112576 151098
rect 112640 124166 112668 151166
rect 112732 126954 112760 151234
rect 112812 150340 112864 150346
rect 112812 150282 112864 150288
rect 112824 132462 112852 150282
rect 112916 133890 112944 151710
rect 116032 151700 116084 151706
rect 116032 151642 116084 151648
rect 115296 151632 115348 151638
rect 115296 151574 115348 151580
rect 113088 151564 113140 151570
rect 113088 151506 113140 151512
rect 112996 150612 113048 150618
rect 112996 150554 113048 150560
rect 113008 137970 113036 150554
rect 113100 140758 113128 151506
rect 115204 150544 115256 150550
rect 115204 150486 115256 150492
rect 113822 144256 113878 144265
rect 113822 144191 113878 144200
rect 113088 140752 113140 140758
rect 113088 140694 113140 140700
rect 112996 137964 113048 137970
rect 112996 137906 113048 137912
rect 112904 133884 112956 133890
rect 112904 133826 112956 133832
rect 112812 132456 112864 132462
rect 112812 132398 112864 132404
rect 112720 126948 112772 126954
rect 112720 126890 112772 126896
rect 112628 124160 112680 124166
rect 112628 124102 112680 124108
rect 112536 122800 112588 122806
rect 112536 122742 112588 122748
rect 112444 118652 112496 118658
rect 112444 118594 112496 118600
rect 111616 117292 111668 117298
rect 111616 117234 111668 117240
rect 111524 114504 111576 114510
rect 111524 114446 111576 114452
rect 111432 113144 111484 113150
rect 111432 113086 111484 113092
rect 111340 111784 111392 111790
rect 111340 111726 111392 111732
rect 111248 92472 111300 92478
rect 111248 92414 111300 92420
rect 111064 89684 111116 89690
rect 111064 89626 111116 89632
rect 113836 88330 113864 144191
rect 115216 135561 115244 150486
rect 115308 141409 115336 151574
rect 116044 143313 116072 151642
rect 116952 151496 117004 151502
rect 116952 151438 117004 151444
rect 116768 151428 116820 151434
rect 116768 151370 116820 151376
rect 116676 151360 116728 151366
rect 116676 151302 116728 151308
rect 116124 150476 116176 150482
rect 116124 150418 116176 150424
rect 116136 145217 116164 150418
rect 116492 150068 116544 150074
rect 116492 150010 116544 150016
rect 116122 145208 116178 145217
rect 116122 145143 116178 145152
rect 116030 143304 116086 143313
rect 116030 143239 116086 143248
rect 115294 141400 115350 141409
rect 115294 141335 115350 141344
rect 116124 140752 116176 140758
rect 116124 140694 116176 140700
rect 116136 139505 116164 140694
rect 116122 139496 116178 139505
rect 116122 139431 116178 139440
rect 116124 137964 116176 137970
rect 116124 137906 116176 137912
rect 116136 137601 116164 137906
rect 116122 137592 116178 137601
rect 116122 137527 116178 137536
rect 115202 135552 115258 135561
rect 115202 135487 115258 135496
rect 116032 133884 116084 133890
rect 116032 133826 116084 133832
rect 116044 133657 116072 133826
rect 116030 133648 116086 133657
rect 116030 133583 116086 133592
rect 114190 132832 114246 132841
rect 114190 132767 114246 132776
rect 114204 132666 114232 132767
rect 114192 132660 114244 132666
rect 114192 132602 114244 132608
rect 115204 132660 115256 132666
rect 115204 132602 115256 132608
rect 113914 121408 113970 121417
rect 113914 121343 113970 121352
rect 113824 88324 113876 88330
rect 113824 88266 113876 88272
rect 113928 83978 113956 121343
rect 114006 110120 114062 110129
rect 114006 110055 114062 110064
rect 113916 83972 113968 83978
rect 113916 83914 113968 83920
rect 114020 82822 114048 110055
rect 114098 98696 114154 98705
rect 114098 98631 114154 98640
rect 114008 82816 114060 82822
rect 114008 82758 114060 82764
rect 114112 80034 114140 98631
rect 114190 87272 114246 87281
rect 114190 87207 114246 87216
rect 114100 80028 114152 80034
rect 114100 79970 114152 79976
rect 114204 78674 114232 87207
rect 115216 85649 115244 132602
rect 116124 132456 116176 132462
rect 116124 132398 116176 132404
rect 116136 131753 116164 132398
rect 116122 131744 116178 131753
rect 116122 131679 116178 131688
rect 116504 129849 116532 150010
rect 116582 149696 116638 149705
rect 116582 149631 116638 149640
rect 116490 129840 116546 129849
rect 116490 129775 116546 129784
rect 116124 126948 116176 126954
rect 116124 126890 116176 126896
rect 116136 126041 116164 126890
rect 116122 126032 116178 126041
rect 116122 125967 116178 125976
rect 116124 124160 116176 124166
rect 116122 124128 116124 124137
rect 116176 124128 116178 124137
rect 116122 124063 116178 124072
rect 115940 122800 115992 122806
rect 115940 122742 115992 122748
rect 115952 122233 115980 122742
rect 115938 122224 115994 122233
rect 115938 122159 115994 122168
rect 116124 121440 116176 121446
rect 116124 121382 116176 121388
rect 116136 120193 116164 121382
rect 116122 120184 116178 120193
rect 116122 120119 116178 120128
rect 116124 118652 116176 118658
rect 116124 118594 116176 118600
rect 116136 118289 116164 118594
rect 116122 118280 116178 118289
rect 116122 118215 116178 118224
rect 116124 117292 116176 117298
rect 116124 117234 116176 117240
rect 116136 116385 116164 117234
rect 116122 116376 116178 116385
rect 116122 116311 116178 116320
rect 116124 114504 116176 114510
rect 116122 114472 116124 114481
rect 116176 114472 116178 114481
rect 116122 114407 116178 114416
rect 115940 113144 115992 113150
rect 115940 113086 115992 113092
rect 115952 112577 115980 113086
rect 115938 112568 115994 112577
rect 115938 112503 115994 112512
rect 116124 111784 116176 111790
rect 116124 111726 116176 111732
rect 116136 110673 116164 111726
rect 116122 110664 116178 110673
rect 116122 110599 116178 110608
rect 116124 108996 116176 109002
rect 116124 108938 116176 108944
rect 116136 108769 116164 108938
rect 116122 108760 116178 108769
rect 116122 108695 116178 108704
rect 116596 93401 116624 149631
rect 116688 95305 116716 151302
rect 116780 97209 116808 151370
rect 116860 150204 116912 150210
rect 116860 150146 116912 150152
rect 116872 99113 116900 150146
rect 116964 102921 116992 151438
rect 117136 150272 117188 150278
rect 117136 150214 117188 150220
rect 117044 148368 117096 148374
rect 117044 148310 117096 148316
rect 116950 102912 117006 102921
rect 116950 102847 117006 102856
rect 117056 101017 117084 148310
rect 117148 104825 117176 150214
rect 117228 150136 117280 150142
rect 117228 150078 117280 150084
rect 117240 132546 117268 150078
rect 118896 149954 118924 157966
rect 119632 153882 119660 158714
rect 120172 156664 120224 156670
rect 120172 156606 120224 156612
rect 119528 153876 119580 153882
rect 119528 153818 119580 153824
rect 119620 153876 119672 153882
rect 119620 153818 119672 153824
rect 119540 149954 119568 153818
rect 120184 149954 120212 156606
rect 120644 152454 120672 163200
rect 121472 156058 121500 163200
rect 121644 158976 121696 158982
rect 121644 158918 121696 158924
rect 121460 156052 121512 156058
rect 121460 155994 121512 156000
rect 121656 153785 121684 158918
rect 122300 155446 122328 163200
rect 123128 159458 123156 163200
rect 123116 159452 123168 159458
rect 123116 159394 123168 159400
rect 122748 159384 122800 159390
rect 122748 159326 122800 159332
rect 122760 158030 122788 159326
rect 124048 158982 124076 163200
rect 124036 158976 124088 158982
rect 124036 158918 124088 158924
rect 122748 158024 122800 158030
rect 122748 157966 122800 157972
rect 123392 158024 123444 158030
rect 123392 157966 123444 157972
rect 122012 155440 122064 155446
rect 122012 155382 122064 155388
rect 122288 155440 122340 155446
rect 122288 155382 122340 155388
rect 121458 153776 121514 153785
rect 121458 153711 121514 153720
rect 121642 153776 121698 153785
rect 121642 153711 121698 153720
rect 120816 152516 120868 152522
rect 120816 152458 120868 152464
rect 120632 152448 120684 152454
rect 120632 152390 120684 152396
rect 120828 149954 120856 152458
rect 121000 152448 121052 152454
rect 121000 152390 121052 152396
rect 121012 151842 121040 152390
rect 121000 151836 121052 151842
rect 121000 151778 121052 151784
rect 121472 149954 121500 153711
rect 122024 149954 122052 155382
rect 122932 155236 122984 155242
rect 122932 155178 122984 155184
rect 122944 149954 122972 155178
rect 123404 149954 123432 157966
rect 124876 155990 124904 163200
rect 125508 158908 125560 158914
rect 125508 158850 125560 158856
rect 124864 155984 124916 155990
rect 124864 155926 124916 155932
rect 124588 155372 124640 155378
rect 124588 155314 124640 155320
rect 124220 153944 124272 153950
rect 124220 153886 124272 153892
rect 124232 149954 124260 153886
rect 124600 149954 124628 155314
rect 125520 153950 125548 158850
rect 125600 155304 125652 155310
rect 125600 155246 125652 155252
rect 125508 153944 125560 153950
rect 125508 153886 125560 153892
rect 125612 150226 125640 155246
rect 125704 155242 125732 163200
rect 126532 159730 126560 163200
rect 126428 159724 126480 159730
rect 126428 159666 126480 159672
rect 126520 159724 126572 159730
rect 126520 159666 126572 159672
rect 126440 159526 126468 159666
rect 126336 159520 126388 159526
rect 126336 159462 126388 159468
rect 126428 159520 126480 159526
rect 126428 159462 126480 159468
rect 126348 159372 126376 159462
rect 126532 159446 127020 159474
rect 126532 159372 126560 159446
rect 126992 159390 127020 159446
rect 126348 159344 126560 159372
rect 126888 159384 126940 159390
rect 126888 159326 126940 159332
rect 126980 159384 127032 159390
rect 126980 159326 127032 159332
rect 125692 155236 125744 155242
rect 125692 155178 125744 155184
rect 126612 154012 126664 154018
rect 126612 153954 126664 153960
rect 125966 152416 126022 152425
rect 125966 152351 126022 152360
rect 125612 150198 125686 150226
rect 118896 149926 119324 149954
rect 119540 149926 119876 149954
rect 120184 149926 120520 149954
rect 120828 149926 121164 149954
rect 121472 149926 121808 149954
rect 122024 149926 122452 149954
rect 122944 149926 123096 149954
rect 123404 149926 123740 149954
rect 124232 149926 124384 149954
rect 124600 149926 125028 149954
rect 125658 149940 125686 150198
rect 125980 149954 126008 152351
rect 126624 149954 126652 153954
rect 126900 152425 126928 159326
rect 127360 158914 127388 163200
rect 127624 159520 127676 159526
rect 127624 159462 127676 159468
rect 127348 158908 127400 158914
rect 127348 158850 127400 158856
rect 127164 156800 127216 156806
rect 127164 156742 127216 156748
rect 126886 152416 126942 152425
rect 126886 152351 126942 152360
rect 127176 149954 127204 156742
rect 127636 154018 127664 159462
rect 127992 158908 128044 158914
rect 127992 158850 128044 158856
rect 127624 154012 127676 154018
rect 127624 153954 127676 153960
rect 128004 152318 128032 158850
rect 128188 156670 128216 163200
rect 128176 156664 128228 156670
rect 128176 156606 128228 156612
rect 129016 155310 129044 163200
rect 129936 159526 129964 163200
rect 129924 159520 129976 159526
rect 129924 159462 129976 159468
rect 130660 159384 130712 159390
rect 130660 159326 130712 159332
rect 129832 156732 129884 156738
rect 129832 156674 129884 156680
rect 129004 155304 129056 155310
rect 129004 155246 129056 155252
rect 129188 154080 129240 154086
rect 129188 154022 129240 154028
rect 128634 152552 128690 152561
rect 128634 152487 128690 152496
rect 127900 152312 127952 152318
rect 127900 152254 127952 152260
rect 127992 152312 128044 152318
rect 127992 152254 128044 152260
rect 127912 149954 127940 152254
rect 128648 149954 128676 152487
rect 129200 149954 129228 154022
rect 129844 149954 129872 156674
rect 130672 151910 130700 159326
rect 130764 158914 130792 163200
rect 131026 159352 131082 159361
rect 131026 159287 131082 159296
rect 130752 158908 130804 158914
rect 130752 158850 130804 158856
rect 130476 151904 130528 151910
rect 130476 151846 130528 151852
rect 130660 151904 130712 151910
rect 130660 151846 130712 151852
rect 130488 149954 130516 151846
rect 131040 151824 131068 159287
rect 131592 158030 131620 163200
rect 131580 158024 131632 158030
rect 131580 157966 131632 157972
rect 132420 154057 132448 163200
rect 133144 159384 133196 159390
rect 133144 159326 133196 159332
rect 133156 158846 133184 159326
rect 133248 158846 133276 163200
rect 133786 159488 133842 159497
rect 133786 159423 133842 159432
rect 133144 158840 133196 158846
rect 133144 158782 133196 158788
rect 133236 158840 133288 158846
rect 133236 158782 133288 158788
rect 132500 156936 132552 156942
rect 132500 156878 132552 156884
rect 131762 154048 131818 154057
rect 131762 153983 131818 153992
rect 132406 154048 132462 154057
rect 132406 153983 132462 153992
rect 131040 151796 131160 151824
rect 131132 149954 131160 151796
rect 131776 149954 131804 153983
rect 132512 149954 132540 156878
rect 133052 154828 133104 154834
rect 133052 154770 133104 154776
rect 132868 154216 132920 154222
rect 132604 154164 132868 154170
rect 132604 154158 132920 154164
rect 132604 154154 132908 154158
rect 132592 154148 132908 154154
rect 132644 154142 132908 154148
rect 132592 154090 132644 154096
rect 133064 149954 133092 154770
rect 133144 154216 133196 154222
rect 133144 154158 133196 154164
rect 133156 153950 133184 154158
rect 133234 154048 133290 154057
rect 133234 153983 133290 153992
rect 133248 153950 133276 153983
rect 133144 153944 133196 153950
rect 133144 153886 133196 153892
rect 133236 153944 133288 153950
rect 133236 153886 133288 153892
rect 133800 151881 133828 159423
rect 134076 152590 134104 163200
rect 134904 156738 134932 163200
rect 135824 156874 135852 163200
rect 136652 163146 136680 163200
rect 136744 163146 136772 163254
rect 136652 163118 136772 163146
rect 137388 159798 137416 163254
rect 137466 163200 137522 164400
rect 138294 163200 138350 164400
rect 139122 163200 139178 164400
rect 139950 163200 140006 164400
rect 140778 163200 140834 164400
rect 141698 163200 141754 164400
rect 142526 163200 142582 164400
rect 143354 163200 143410 164400
rect 144182 163200 144238 164400
rect 145010 163200 145066 164400
rect 145838 163200 145894 164400
rect 146666 163200 146722 164400
rect 147586 163200 147642 164400
rect 148414 163200 148470 164400
rect 149242 163200 149298 164400
rect 150070 163200 150126 164400
rect 150898 163200 150954 164400
rect 151726 163200 151782 164400
rect 152554 163200 152610 164400
rect 153474 163200 153530 164400
rect 154302 163200 154358 164400
rect 155130 163200 155186 164400
rect 155958 163200 156014 164400
rect 156786 163200 156842 164400
rect 157614 163200 157670 164400
rect 158442 163200 158498 164400
rect 159362 163200 159418 164400
rect 160190 163200 160246 164400
rect 161018 163200 161074 164400
rect 161846 163200 161902 164400
rect 162674 163200 162730 164400
rect 163502 163200 163558 164400
rect 164330 163200 164386 164400
rect 165250 163200 165306 164400
rect 166078 163200 166134 164400
rect 166906 163200 166962 164400
rect 167734 163200 167790 164400
rect 168562 163200 168618 164400
rect 169390 163200 169446 164400
rect 170218 163200 170274 164400
rect 171138 163200 171194 164400
rect 171966 163200 172022 164400
rect 172794 163200 172850 164400
rect 173622 163200 173678 164400
rect 174450 163200 174506 164400
rect 175278 163200 175334 164400
rect 176106 163200 176162 164400
rect 177026 163200 177082 164400
rect 177854 163200 177910 164400
rect 178682 163200 178738 164400
rect 179510 163200 179566 164400
rect 180338 163200 180394 164400
rect 181166 163200 181222 164400
rect 181994 163200 182050 164400
rect 182914 163200 182970 164400
rect 183742 163200 183798 164400
rect 184570 163200 184626 164400
rect 185398 163200 185454 164400
rect 186226 163200 186282 164400
rect 187054 163200 187110 164400
rect 187882 163200 187938 164400
rect 188802 163200 188858 164400
rect 189630 163200 189686 164400
rect 190458 163200 190514 164400
rect 191286 163200 191342 164400
rect 192114 163200 192170 164400
rect 192942 163200 192998 164400
rect 193770 163200 193826 164400
rect 194690 163200 194746 164400
rect 195518 163200 195574 164400
rect 196346 163200 196402 164400
rect 197174 163200 197230 164400
rect 198002 163200 198058 164400
rect 198830 163200 198886 164400
rect 199658 163200 199714 164400
rect 200578 163200 200634 164400
rect 201406 163200 201462 164400
rect 202234 163200 202290 164400
rect 203062 163200 203118 164400
rect 203890 163200 203946 164400
rect 204718 163200 204774 164400
rect 205546 163200 205602 164400
rect 206466 163200 206522 164400
rect 207294 163200 207350 164400
rect 208122 163200 208178 164400
rect 208950 163200 209006 164400
rect 209778 163200 209834 164400
rect 210606 163200 210662 164400
rect 211434 163200 211490 164400
rect 212354 163200 212410 164400
rect 213182 163200 213238 164400
rect 214010 163200 214066 164400
rect 214838 163200 214894 164400
rect 215666 163200 215722 164400
rect 216494 163200 216550 164400
rect 217322 163200 217378 164400
rect 218242 163200 218298 164400
rect 219070 163200 219126 164400
rect 219176 163254 219388 163282
rect 137284 159792 137336 159798
rect 137284 159734 137336 159740
rect 137376 159792 137428 159798
rect 137376 159734 137428 159740
rect 137296 159594 137324 159734
rect 137100 159588 137152 159594
rect 137100 159530 137152 159536
rect 137284 159588 137336 159594
rect 137284 159530 137336 159536
rect 135260 156868 135312 156874
rect 135260 156810 135312 156816
rect 135812 156868 135864 156874
rect 135812 156810 135864 156816
rect 134892 156732 134944 156738
rect 134892 156674 134944 156680
rect 134338 153912 134394 153921
rect 134338 153847 134394 153856
rect 133880 152584 133932 152590
rect 133880 152526 133932 152532
rect 134064 152584 134116 152590
rect 134064 152526 134116 152532
rect 133786 151872 133842 151881
rect 133786 151807 133842 151816
rect 133892 149954 133920 152526
rect 134352 149954 134380 153847
rect 135272 150226 135300 156810
rect 136916 154080 136968 154086
rect 136916 154022 136968 154028
rect 135628 152652 135680 152658
rect 135628 152594 135680 152600
rect 135272 150198 135346 150226
rect 125980 149926 126316 149954
rect 126624 149926 126960 149954
rect 127176 149926 127604 149954
rect 127912 149926 128248 149954
rect 128648 149926 128892 149954
rect 129200 149926 129536 149954
rect 129844 149926 130180 149954
rect 130488 149926 130824 149954
rect 131132 149926 131468 149954
rect 131776 149926 132112 149954
rect 132512 149926 132756 149954
rect 133064 149926 133400 149954
rect 133892 149926 134044 149954
rect 134352 149926 134688 149954
rect 135318 149940 135346 150198
rect 135640 149954 135668 152594
rect 136270 151872 136326 151881
rect 136270 151807 136326 151816
rect 136284 149954 136312 151807
rect 136928 149954 136956 154022
rect 137112 152658 137140 159530
rect 137480 159390 137508 163200
rect 138018 159624 138074 159633
rect 138018 159559 138074 159568
rect 137376 159384 137428 159390
rect 137376 159326 137428 159332
rect 137468 159384 137520 159390
rect 137468 159326 137520 159332
rect 137388 154086 137416 159326
rect 137560 157004 137612 157010
rect 137560 156946 137612 156952
rect 137376 154080 137428 154086
rect 137376 154022 137428 154028
rect 137100 152652 137152 152658
rect 137100 152594 137152 152600
rect 137572 149954 137600 156946
rect 138032 151842 138060 159559
rect 138308 156942 138336 163200
rect 138296 156936 138348 156942
rect 138296 156878 138348 156884
rect 139136 156806 139164 163200
rect 139584 159792 139636 159798
rect 139584 159734 139636 159740
rect 139860 159792 139912 159798
rect 139860 159734 139912 159740
rect 139124 156800 139176 156806
rect 139124 156742 139176 156748
rect 139308 154964 139360 154970
rect 139308 154906 139360 154912
rect 138848 152788 138900 152794
rect 138848 152730 138900 152736
rect 138296 151972 138348 151978
rect 138296 151914 138348 151920
rect 138020 151836 138072 151842
rect 138020 151778 138072 151784
rect 138308 149954 138336 151914
rect 138860 149954 138888 152730
rect 139320 151978 139348 154906
rect 139596 154154 139624 159734
rect 139872 159594 139900 159734
rect 139964 159594 139992 163200
rect 139860 159588 139912 159594
rect 139860 159530 139912 159536
rect 139952 159588 140004 159594
rect 139952 159530 140004 159536
rect 140792 157334 140820 163200
rect 141712 157418 141740 163200
rect 141884 160064 141936 160070
rect 141884 160006 141936 160012
rect 141896 159526 141924 160006
rect 141884 159520 141936 159526
rect 141884 159462 141936 159468
rect 141700 157412 141752 157418
rect 141700 157354 141752 157360
rect 140792 157306 140912 157334
rect 140134 156632 140190 156641
rect 140134 156567 140190 156576
rect 139492 154148 139544 154154
rect 139492 154090 139544 154096
rect 139584 154148 139636 154154
rect 139584 154090 139636 154096
rect 139308 151972 139360 151978
rect 139308 151914 139360 151920
rect 139504 149954 139532 154090
rect 140148 149954 140176 156567
rect 140884 152726 140912 157306
rect 142540 155378 142568 163200
rect 143368 159662 143396 163200
rect 143264 159656 143316 159662
rect 143264 159598 143316 159604
rect 143356 159656 143408 159662
rect 143356 159598 143408 159604
rect 142710 156768 142766 156777
rect 142710 156703 142766 156712
rect 142528 155372 142580 155378
rect 142528 155314 142580 155320
rect 142528 154488 142580 154494
rect 142528 154430 142580 154436
rect 142620 154488 142672 154494
rect 142620 154430 142672 154436
rect 142158 154184 142214 154193
rect 142158 154119 142214 154128
rect 142344 154148 142396 154154
rect 140780 152720 140832 152726
rect 140780 152662 140832 152668
rect 140872 152720 140924 152726
rect 140872 152662 140924 152668
rect 140792 149954 140820 152662
rect 141424 151836 141476 151842
rect 141424 151778 141476 151784
rect 141436 149954 141464 151778
rect 142172 149954 142200 154119
rect 142344 154090 142396 154096
rect 142356 154057 142384 154090
rect 142342 154048 142398 154057
rect 142540 154018 142568 154430
rect 142632 154222 142660 154430
rect 142620 154216 142672 154222
rect 142620 154158 142672 154164
rect 142342 153983 142398 153992
rect 142436 154012 142488 154018
rect 142436 153954 142488 153960
rect 142528 154012 142580 154018
rect 142528 153954 142580 153960
rect 142448 153270 142476 153954
rect 142344 153264 142396 153270
rect 142344 153206 142396 153212
rect 142436 153264 142488 153270
rect 142436 153206 142488 153212
rect 142356 152794 142384 153206
rect 142344 152788 142396 152794
rect 142344 152730 142396 152736
rect 142252 152652 142304 152658
rect 142252 152594 142304 152600
rect 142264 151842 142292 152594
rect 142252 151836 142304 151842
rect 142252 151778 142304 151784
rect 142724 149954 142752 156703
rect 142804 154420 142856 154426
rect 142804 154362 142856 154368
rect 142896 154420 142948 154426
rect 142896 154362 142948 154368
rect 142816 154222 142844 154362
rect 142804 154216 142856 154222
rect 142804 154158 142856 154164
rect 142908 154086 142936 154362
rect 142896 154080 142948 154086
rect 142896 154022 142948 154028
rect 143078 154048 143134 154057
rect 143078 153983 143080 153992
rect 143132 153983 143134 153992
rect 143080 153954 143132 153960
rect 143276 152726 143304 159598
rect 144196 159526 144224 163200
rect 144920 160132 144972 160138
rect 144920 160074 144972 160080
rect 144932 159798 144960 160074
rect 144828 159792 144880 159798
rect 144828 159734 144880 159740
rect 144920 159792 144972 159798
rect 144920 159734 144972 159740
rect 144184 159520 144236 159526
rect 144184 159462 144236 159468
rect 144840 152862 144868 159734
rect 144918 157992 144974 158001
rect 144918 157927 144974 157936
rect 144000 152856 144052 152862
rect 144000 152798 144052 152804
rect 144828 152856 144880 152862
rect 144828 152798 144880 152804
rect 143264 152720 143316 152726
rect 143264 152662 143316 152668
rect 143538 152416 143594 152425
rect 143538 152351 143594 152360
rect 143552 149954 143580 152351
rect 144012 149954 144040 152798
rect 144932 150226 144960 157927
rect 145024 157078 145052 163200
rect 145852 157334 145880 163200
rect 146680 159798 146708 163200
rect 146484 159792 146536 159798
rect 146484 159734 146536 159740
rect 146668 159792 146720 159798
rect 146668 159734 146720 159740
rect 145852 157306 145972 157334
rect 145012 157072 145064 157078
rect 145012 157014 145064 157020
rect 145944 154970 145972 157306
rect 146024 157004 146076 157010
rect 146024 156946 146076 156952
rect 145932 154964 145984 154970
rect 145932 154906 145984 154912
rect 145288 152788 145340 152794
rect 145288 152730 145340 152736
rect 144932 150198 145006 150226
rect 135640 149926 135976 149954
rect 136284 149926 136620 149954
rect 136928 149926 137264 149954
rect 137572 149926 137908 149954
rect 138308 149926 138552 149954
rect 138860 149926 139196 149954
rect 139504 149926 139840 149954
rect 140148 149926 140484 149954
rect 140792 149926 141128 149954
rect 141436 149926 141772 149954
rect 142172 149926 142416 149954
rect 142724 149926 143060 149954
rect 143552 149926 143704 149954
rect 144012 149926 144348 149954
rect 144978 149940 145006 150198
rect 145300 149954 145328 152730
rect 146036 149954 146064 156946
rect 146496 154578 146524 159734
rect 147600 159610 147628 163200
rect 147508 159582 147628 159610
rect 147402 159488 147458 159497
rect 147402 159423 147404 159432
rect 147456 159423 147458 159432
rect 147404 159394 147456 159400
rect 147508 158778 147536 159582
rect 147678 159488 147734 159497
rect 147678 159423 147734 159432
rect 147404 158772 147456 158778
rect 147404 158714 147456 158720
rect 147496 158772 147548 158778
rect 147496 158714 147548 158720
rect 147128 158092 147180 158098
rect 147128 158034 147180 158040
rect 146496 154550 146708 154578
rect 146680 151910 146708 154550
rect 146576 151904 146628 151910
rect 146576 151846 146628 151852
rect 146668 151904 146720 151910
rect 146668 151846 146720 151852
rect 146588 149954 146616 151846
rect 147140 149954 147168 158034
rect 147416 157334 147444 158714
rect 147416 157306 147628 157334
rect 147600 154154 147628 157306
rect 147692 154290 147720 159423
rect 148428 158098 148456 163200
rect 149060 158772 149112 158778
rect 149060 158714 149112 158720
rect 148416 158092 148468 158098
rect 148416 158034 148468 158040
rect 148232 157208 148284 157214
rect 148232 157150 148284 157156
rect 147680 154284 147732 154290
rect 147680 154226 147732 154232
rect 147496 154148 147548 154154
rect 147496 154090 147548 154096
rect 147588 154148 147640 154154
rect 147588 154090 147640 154096
rect 147508 154057 147536 154090
rect 147494 154048 147550 154057
rect 147494 153983 147550 153992
rect 147862 154048 147918 154057
rect 147862 153983 147918 153992
rect 147876 149954 147904 153983
rect 148244 151814 148272 157150
rect 149072 152794 149100 158714
rect 149256 154834 149284 163200
rect 149610 158128 149666 158137
rect 149610 158063 149666 158072
rect 149244 154828 149296 154834
rect 149244 154770 149296 154776
rect 149060 152788 149112 152794
rect 149060 152730 149112 152736
rect 149152 152108 149204 152114
rect 149152 152050 149204 152056
rect 148244 151786 148456 151814
rect 148428 149954 148456 151786
rect 149164 149954 149192 152050
rect 149624 149954 149652 158063
rect 150084 157010 150112 163200
rect 150912 159458 150940 163200
rect 150900 159452 150952 159458
rect 150900 159394 150952 159400
rect 151740 157146 151768 163200
rect 152186 158264 152242 158273
rect 152186 158199 152242 158208
rect 150900 157140 150952 157146
rect 150900 157082 150952 157088
rect 151728 157140 151780 157146
rect 151728 157082 151780 157088
rect 150072 157004 150124 157010
rect 150072 156946 150124 156952
rect 150440 154216 150492 154222
rect 150440 154158 150492 154164
rect 150452 149954 150480 154158
rect 150912 149954 150940 157082
rect 151820 151836 151872 151842
rect 151820 151778 151872 151784
rect 151832 149954 151860 151778
rect 152200 149954 152228 158199
rect 152568 154222 152596 163200
rect 153488 159798 153516 163200
rect 153292 159792 153344 159798
rect 153292 159734 153344 159740
rect 153476 159792 153528 159798
rect 153476 159734 153528 159740
rect 153304 158778 153332 159734
rect 153292 158772 153344 158778
rect 153292 158714 153344 158720
rect 153476 157276 153528 157282
rect 153476 157218 153528 157224
rect 152556 154216 152608 154222
rect 152556 154158 152608 154164
rect 153200 154080 153252 154086
rect 153200 154022 153252 154028
rect 153212 150226 153240 154022
rect 153212 150198 153286 150226
rect 145300 149926 145636 149954
rect 146036 149926 146280 149954
rect 146588 149926 146924 149954
rect 147140 149926 147568 149954
rect 147876 149926 148212 149954
rect 148428 149926 148856 149954
rect 149164 149926 149500 149954
rect 149624 149926 150052 149954
rect 150452 149926 150696 149954
rect 150912 149926 151340 149954
rect 151832 149926 151984 149954
rect 152200 149926 152628 149954
rect 153258 149940 153286 150198
rect 153488 149954 153516 157218
rect 154212 152040 154264 152046
rect 154212 151982 154264 151988
rect 154224 149954 154252 151982
rect 154316 151842 154344 163200
rect 154488 160064 154540 160070
rect 154488 160006 154540 160012
rect 154500 154630 154528 160006
rect 155144 158166 155172 163200
rect 154764 158160 154816 158166
rect 154764 158102 154816 158108
rect 155132 158160 155184 158166
rect 155132 158102 155184 158108
rect 154488 154624 154540 154630
rect 154488 154566 154540 154572
rect 154304 151836 154356 151842
rect 154304 151778 154356 151784
rect 154776 149954 154804 158102
rect 155972 154766 156000 163200
rect 156800 160070 156828 163200
rect 156788 160064 156840 160070
rect 156788 160006 156840 160012
rect 156432 159854 156644 159882
rect 156328 159724 156380 159730
rect 156328 159666 156380 159672
rect 156340 157350 156368 159666
rect 156432 159662 156460 159854
rect 156616 159746 156644 159854
rect 156880 159860 156932 159866
rect 156880 159802 156932 159808
rect 156616 159718 156828 159746
rect 156800 159662 156828 159718
rect 156420 159656 156472 159662
rect 156420 159598 156472 159604
rect 156788 159656 156840 159662
rect 156788 159598 156840 159604
rect 156052 157344 156104 157350
rect 156052 157286 156104 157292
rect 156328 157344 156380 157350
rect 156328 157286 156380 157292
rect 155960 154760 156012 154766
rect 155960 154702 156012 154708
rect 154948 154556 155000 154562
rect 154948 154498 155000 154504
rect 154960 154086 154988 154498
rect 154948 154080 155000 154086
rect 154948 154022 155000 154028
rect 155500 153808 155552 153814
rect 155500 153750 155552 153756
rect 155512 149954 155540 153750
rect 156064 149954 156092 157286
rect 156420 154556 156472 154562
rect 156420 154498 156472 154504
rect 156604 154556 156656 154562
rect 156604 154498 156656 154504
rect 156328 154148 156380 154154
rect 156328 154090 156380 154096
rect 156340 153490 156368 154090
rect 156432 153814 156460 154498
rect 156616 154290 156644 154498
rect 156604 154284 156656 154290
rect 156604 154226 156656 154232
rect 156788 154216 156840 154222
rect 156788 154158 156840 154164
rect 156420 153808 156472 153814
rect 156800 153762 156828 154158
rect 156420 153750 156472 153756
rect 156524 153734 156828 153762
rect 156524 153678 156552 153734
rect 156512 153672 156564 153678
rect 156512 153614 156564 153620
rect 156604 153672 156656 153678
rect 156604 153614 156656 153620
rect 156616 153490 156644 153614
rect 156340 153462 156644 153490
rect 156788 152720 156840 152726
rect 156788 152662 156840 152668
rect 156800 149954 156828 152662
rect 156892 152114 156920 159802
rect 157628 159594 157656 163200
rect 157616 159588 157668 159594
rect 157616 159530 157668 159536
rect 158456 158234 158484 163200
rect 158720 158840 158772 158846
rect 158720 158782 158772 158788
rect 157340 158228 157392 158234
rect 157340 158170 157392 158176
rect 158444 158228 158496 158234
rect 158444 158170 158496 158176
rect 156880 152108 156932 152114
rect 156880 152050 156932 152056
rect 157352 149954 157380 158170
rect 158732 156602 158760 158782
rect 158628 156596 158680 156602
rect 158628 156538 158680 156544
rect 158720 156596 158772 156602
rect 158720 156538 158772 156544
rect 158640 156482 158668 156538
rect 158640 156454 158852 156482
rect 158076 154080 158128 154086
rect 158076 154022 158128 154028
rect 158088 149954 158116 154022
rect 158824 149954 158852 156454
rect 159376 154630 159404 163200
rect 160100 159656 160152 159662
rect 160100 159598 160152 159604
rect 160112 157214 160140 159598
rect 160100 157208 160152 157214
rect 160100 157150 160152 157156
rect 159364 154624 159416 154630
rect 159364 154566 159416 154572
rect 160204 154154 160232 163200
rect 161032 159662 161060 163200
rect 161020 159656 161072 159662
rect 161020 159598 161072 159604
rect 161860 158302 161888 163200
rect 162492 159928 162544 159934
rect 162492 159870 162544 159876
rect 160284 158296 160336 158302
rect 160284 158238 160336 158244
rect 161848 158296 161900 158302
rect 161848 158238 161900 158244
rect 160192 154148 160244 154154
rect 160192 154090 160244 154096
rect 159364 153196 159416 153202
rect 159364 153138 159416 153144
rect 159376 149954 159404 153138
rect 160296 150226 160324 158238
rect 161570 156904 161626 156913
rect 161570 156839 161626 156848
rect 160650 154320 160706 154329
rect 160650 154255 160706 154264
rect 160296 150198 160370 150226
rect 153488 149926 153916 149954
rect 154224 149926 154560 149954
rect 154776 149926 155204 149954
rect 155512 149926 155848 149954
rect 156064 149926 156492 149954
rect 156800 149926 157136 149954
rect 157352 149926 157780 149954
rect 158088 149926 158424 149954
rect 158824 149926 159068 149954
rect 159376 149926 159712 149954
rect 160342 149940 160370 150198
rect 160664 149954 160692 154255
rect 161584 150226 161612 156839
rect 161940 152856 161992 152862
rect 161940 152798 161992 152804
rect 161584 150198 161658 150226
rect 160664 149926 161000 149954
rect 161630 149940 161658 150198
rect 161952 149954 161980 152798
rect 162504 152046 162532 159870
rect 162688 154698 162716 163200
rect 163516 158846 163544 163200
rect 164344 161474 164372 163200
rect 164344 161446 164464 161474
rect 164148 159724 164200 159730
rect 164148 159666 164200 159672
rect 163504 158840 163556 158846
rect 163504 158782 163556 158788
rect 162858 158400 162914 158409
rect 162858 158335 162914 158344
rect 162676 154692 162728 154698
rect 162676 154634 162728 154640
rect 162492 152040 162544 152046
rect 162492 151982 162544 151988
rect 162872 150226 162900 158335
rect 164160 157298 164188 159666
rect 164160 157270 164372 157298
rect 164056 157208 164108 157214
rect 164056 157150 164108 157156
rect 164148 157208 164200 157214
rect 164148 157150 164200 157156
rect 164068 156534 164096 157150
rect 163780 156528 163832 156534
rect 163780 156470 163832 156476
rect 164056 156528 164108 156534
rect 164056 156470 164108 156476
rect 163228 154216 163280 154222
rect 163228 154158 163280 154164
rect 162872 150198 162946 150226
rect 161952 149926 162288 149954
rect 162918 149940 162946 150198
rect 163240 149954 163268 154158
rect 163792 149954 163820 156470
rect 164160 156466 164188 157150
rect 164344 156534 164372 157270
rect 164332 156528 164384 156534
rect 164332 156470 164384 156476
rect 164148 156460 164200 156466
rect 164148 156402 164200 156408
rect 164436 152862 164464 161446
rect 165264 158438 165292 163200
rect 165068 158432 165120 158438
rect 165068 158374 165120 158380
rect 165252 158432 165304 158438
rect 165252 158374 165304 158380
rect 164424 152856 164476 152862
rect 164424 152798 164476 152804
rect 164516 152176 164568 152182
rect 164516 152118 164568 152124
rect 164528 149954 164556 152118
rect 165080 149954 165108 158374
rect 166092 154222 166120 163200
rect 166920 159934 166948 163200
rect 166908 159928 166960 159934
rect 166908 159870 166960 159876
rect 166264 159860 166316 159866
rect 166264 159802 166316 159808
rect 166276 159118 166304 159802
rect 167748 159730 167776 163200
rect 167736 159724 167788 159730
rect 167736 159666 167788 159672
rect 167000 159316 167052 159322
rect 167000 159258 167052 159264
rect 166264 159112 166316 159118
rect 166264 159054 166316 159060
rect 166354 155544 166410 155553
rect 166354 155479 166410 155488
rect 166080 154216 166132 154222
rect 166080 154158 166132 154164
rect 165804 153740 165856 153746
rect 165804 153682 165856 153688
rect 165816 149954 165844 153682
rect 166368 149954 166396 155479
rect 167012 152182 167040 159258
rect 168576 158370 168604 163200
rect 167552 158364 167604 158370
rect 167552 158306 167604 158312
rect 168564 158364 168616 158370
rect 168564 158306 168616 158312
rect 167000 152176 167052 152182
rect 167000 152118 167052 152124
rect 167092 151904 167144 151910
rect 167092 151846 167144 151852
rect 167104 149954 167132 151846
rect 167564 151814 167592 158306
rect 169404 155514 169432 163200
rect 170232 159322 170260 163200
rect 170220 159316 170272 159322
rect 170220 159258 170272 159264
rect 171152 159186 171180 163200
rect 169944 159180 169996 159186
rect 169944 159122 169996 159128
rect 171140 159180 171192 159186
rect 171140 159122 171192 159128
rect 168380 155508 168432 155514
rect 168380 155450 168432 155456
rect 169392 155508 169444 155514
rect 169392 155450 169444 155456
rect 167564 151786 167684 151814
rect 167656 149954 167684 151786
rect 168392 149954 168420 155450
rect 168930 155272 168986 155281
rect 168930 155207 168986 155216
rect 168944 149954 168972 155207
rect 169760 152244 169812 152250
rect 169760 152186 169812 152192
rect 169772 149954 169800 152186
rect 169956 152182 169984 159122
rect 171980 158506 172008 163200
rect 172428 159860 172480 159866
rect 172428 159802 172480 159808
rect 170220 158500 170272 158506
rect 170220 158442 170272 158448
rect 171968 158500 172020 158506
rect 171968 158442 172020 158448
rect 169944 152176 169996 152182
rect 169944 152118 169996 152124
rect 170232 149954 170260 158442
rect 171600 157208 171652 157214
rect 171600 157150 171652 157156
rect 171230 155408 171286 155417
rect 171230 155343 171286 155352
rect 171244 150226 171272 155343
rect 171244 150198 171318 150226
rect 163240 149926 163576 149954
rect 163792 149926 164220 149954
rect 164528 149926 164864 149954
rect 165080 149926 165508 149954
rect 165816 149926 166152 149954
rect 166368 149926 166796 149954
rect 167104 149926 167440 149954
rect 167656 149926 168084 149954
rect 168392 149926 168728 149954
rect 168944 149926 169372 149954
rect 169772 149926 170016 149954
rect 170232 149926 170660 149954
rect 171290 149940 171318 150198
rect 171612 149954 171640 157150
rect 172440 152726 172468 159802
rect 172520 159180 172572 159186
rect 172520 159122 172572 159128
rect 172532 153202 172560 159122
rect 172704 158568 172756 158574
rect 172704 158510 172756 158516
rect 172520 153196 172572 153202
rect 172520 153138 172572 153144
rect 172428 152720 172480 152726
rect 172428 152662 172480 152668
rect 172520 152108 172572 152114
rect 172520 152050 172572 152056
rect 172532 150226 172560 152050
rect 172716 151814 172744 158510
rect 172808 154290 172836 163200
rect 173636 159186 173664 163200
rect 173624 159180 173676 159186
rect 173624 159122 173676 159128
rect 174360 159044 174412 159050
rect 174360 158986 174412 158992
rect 174372 158778 174400 158986
rect 174464 158778 174492 163200
rect 174360 158772 174412 158778
rect 174360 158714 174412 158720
rect 174452 158772 174504 158778
rect 174452 158714 174504 158720
rect 174912 158772 174964 158778
rect 174912 158714 174964 158720
rect 174082 157040 174138 157049
rect 174082 156975 174138 156984
rect 173072 155576 173124 155582
rect 173072 155518 173124 155524
rect 172796 154284 172848 154290
rect 172796 154226 172848 154232
rect 173084 151814 173112 155518
rect 172716 151786 172836 151814
rect 173084 151786 173480 151814
rect 172532 150198 172606 150226
rect 171612 149926 171948 149954
rect 172578 149940 172606 150198
rect 172808 149954 172836 151786
rect 173452 149954 173480 151786
rect 174096 149954 174124 156975
rect 174924 153066 174952 158714
rect 175292 158642 175320 163200
rect 176120 161474 176148 163200
rect 176120 161446 176332 161474
rect 175188 158636 175240 158642
rect 175188 158578 175240 158584
rect 175280 158636 175332 158642
rect 175280 158578 175332 158584
rect 175200 158522 175228 158578
rect 175200 158494 175320 158522
rect 174820 153060 174872 153066
rect 174820 153002 174872 153008
rect 174912 153060 174964 153066
rect 174912 153002 174964 153008
rect 174832 149954 174860 153002
rect 175292 151814 175320 158494
rect 176200 157956 176252 157962
rect 176200 157898 176252 157904
rect 175924 157888 175976 157894
rect 176212 157842 176240 157898
rect 175976 157836 176240 157842
rect 175924 157830 176240 157836
rect 175936 157814 176240 157830
rect 176016 155644 176068 155650
rect 176016 155586 176068 155592
rect 175292 151786 175412 151814
rect 175384 149954 175412 151786
rect 176028 149954 176056 155586
rect 176304 155582 176332 161446
rect 176660 159044 176712 159050
rect 176660 158986 176712 158992
rect 176292 155576 176344 155582
rect 176292 155518 176344 155524
rect 176672 153678 176700 158986
rect 177040 157214 177068 163200
rect 177868 159798 177896 163200
rect 177856 159792 177908 159798
rect 177856 159734 177908 159740
rect 178696 158574 178724 163200
rect 178684 158568 178736 158574
rect 178684 158510 178736 158516
rect 178040 157888 178092 157894
rect 178040 157830 178092 157836
rect 177028 157208 177080 157214
rect 177028 157150 177080 157156
rect 176842 155816 176898 155825
rect 176842 155751 176898 155760
rect 176660 153672 176712 153678
rect 176660 153614 176712 153620
rect 176108 152720 176160 152726
rect 176108 152662 176160 152668
rect 176120 152250 176148 152662
rect 176108 152244 176160 152250
rect 176108 152186 176160 152192
rect 176856 149954 176884 155751
rect 177396 152040 177448 152046
rect 177396 151982 177448 151988
rect 177408 149954 177436 151982
rect 178052 149954 178080 157830
rect 178682 155680 178738 155689
rect 179524 155650 179552 163200
rect 180352 158778 180380 163200
rect 180708 159860 180760 159866
rect 180708 159802 180760 159808
rect 180720 158794 180748 159802
rect 180340 158772 180392 158778
rect 180720 158766 180932 158794
rect 180340 158714 180392 158720
rect 180904 158710 180932 158766
rect 180800 158704 180852 158710
rect 180800 158646 180852 158652
rect 180892 158704 180944 158710
rect 180892 158646 180944 158652
rect 178682 155615 178738 155624
rect 179512 155644 179564 155650
rect 178696 149954 178724 155615
rect 179512 155586 179564 155592
rect 179420 153604 179472 153610
rect 179420 153546 179472 153552
rect 179432 149954 179460 153546
rect 179972 152380 180024 152386
rect 179972 152322 180024 152328
rect 179984 149954 180012 152322
rect 180812 150226 180840 158646
rect 181180 157334 181208 163200
rect 182008 158710 182036 163200
rect 181904 158704 181956 158710
rect 181904 158646 181956 158652
rect 181996 158704 182048 158710
rect 181996 158646 182048 158652
rect 181272 157950 181576 157978
rect 181272 157758 181300 157950
rect 181548 157894 181576 157950
rect 181536 157888 181588 157894
rect 181536 157830 181588 157836
rect 181628 157820 181680 157826
rect 181628 157762 181680 157768
rect 181812 157820 181864 157826
rect 181812 157762 181864 157768
rect 181260 157752 181312 157758
rect 181260 157694 181312 157700
rect 181640 157706 181668 157762
rect 181640 157690 181760 157706
rect 181536 157684 181588 157690
rect 181640 157684 181772 157690
rect 181640 157678 181720 157684
rect 181536 157626 181588 157632
rect 181720 157626 181772 157632
rect 181548 157570 181576 157626
rect 181824 157570 181852 157762
rect 181916 157758 181944 158646
rect 182824 157956 182876 157962
rect 182824 157898 182876 157904
rect 181904 157752 181956 157758
rect 181904 157694 181956 157700
rect 181548 157542 181852 157570
rect 181180 157306 181300 157334
rect 181168 155712 181220 155718
rect 181168 155654 181220 155660
rect 181076 154352 181128 154358
rect 181074 154320 181076 154329
rect 181128 154320 181130 154329
rect 181074 154255 181130 154264
rect 180812 150198 180886 150226
rect 172808 149926 173236 149954
rect 173452 149926 173880 149954
rect 174096 149926 174524 149954
rect 174832 149926 175168 149954
rect 175384 149926 175812 149954
rect 176028 149926 176456 149954
rect 176856 149926 177100 149954
rect 177408 149926 177744 149954
rect 178052 149926 178388 149954
rect 178696 149926 179032 149954
rect 179432 149926 179676 149954
rect 179984 149926 180320 149954
rect 180858 149940 180886 150198
rect 181180 149954 181208 155654
rect 181272 152386 181300 157306
rect 181812 156392 181864 156398
rect 181812 156334 181864 156340
rect 181444 154420 181496 154426
rect 181444 154362 181496 154368
rect 181456 154329 181484 154362
rect 181442 154320 181498 154329
rect 181442 154255 181498 154264
rect 181260 152380 181312 152386
rect 181260 152322 181312 152328
rect 181824 149954 181852 156334
rect 182456 152176 182508 152182
rect 182456 152118 182508 152124
rect 182468 149954 182496 152118
rect 182836 150090 182864 157898
rect 182928 153678 182956 163200
rect 183468 159112 183520 159118
rect 183468 159054 183520 159060
rect 182916 153672 182968 153678
rect 182916 153614 182968 153620
rect 183480 152182 183508 159054
rect 183756 159050 183784 163200
rect 184584 159866 184612 163200
rect 184572 159860 184624 159866
rect 184572 159802 184624 159808
rect 184664 159248 184716 159254
rect 184664 159190 184716 159196
rect 183744 159044 183796 159050
rect 183744 158986 183796 158992
rect 183742 155952 183798 155961
rect 183742 155887 183798 155896
rect 183468 152176 183520 152182
rect 183468 152118 183520 152124
rect 182836 150062 183048 150090
rect 183020 149954 183048 150062
rect 183756 149954 183784 155887
rect 184386 154456 184442 154465
rect 184386 154391 184442 154400
rect 184400 149954 184428 154391
rect 184676 152046 184704 159190
rect 185412 157962 185440 163200
rect 185400 157956 185452 157962
rect 185400 157898 185452 157904
rect 185584 157684 185636 157690
rect 185584 157626 185636 157632
rect 185032 152108 185084 152114
rect 185032 152050 185084 152056
rect 184664 152040 184716 152046
rect 184664 151982 184716 151988
rect 185044 149954 185072 152050
rect 185596 149954 185624 157626
rect 186240 155718 186268 163200
rect 186412 159928 186464 159934
rect 186412 159870 186464 159876
rect 186424 157334 186452 159870
rect 187068 159254 187096 163200
rect 187056 159248 187108 159254
rect 187056 159190 187108 159196
rect 186424 157306 186728 157334
rect 186412 155848 186464 155854
rect 186412 155790 186464 155796
rect 186228 155712 186280 155718
rect 186228 155654 186280 155660
rect 186318 155136 186374 155145
rect 186318 155071 186374 155080
rect 186332 155038 186360 155071
rect 186320 155032 186372 155038
rect 186320 154974 186372 154980
rect 186424 149954 186452 155790
rect 186700 154902 186728 157306
rect 186964 155916 187016 155922
rect 186964 155858 187016 155864
rect 186780 155100 186832 155106
rect 186780 155042 186832 155048
rect 186596 154896 186648 154902
rect 186596 154838 186648 154844
rect 186688 154896 186740 154902
rect 186688 154838 186740 154844
rect 186608 154714 186636 154838
rect 186792 154714 186820 155042
rect 186608 154686 186820 154714
rect 186976 149954 187004 155858
rect 187896 152930 187924 163200
rect 188816 157894 188844 163200
rect 188160 157888 188212 157894
rect 188160 157830 188212 157836
rect 188804 157888 188856 157894
rect 188804 157830 188856 157836
rect 187700 152924 187752 152930
rect 187700 152866 187752 152872
rect 187884 152924 187936 152930
rect 187884 152866 187936 152872
rect 187712 149954 187740 152866
rect 188172 149954 188200 157830
rect 189644 155854 189672 163200
rect 190472 157758 190500 163200
rect 191300 159934 191328 163200
rect 191748 160064 191800 160070
rect 191748 160006 191800 160012
rect 191656 159996 191708 160002
rect 191656 159938 191708 159944
rect 191288 159928 191340 159934
rect 191288 159870 191340 159876
rect 190644 157820 190696 157826
rect 190644 157762 190696 157768
rect 190460 157752 190512 157758
rect 190460 157694 190512 157700
rect 190656 157334 190684 157762
rect 190656 157306 190776 157334
rect 189632 155848 189684 155854
rect 189632 155790 189684 155796
rect 189080 155168 189132 155174
rect 189172 155168 189224 155174
rect 189080 155110 189132 155116
rect 189170 155136 189172 155145
rect 189224 155136 189226 155145
rect 189092 149954 189120 155110
rect 189170 155071 189226 155080
rect 189540 154420 189592 154426
rect 189540 154362 189592 154368
rect 189552 149954 189580 154362
rect 190184 152244 190236 152250
rect 190184 152186 190236 152192
rect 190196 149954 190224 152186
rect 190748 149954 190776 157306
rect 191472 155032 191524 155038
rect 191472 154974 191524 154980
rect 191024 154550 191328 154578
rect 191024 154494 191052 154550
rect 191012 154488 191064 154494
rect 191012 154430 191064 154436
rect 191196 154420 191248 154426
rect 191196 154362 191248 154368
rect 191208 153678 191236 154362
rect 191300 153678 191328 154550
rect 191380 154352 191432 154358
rect 191380 154294 191432 154300
rect 191196 153672 191248 153678
rect 191196 153614 191248 153620
rect 191288 153672 191340 153678
rect 191288 153614 191340 153620
rect 191392 153406 191420 154294
rect 191380 153400 191432 153406
rect 191380 153342 191432 153348
rect 191484 149954 191512 154974
rect 191668 152182 191696 159938
rect 191760 153406 191788 160006
rect 192128 157282 192156 163200
rect 192116 157276 192168 157282
rect 192116 157218 192168 157224
rect 192956 155922 192984 163200
rect 193784 159118 193812 163200
rect 193772 159112 193824 159118
rect 193772 159054 193824 159060
rect 194704 158982 194732 163200
rect 194508 158976 194560 158982
rect 194508 158918 194560 158924
rect 194692 158976 194744 158982
rect 194692 158918 194744 158924
rect 193220 157616 193272 157622
rect 193220 157558 193272 157564
rect 193232 157334 193260 157558
rect 193232 157306 193352 157334
rect 192944 155916 192996 155922
rect 192944 155858 192996 155864
rect 192114 153776 192170 153785
rect 192114 153711 192170 153720
rect 191748 153400 191800 153406
rect 191748 153342 191800 153348
rect 191656 152176 191708 152182
rect 191656 152118 191708 152124
rect 192128 149954 192156 153711
rect 192760 152992 192812 152998
rect 192760 152934 192812 152940
rect 192772 149954 192800 152934
rect 193324 149954 193352 157306
rect 194048 155168 194100 155174
rect 194048 155110 194100 155116
rect 194060 149954 194088 155110
rect 194520 152250 194548 158918
rect 194968 158908 195020 158914
rect 194968 158850 195020 158856
rect 194692 156256 194744 156262
rect 194692 156198 194744 156204
rect 194508 152244 194560 152250
rect 194508 152186 194560 152192
rect 194704 149954 194732 156198
rect 194980 152998 195008 158850
rect 195532 157826 195560 163200
rect 196072 158840 196124 158846
rect 196072 158782 196124 158788
rect 195520 157820 195572 157826
rect 195520 157762 195572 157768
rect 196084 157334 196112 158782
rect 196084 157306 196296 157334
rect 196164 156324 196216 156330
rect 196164 156266 196216 156272
rect 195980 153672 196032 153678
rect 195886 153640 195942 153649
rect 196072 153672 196124 153678
rect 195980 153614 196032 153620
rect 196070 153640 196072 153649
rect 196124 153640 196126 153649
rect 195886 153575 195942 153584
rect 195900 153406 195928 153575
rect 195992 153406 196020 153614
rect 196070 153575 196126 153584
rect 195888 153400 195940 153406
rect 195888 153342 195940 153348
rect 195980 153400 196032 153406
rect 195980 153342 196032 153348
rect 194968 152992 195020 152998
rect 194968 152934 195020 152940
rect 195336 152040 195388 152046
rect 195336 151982 195388 151988
rect 195348 149954 195376 151982
rect 196176 149954 196204 156266
rect 196268 154986 196296 157306
rect 196360 155174 196388 163200
rect 197188 160070 197216 163200
rect 197176 160064 197228 160070
rect 197176 160006 197228 160012
rect 198016 160002 198044 163200
rect 198004 159996 198056 160002
rect 198004 159938 198056 159944
rect 197360 159180 197412 159186
rect 197360 159122 197412 159128
rect 197372 157622 197400 159122
rect 198738 158536 198794 158545
rect 198738 158471 198794 158480
rect 197360 157616 197412 157622
rect 197360 157558 197412 157564
rect 196348 155168 196400 155174
rect 196348 155110 196400 155116
rect 196268 154958 196756 154986
rect 196728 153542 196756 154958
rect 196624 153536 196676 153542
rect 196624 153478 196676 153484
rect 196716 153536 196768 153542
rect 196716 153478 196768 153484
rect 196636 149954 196664 153478
rect 197280 153474 197676 153490
rect 197268 153468 197688 153474
rect 197320 153462 197636 153468
rect 197268 153410 197320 153416
rect 197636 153410 197688 153416
rect 197360 153400 197412 153406
rect 197360 153342 197412 153348
rect 197372 149954 197400 153342
rect 197912 153128 197964 153134
rect 197912 153070 197964 153076
rect 197924 149954 197952 153070
rect 198752 149954 198780 158471
rect 198844 156398 198872 163200
rect 199292 159316 199344 159322
rect 199292 159258 199344 159264
rect 198832 156392 198884 156398
rect 198832 156334 198884 156340
rect 199304 153474 199332 159258
rect 199672 155106 199700 163200
rect 200592 159050 200620 163200
rect 201420 159322 201448 163200
rect 201408 159316 201460 159322
rect 201408 159258 201460 159264
rect 200488 159044 200540 159050
rect 200488 158986 200540 158992
rect 200580 159044 200632 159050
rect 200580 158986 200632 158992
rect 199660 155100 199712 155106
rect 199660 155042 199712 155048
rect 200120 155032 200172 155038
rect 200120 154974 200172 154980
rect 199200 153468 199252 153474
rect 199200 153410 199252 153416
rect 199292 153468 199344 153474
rect 199292 153410 199344 153416
rect 199212 149954 199240 153410
rect 200132 150226 200160 154974
rect 200500 153542 200528 158986
rect 200948 156392 201000 156398
rect 200948 156334 201000 156340
rect 200764 156324 200816 156330
rect 200764 156266 200816 156272
rect 200672 156188 200724 156194
rect 200672 156130 200724 156136
rect 200488 153536 200540 153542
rect 200488 153478 200540 153484
rect 200488 152108 200540 152114
rect 200488 152050 200540 152056
rect 200132 150198 200206 150226
rect 181180 149926 181516 149954
rect 181824 149926 182160 149954
rect 182468 149926 182804 149954
rect 183020 149926 183448 149954
rect 183756 149926 184092 149954
rect 184400 149926 184736 149954
rect 185044 149926 185380 149954
rect 185596 149926 186024 149954
rect 186424 149926 186668 149954
rect 186976 149926 187312 149954
rect 187712 149926 187956 149954
rect 188172 149926 188600 149954
rect 189092 149926 189244 149954
rect 189552 149926 189888 149954
rect 190196 149926 190532 149954
rect 190748 149926 191176 149954
rect 191484 149926 191820 149954
rect 192128 149926 192464 149954
rect 192772 149926 193108 149954
rect 193324 149926 193752 149954
rect 194060 149926 194396 149954
rect 194704 149926 195040 149954
rect 195348 149926 195684 149954
rect 196176 149926 196328 149954
rect 196636 149926 196972 149954
rect 197372 149926 197616 149954
rect 197924 149926 198260 149954
rect 198752 149926 198904 149954
rect 199212 149926 199548 149954
rect 200178 149940 200206 150198
rect 200500 149954 200528 152050
rect 200684 150090 200712 156130
rect 200776 156058 200804 156266
rect 200960 156126 200988 156334
rect 200948 156120 201000 156126
rect 200948 156062 201000 156068
rect 202248 156058 202276 163200
rect 203076 156262 203104 163200
rect 203904 159186 203932 163200
rect 204732 159361 204760 163200
rect 204718 159352 204774 159361
rect 204718 159287 204774 159296
rect 203892 159180 203944 159186
rect 203892 159122 203944 159128
rect 203708 158976 203760 158982
rect 203708 158918 203760 158924
rect 203432 157548 203484 157554
rect 203432 157490 203484 157496
rect 203444 157334 203472 157490
rect 203444 157306 203656 157334
rect 203064 156256 203116 156262
rect 203064 156198 203116 156204
rect 200764 156052 200816 156058
rect 200764 155994 200816 156000
rect 202236 156052 202288 156058
rect 202236 155994 202288 156000
rect 202420 154488 202472 154494
rect 202420 154430 202472 154436
rect 201776 154352 201828 154358
rect 201776 154294 201828 154300
rect 200684 150062 201080 150090
rect 201052 149954 201080 150062
rect 201788 149954 201816 154294
rect 202432 149954 202460 154430
rect 203064 151972 203116 151978
rect 203064 151914 203116 151920
rect 203076 149954 203104 151914
rect 203628 149954 203656 157306
rect 203720 153134 203748 158918
rect 204904 158772 204956 158778
rect 204904 158714 204956 158720
rect 204916 157554 204944 158714
rect 204904 157548 204956 157554
rect 204904 157490 204956 157496
rect 204352 155780 204404 155786
rect 204352 155722 204404 155728
rect 203708 153128 203760 153134
rect 203708 153070 203760 153076
rect 204364 149954 204392 155722
rect 205560 154358 205588 163200
rect 206192 157480 206244 157486
rect 206192 157422 206244 157428
rect 205548 154352 205600 154358
rect 205548 154294 205600 154300
rect 204996 153264 205048 153270
rect 204996 153206 205048 153212
rect 205008 149954 205036 153206
rect 205640 152448 205692 152454
rect 205640 152390 205692 152396
rect 205652 149954 205680 152390
rect 206204 149954 206232 157422
rect 206480 155786 206508 163200
rect 207112 160064 207164 160070
rect 207112 160006 207164 160012
rect 207018 157176 207074 157185
rect 207018 157111 207074 157120
rect 206468 155780 206520 155786
rect 206468 155722 206520 155728
rect 207032 149954 207060 157111
rect 207124 155038 207152 160006
rect 207308 158846 207336 163200
rect 208136 158982 208164 163200
rect 208124 158976 208176 158982
rect 208124 158918 208176 158924
rect 207296 158840 207348 158846
rect 207296 158782 207348 158788
rect 208768 156188 208820 156194
rect 208768 156130 208820 156136
rect 207112 155032 207164 155038
rect 207112 154974 207164 154980
rect 207572 153332 207624 153338
rect 207572 153274 207624 153280
rect 207584 149954 207612 153274
rect 208400 152176 208452 152182
rect 208400 152118 208452 152124
rect 208412 149954 208440 152118
rect 208780 149954 208808 156130
rect 208964 154494 208992 163200
rect 209792 156398 209820 163200
rect 210620 158778 210648 163200
rect 211448 160070 211476 163200
rect 211436 160064 211488 160070
rect 211436 160006 211488 160012
rect 210608 158772 210660 158778
rect 210608 158714 210660 158720
rect 209780 156392 209832 156398
rect 209780 156334 209832 156340
rect 211344 156324 211396 156330
rect 211344 156266 211396 156272
rect 208952 154488 209004 154494
rect 208952 154430 209004 154436
rect 209780 153876 209832 153882
rect 209780 153818 209832 153824
rect 209792 150226 209820 153818
rect 210148 153740 210200 153746
rect 210148 153682 210200 153688
rect 209792 150198 209866 150226
rect 200500 149926 200836 149954
rect 201052 149926 201480 149954
rect 201788 149926 202124 149954
rect 202432 149926 202768 149954
rect 203076 149926 203412 149954
rect 203628 149926 204056 149954
rect 204364 149926 204700 149954
rect 205008 149926 205344 149954
rect 205652 149926 205988 149954
rect 206204 149926 206632 149954
rect 207032 149926 207276 149954
rect 207584 149926 207920 149954
rect 208412 149926 208564 149954
rect 208780 149926 209208 149954
rect 209838 149940 209866 150198
rect 210160 149954 210188 153682
rect 210792 152516 210844 152522
rect 210792 152458 210844 152464
rect 210804 149954 210832 152458
rect 211356 149954 211384 156266
rect 211988 155440 212040 155446
rect 211988 155382 212040 155388
rect 212000 149954 212028 155382
rect 212368 153785 212396 163200
rect 213092 159316 213144 159322
rect 213092 159258 213144 159264
rect 212448 158976 212500 158982
rect 212448 158918 212500 158924
rect 212354 153776 212410 153785
rect 212354 153711 212410 153720
rect 212460 152522 212488 158918
rect 212540 157344 212592 157350
rect 212540 157286 212592 157292
rect 212552 156330 212580 157286
rect 212540 156324 212592 156330
rect 212540 156266 212592 156272
rect 212724 154556 212776 154562
rect 212724 154498 212776 154504
rect 212448 152516 212500 152522
rect 212448 152458 212500 152464
rect 212736 149954 212764 154498
rect 213104 151978 213132 159258
rect 213196 157350 213224 163200
rect 214024 159322 214052 163200
rect 214012 159316 214064 159322
rect 214012 159258 214064 159264
rect 214104 159248 214156 159254
rect 214104 159190 214156 159196
rect 213644 159180 213696 159186
rect 213644 159122 213696 159128
rect 213184 157344 213236 157350
rect 213184 157286 213236 157292
rect 213276 152244 213328 152250
rect 213276 152186 213328 152192
rect 213092 151972 213144 151978
rect 213092 151914 213144 151920
rect 213288 149954 213316 152186
rect 213656 152182 213684 159122
rect 213920 155984 213972 155990
rect 213920 155926 213972 155932
rect 213644 152176 213696 152182
rect 213644 152118 213696 152124
rect 213932 149954 213960 155926
rect 214116 155446 214144 159190
rect 214852 158846 214880 163200
rect 214840 158840 214892 158846
rect 214840 158782 214892 158788
rect 215300 158772 215352 158778
rect 215300 158714 215352 158720
rect 214300 156058 214604 156074
rect 214288 156052 214616 156058
rect 214340 156046 214564 156052
rect 214288 155994 214340 156000
rect 214564 155994 214616 156000
rect 214104 155440 214156 155446
rect 214104 155382 214156 155388
rect 214472 155236 214524 155242
rect 214472 155178 214524 155184
rect 214484 149954 214512 155178
rect 215312 152454 215340 158714
rect 215392 156324 215444 156330
rect 215392 156266 215444 156272
rect 215300 152448 215352 152454
rect 215300 152390 215352 152396
rect 215404 149954 215432 156266
rect 215680 153882 215708 163200
rect 216508 156330 216536 163200
rect 217336 158914 217364 163200
rect 218256 159254 218284 163200
rect 219084 163146 219112 163200
rect 219176 163146 219204 163254
rect 219084 163118 219204 163146
rect 218244 159248 218296 159254
rect 218244 159190 218296 159196
rect 218060 159112 218112 159118
rect 218060 159054 218112 159060
rect 217324 158908 217376 158914
rect 217324 158850 217376 158856
rect 216680 156664 216732 156670
rect 216680 156606 216732 156612
rect 216496 156324 216548 156330
rect 216496 156266 216548 156272
rect 215668 153876 215720 153882
rect 215668 153818 215720 153824
rect 215852 152312 215904 152318
rect 215852 152254 215904 152260
rect 215864 149954 215892 152254
rect 216692 149954 216720 156606
rect 218072 156194 218100 159054
rect 218980 158024 219032 158030
rect 218980 157966 219032 157972
rect 218060 156188 218112 156194
rect 218060 156130 218112 156136
rect 217048 155304 217100 155310
rect 217048 155246 217100 155252
rect 217060 149954 217088 155246
rect 218060 153808 218112 153814
rect 218060 153750 218112 153756
rect 218072 150226 218100 153750
rect 218428 152992 218480 152998
rect 218428 152934 218480 152940
rect 218072 150198 218146 150226
rect 210160 149926 210496 149954
rect 210804 149926 211140 149954
rect 211356 149926 211692 149954
rect 212000 149926 212336 149954
rect 212736 149926 212980 149954
rect 213288 149926 213624 149954
rect 213932 149926 214268 149954
rect 214484 149926 214912 149954
rect 215404 149926 215556 149954
rect 215864 149926 216200 149954
rect 216692 149926 216844 149954
rect 217060 149926 217488 149954
rect 218118 149940 218146 150198
rect 218440 149954 218468 152934
rect 218992 149954 219020 157966
rect 219360 154562 219388 163254
rect 219898 163200 219954 164400
rect 220726 163200 220782 164400
rect 221554 163200 221610 164400
rect 222382 163200 222438 164400
rect 223210 163200 223266 164400
rect 224130 163200 224186 164400
rect 224958 163200 225014 164400
rect 225786 163200 225842 164400
rect 226614 163200 226670 164400
rect 227442 163200 227498 164400
rect 228270 163200 228326 164400
rect 229098 163200 229154 164400
rect 230018 163200 230074 164400
rect 230846 163200 230902 164400
rect 231674 163200 231730 164400
rect 232502 163200 232558 164400
rect 233330 163200 233386 164400
rect 234158 163200 234214 164400
rect 234264 163254 234568 163282
rect 219912 156262 219940 163200
rect 220740 159186 220768 163200
rect 220728 159180 220780 159186
rect 220728 159122 220780 159128
rect 220728 158908 220780 158914
rect 220728 158850 220780 158856
rect 219992 156596 220044 156602
rect 219992 156538 220044 156544
rect 219900 156256 219952 156262
rect 219900 156198 219952 156204
rect 219348 154556 219400 154562
rect 219348 154498 219400 154504
rect 219716 153944 219768 153950
rect 219716 153886 219768 153892
rect 219728 149954 219756 153886
rect 220004 151814 220032 156538
rect 220740 152726 220768 158850
rect 221568 158778 221596 163200
rect 221740 158840 221792 158846
rect 221740 158782 221792 158788
rect 221556 158772 221608 158778
rect 221556 158714 221608 158720
rect 221372 156732 221424 156738
rect 221372 156674 221424 156680
rect 220728 152720 220780 152726
rect 220728 152662 220780 152668
rect 221004 152584 221056 152590
rect 221004 152526 221056 152532
rect 220004 151786 220308 151814
rect 220280 149954 220308 151786
rect 221016 149954 221044 152526
rect 221384 151814 221412 156674
rect 221752 152250 221780 158782
rect 222200 156868 222252 156874
rect 222200 156810 222252 156816
rect 221740 152244 221792 152250
rect 221740 152186 221792 152192
rect 221384 151786 221596 151814
rect 221568 149954 221596 151786
rect 222212 149954 222240 156810
rect 222396 153950 222424 163200
rect 223224 156670 223252 163200
rect 223580 159384 223632 159390
rect 223580 159326 223632 159332
rect 223212 156664 223264 156670
rect 223212 156606 223264 156612
rect 222936 154012 222988 154018
rect 222936 153954 222988 153960
rect 222384 153944 222436 153950
rect 222384 153886 222436 153892
rect 222948 149954 222976 153954
rect 223592 149954 223620 159326
rect 224144 159118 224172 163200
rect 224972 159390 225000 163200
rect 225144 159520 225196 159526
rect 225144 159462 225196 159468
rect 224960 159384 225012 159390
rect 224960 159326 225012 159332
rect 224132 159112 224184 159118
rect 224132 159054 224184 159060
rect 224960 159044 225012 159050
rect 224960 158986 225012 158992
rect 223856 158772 223908 158778
rect 223856 158714 223908 158720
rect 223868 152318 223896 158714
rect 224132 156936 224184 156942
rect 224132 156878 224184 156884
rect 223856 152312 223908 152318
rect 223856 152254 223908 152260
rect 224144 149954 224172 156878
rect 224972 156874 225000 158986
rect 224960 156868 225012 156874
rect 224960 156810 225012 156816
rect 225052 156800 225104 156806
rect 225052 156742 225104 156748
rect 225064 149954 225092 156742
rect 225156 152998 225184 159462
rect 225512 156528 225564 156534
rect 225512 156470 225564 156476
rect 225144 152992 225196 152998
rect 225144 152934 225196 152940
rect 225524 149954 225552 156470
rect 225800 153950 225828 163200
rect 226628 156806 226656 163200
rect 226708 157412 226760 157418
rect 226708 157354 226760 157360
rect 226616 156800 226668 156806
rect 226616 156742 226668 156748
rect 225788 153944 225840 153950
rect 225788 153886 225840 153892
rect 226340 152652 226392 152658
rect 226340 152594 226392 152600
rect 226352 149954 226380 152594
rect 226720 149954 226748 157354
rect 227456 152425 227484 163200
rect 227996 156460 228048 156466
rect 227996 156402 228048 156408
rect 227812 155372 227864 155378
rect 227812 155314 227864 155320
rect 227442 152416 227498 152425
rect 227442 152351 227498 152360
rect 227824 150226 227852 155314
rect 227778 150198 227852 150226
rect 218440 149926 218776 149954
rect 218992 149926 219420 149954
rect 219728 149926 220064 149954
rect 220280 149926 220708 149954
rect 221016 149926 221352 149954
rect 221568 149926 221996 149954
rect 222212 149926 222640 149954
rect 222948 149926 223284 149954
rect 223592 149926 223928 149954
rect 224144 149926 224572 149954
rect 225064 149926 225216 149954
rect 225524 149926 225860 149954
rect 226352 149926 226504 149954
rect 226720 149926 227148 149954
rect 227778 149940 227806 150198
rect 228008 149954 228036 156402
rect 228284 152590 228312 163200
rect 229112 153746 229140 163200
rect 229284 157072 229336 157078
rect 229284 157014 229336 157020
rect 229100 153740 229152 153746
rect 229100 153682 229152 153688
rect 228732 152992 228784 152998
rect 228732 152934 228784 152940
rect 228824 152992 228876 152998
rect 228824 152934 228876 152940
rect 228272 152584 228324 152590
rect 228272 152526 228324 152532
rect 228744 149954 228772 152934
rect 228836 152726 228864 152934
rect 228824 152720 228876 152726
rect 228824 152662 228876 152668
rect 229296 149954 229324 157014
rect 230032 156738 230060 163200
rect 230860 159050 230888 163200
rect 231688 159526 231716 163200
rect 232516 161474 232544 163200
rect 232516 161446 232636 161474
rect 231676 159520 231728 159526
rect 231676 159462 231728 159468
rect 230848 159044 230900 159050
rect 230848 158986 230900 158992
rect 231032 158976 231084 158982
rect 231032 158918 231084 158924
rect 231044 157078 231072 158918
rect 231860 158092 231912 158098
rect 231860 158034 231912 158040
rect 231032 157072 231084 157078
rect 231032 157014 231084 157020
rect 230020 156732 230072 156738
rect 230020 156674 230072 156680
rect 230020 154964 230072 154970
rect 230020 154906 230072 154912
rect 230032 149954 230060 154906
rect 230664 153604 230716 153610
rect 230664 153546 230716 153552
rect 230676 149954 230704 153546
rect 231308 152788 231360 152794
rect 231308 152730 231360 152736
rect 231320 149954 231348 152730
rect 231872 149954 231900 158034
rect 232504 154828 232556 154834
rect 232504 154770 232556 154776
rect 232516 149954 232544 154770
rect 232608 153814 232636 161446
rect 233240 157004 233292 157010
rect 233240 156946 233292 156952
rect 232596 153808 232648 153814
rect 232596 153750 232648 153756
rect 233252 149954 233280 156946
rect 233344 155310 233372 163200
rect 234172 163146 234200 163200
rect 234264 163146 234292 163254
rect 234172 163118 234292 163146
rect 233792 159452 233844 159458
rect 233792 159394 233844 159400
rect 233332 155304 233384 155310
rect 233332 155246 233384 155252
rect 233804 149954 233832 159394
rect 234540 152658 234568 163254
rect 234986 163200 235042 164400
rect 235906 163200 235962 164400
rect 236734 163200 236790 164400
rect 237562 163200 237618 164400
rect 238390 163200 238446 164400
rect 239218 163200 239274 164400
rect 240046 163200 240102 164400
rect 240874 163200 240930 164400
rect 241794 163200 241850 164400
rect 242622 163200 242678 164400
rect 243450 163200 243506 164400
rect 244278 163200 244334 164400
rect 245106 163200 245162 164400
rect 245934 163200 245990 164400
rect 246762 163200 246818 164400
rect 247682 163200 247738 164400
rect 248510 163200 248566 164400
rect 249338 163200 249394 164400
rect 249444 163254 249748 163282
rect 235000 159458 235028 163200
rect 234988 159452 235040 159458
rect 234988 159394 235040 159400
rect 234620 157140 234672 157146
rect 234620 157082 234672 157088
rect 234528 152652 234580 152658
rect 234528 152594 234580 152600
rect 234632 149954 234660 157082
rect 235920 154086 235948 163200
rect 236748 158030 236776 163200
rect 237576 158982 237604 163200
rect 237564 158976 237616 158982
rect 237564 158918 237616 158924
rect 238404 158846 238432 163200
rect 238944 159588 238996 159594
rect 238944 159530 238996 159536
rect 238392 158840 238444 158846
rect 238392 158782 238444 158788
rect 237380 158160 237432 158166
rect 237380 158102 237432 158108
rect 236736 158024 236788 158030
rect 236736 157966 236788 157972
rect 236092 157684 236144 157690
rect 236092 157626 236144 157632
rect 235172 154080 235224 154086
rect 235172 154022 235224 154028
rect 235908 154080 235960 154086
rect 235908 154022 235960 154028
rect 235184 149954 235212 154022
rect 236104 150226 236132 157626
rect 236460 151836 236512 151842
rect 236460 151778 236512 151784
rect 236104 150198 236178 150226
rect 228008 149926 228436 149954
rect 228744 149926 229080 149954
rect 229296 149926 229724 149954
rect 230032 149926 230368 149954
rect 230676 149926 231012 149954
rect 231320 149926 231656 149954
rect 231872 149926 232300 149954
rect 232516 149926 232944 149954
rect 233252 149926 233588 149954
rect 233804 149926 234232 149954
rect 234632 149926 234876 149954
rect 235184 149926 235520 149954
rect 236150 149940 236178 150198
rect 236472 149954 236500 151778
rect 237392 150226 237420 158102
rect 237656 154760 237708 154766
rect 237656 154702 237708 154708
rect 237392 150198 237466 150226
rect 236472 149926 236808 149954
rect 237438 149940 237466 150198
rect 237668 149954 237696 154702
rect 238392 153672 238444 153678
rect 238392 153614 238444 153620
rect 238404 149954 238432 153614
rect 238956 149954 238984 159530
rect 239232 153678 239260 163200
rect 239680 158228 239732 158234
rect 239680 158170 239732 158176
rect 239220 153672 239272 153678
rect 239220 153614 239272 153620
rect 239692 149954 239720 158170
rect 240060 155242 240088 163200
rect 240888 158778 240916 163200
rect 241428 159656 241480 159662
rect 241428 159598 241480 159604
rect 240876 158772 240928 158778
rect 240876 158714 240928 158720
rect 240048 155236 240100 155242
rect 240048 155178 240100 155184
rect 240232 154624 240284 154630
rect 240232 154566 240284 154572
rect 240244 149954 240272 154566
rect 240968 154148 241020 154154
rect 240968 154090 241020 154096
rect 240980 149954 241008 154090
rect 241440 151814 241468 159598
rect 241808 159594 241836 163200
rect 241796 159588 241848 159594
rect 241796 159530 241848 159536
rect 242072 158296 242124 158302
rect 242072 158238 242124 158244
rect 241440 151786 241560 151814
rect 241532 149954 241560 151786
rect 242084 149954 242112 158238
rect 242636 154154 242664 163200
rect 242808 158840 242860 158846
rect 242808 158782 242860 158788
rect 242624 154148 242676 154154
rect 242624 154090 242676 154096
rect 242820 152114 242848 158782
rect 243360 158772 243412 158778
rect 243360 158714 243412 158720
rect 242900 154692 242952 154698
rect 242900 154634 242952 154640
rect 242808 152108 242860 152114
rect 242808 152050 242860 152056
rect 242912 149954 242940 154634
rect 243372 152046 243400 158714
rect 243464 158098 243492 163200
rect 244292 159662 244320 163200
rect 244280 159656 244332 159662
rect 244280 159598 244332 159604
rect 244648 158432 244700 158438
rect 244648 158374 244700 158380
rect 243452 158092 243504 158098
rect 243452 158034 243504 158040
rect 243452 153400 243504 153406
rect 243452 153342 243504 153348
rect 243360 152040 243412 152046
rect 243360 151982 243412 151988
rect 243464 149954 243492 153342
rect 244280 152856 244332 152862
rect 244280 152798 244332 152804
rect 244292 149954 244320 152798
rect 244660 149954 244688 158374
rect 245120 152794 245148 163200
rect 245948 161474 245976 163200
rect 245948 161446 246068 161474
rect 245936 154896 245988 154902
rect 245936 154838 245988 154844
rect 245660 154216 245712 154222
rect 245660 154158 245712 154164
rect 245108 152788 245160 152794
rect 245108 152730 245160 152736
rect 245672 150226 245700 154158
rect 245672 150198 245746 150226
rect 237668 149926 238096 149954
rect 238404 149926 238740 149954
rect 238956 149926 239384 149954
rect 239692 149926 240028 149954
rect 240244 149926 240672 149954
rect 240980 149926 241316 149954
rect 241532 149926 241960 149954
rect 242084 149926 242512 149954
rect 242912 149926 243156 149954
rect 243464 149926 243800 149954
rect 244292 149926 244444 149954
rect 244660 149926 245088 149954
rect 245718 149940 245746 150198
rect 245948 149954 245976 154838
rect 246040 153610 246068 161446
rect 246672 159724 246724 159730
rect 246672 159666 246724 159672
rect 246028 153604 246080 153610
rect 246028 153546 246080 153552
rect 246684 149954 246712 159666
rect 246776 158166 246804 163200
rect 247224 158364 247276 158370
rect 247224 158306 247276 158312
rect 246764 158160 246816 158166
rect 246764 158102 246816 158108
rect 247236 149954 247264 158306
rect 247696 152726 247724 163200
rect 248524 158914 248552 163200
rect 249352 163146 249380 163200
rect 249444 163146 249472 163254
rect 249352 163118 249472 163146
rect 248512 158908 248564 158914
rect 248512 158850 248564 158856
rect 247960 155508 248012 155514
rect 247960 155450 248012 155456
rect 247684 152720 247736 152726
rect 247684 152662 247736 152668
rect 247972 149954 248000 155450
rect 249720 154222 249748 163254
rect 250166 163200 250222 164400
rect 250994 163200 251050 164400
rect 251822 163200 251878 164400
rect 252650 163200 252706 164400
rect 253570 163200 253626 164400
rect 254398 163200 254454 164400
rect 255226 163200 255282 164400
rect 256054 163200 256110 164400
rect 256882 163200 256938 164400
rect 257710 163200 257766 164400
rect 258538 163200 258594 164400
rect 259458 163200 259514 164400
rect 260286 163200 260342 164400
rect 261114 163200 261170 164400
rect 261942 163200 261998 164400
rect 262770 163200 262826 164400
rect 263598 163200 263654 164400
rect 264426 163200 264482 164400
rect 265346 163200 265402 164400
rect 266174 163200 266230 164400
rect 267002 163200 267058 164400
rect 267830 163200 267886 164400
rect 268658 163200 268714 164400
rect 269486 163200 269542 164400
rect 270314 163200 270370 164400
rect 271234 163200 271290 164400
rect 272062 163200 272118 164400
rect 272168 163254 272656 163282
rect 249800 158500 249852 158506
rect 249800 158442 249852 158448
rect 249708 154216 249760 154222
rect 249708 154158 249760 154164
rect 248604 153468 248656 153474
rect 248604 153410 248656 153416
rect 248616 149954 248644 153410
rect 249248 153196 249300 153202
rect 249248 153138 249300 153144
rect 249260 149954 249288 153138
rect 249812 149954 249840 158442
rect 250180 154970 250208 163200
rect 251008 159730 251036 163200
rect 251836 161474 251864 163200
rect 251836 161446 251956 161474
rect 250996 159724 251048 159730
rect 250996 159666 251048 159672
rect 251272 157616 251324 157622
rect 251272 157558 251324 157564
rect 250168 154964 250220 154970
rect 250168 154906 250220 154912
rect 250536 154284 250588 154290
rect 250536 154226 250588 154232
rect 250548 149954 250576 154226
rect 251284 149954 251312 157558
rect 251824 153060 251876 153066
rect 251824 153002 251876 153008
rect 251836 149954 251864 153002
rect 251928 152862 251956 161446
rect 252560 158636 252612 158642
rect 252560 158578 252612 158584
rect 251916 152856 251968 152862
rect 251916 152798 251968 152804
rect 252572 149954 252600 158578
rect 252664 153474 252692 163200
rect 253020 155576 253072 155582
rect 253020 155518 253072 155524
rect 252652 153468 252704 153474
rect 252652 153410 252704 153416
rect 253032 149954 253060 155518
rect 253584 155378 253612 163200
rect 254308 159792 254360 159798
rect 254308 159734 254360 159740
rect 254032 157208 254084 157214
rect 254032 157150 254084 157156
rect 253572 155372 253624 155378
rect 253572 155314 253624 155320
rect 254044 150226 254072 157150
rect 254044 150198 254118 150226
rect 245948 149926 246376 149954
rect 246684 149926 247020 149954
rect 247236 149926 247664 149954
rect 247972 149926 248308 149954
rect 248616 149926 248952 149954
rect 249260 149926 249596 149954
rect 249812 149926 250240 149954
rect 250548 149926 250884 149954
rect 251284 149926 251528 149954
rect 251836 149926 252172 149954
rect 252572 149926 252816 149954
rect 253032 149926 253460 149954
rect 254090 149940 254118 150198
rect 254320 149954 254348 159734
rect 254412 158778 254440 163200
rect 255240 159798 255268 163200
rect 255228 159792 255280 159798
rect 255228 159734 255280 159740
rect 254400 158772 254452 158778
rect 254400 158714 254452 158720
rect 255320 158772 255372 158778
rect 255320 158714 255372 158720
rect 255332 153202 255360 158714
rect 255412 158568 255464 158574
rect 255412 158510 255464 158516
rect 255320 153196 255372 153202
rect 255320 153138 255372 153144
rect 255424 150226 255452 158510
rect 255596 155644 255648 155650
rect 255596 155586 255648 155592
rect 255378 150198 255452 150226
rect 254320 149926 254748 149954
rect 255378 149940 255406 150198
rect 255608 149954 255636 155586
rect 256068 154290 256096 163200
rect 256896 158234 256924 163200
rect 257528 158704 257580 158710
rect 257528 158646 257580 158652
rect 256884 158228 256936 158234
rect 256884 158170 256936 158176
rect 256332 157548 256384 157554
rect 256332 157490 256384 157496
rect 256056 154284 256108 154290
rect 256056 154226 256108 154232
rect 256344 149954 256372 157490
rect 256976 152380 257028 152386
rect 256976 152322 257028 152328
rect 256988 149954 257016 152322
rect 257540 149954 257568 158646
rect 257724 153066 257752 163200
rect 258552 158778 258580 163200
rect 258540 158772 258592 158778
rect 258540 158714 258592 158720
rect 258264 154420 258316 154426
rect 258264 154362 258316 154368
rect 257712 153060 257764 153066
rect 257712 153002 257764 153008
rect 258276 149954 258304 154362
rect 258908 153536 258960 153542
rect 258908 153478 258960 153484
rect 258920 149954 258948 153478
rect 259472 153406 259500 163200
rect 259644 159860 259696 159866
rect 259644 159802 259696 159808
rect 259460 153400 259512 153406
rect 259460 153342 259512 153348
rect 259656 149954 259684 159802
rect 260196 157956 260248 157962
rect 260196 157898 260248 157904
rect 260208 149954 260236 157898
rect 260300 155514 260328 163200
rect 261128 158846 261156 163200
rect 261956 159866 261984 163200
rect 261944 159860 261996 159866
rect 261944 159802 261996 159808
rect 261116 158840 261168 158846
rect 261116 158782 261168 158788
rect 260932 158772 260984 158778
rect 260932 158714 260984 158720
rect 260840 155712 260892 155718
rect 260840 155654 260892 155660
rect 260288 155508 260340 155514
rect 260288 155450 260340 155456
rect 260852 149954 260880 155654
rect 260944 152386 260972 158714
rect 262680 157888 262732 157894
rect 262680 157830 262732 157836
rect 261392 155440 261444 155446
rect 261392 155382 261444 155388
rect 260932 152380 260984 152386
rect 260932 152322 260984 152328
rect 261404 149954 261432 155382
rect 262220 152924 262272 152930
rect 262220 152866 262272 152872
rect 262232 149954 262260 152866
rect 262692 149954 262720 157830
rect 262784 153542 262812 163200
rect 263612 155582 263640 163200
rect 264440 158778 264468 163200
rect 264888 159928 264940 159934
rect 264888 159870 264940 159876
rect 264428 158772 264480 158778
rect 264428 158714 264480 158720
rect 264060 157752 264112 157758
rect 264060 157694 264112 157700
rect 263692 155848 263744 155854
rect 263692 155790 263744 155796
rect 263600 155576 263652 155582
rect 263600 155518 263652 155524
rect 262772 153536 262824 153542
rect 262772 153478 262824 153484
rect 263704 150226 263732 155790
rect 263704 150198 263778 150226
rect 255608 149926 256036 149954
rect 256344 149926 256680 149954
rect 256988 149926 257324 149954
rect 257540 149926 257968 149954
rect 258276 149926 258612 149954
rect 258920 149926 259256 149954
rect 259656 149926 259900 149954
rect 260208 149926 260544 149954
rect 260852 149926 261188 149954
rect 261404 149926 261832 149954
rect 262232 149926 262476 149954
rect 262692 149926 263120 149954
rect 263750 149940 263778 150198
rect 264072 149954 264100 157694
rect 264900 151814 264928 159870
rect 265164 157276 265216 157282
rect 265164 157218 265216 157224
rect 265176 151814 265204 157218
rect 265360 152930 265388 163200
rect 265900 155916 265952 155922
rect 265900 155858 265952 155864
rect 265348 152924 265400 152930
rect 265348 152866 265400 152872
rect 264900 151786 265020 151814
rect 265176 151786 265296 151814
rect 264992 150226 265020 151786
rect 264992 150198 265066 150226
rect 264072 149926 264408 149954
rect 265038 149940 265066 150198
rect 265268 149954 265296 151786
rect 265912 149954 265940 155858
rect 266188 154426 266216 163200
rect 266544 156188 266596 156194
rect 266544 156130 266596 156136
rect 266176 154420 266228 154426
rect 266176 154362 266228 154368
rect 266556 149954 266584 156130
rect 267016 155718 267044 163200
rect 267844 158778 267872 163200
rect 268672 159934 268700 163200
rect 268660 159928 268712 159934
rect 268660 159870 268712 159876
rect 267096 158772 267148 158778
rect 267096 158714 267148 158720
rect 267832 158772 267884 158778
rect 267832 158714 267884 158720
rect 267004 155712 267056 155718
rect 267004 155654 267056 155660
rect 267108 153134 267136 158714
rect 267740 157820 267792 157826
rect 267740 157762 267792 157768
rect 266912 153128 266964 153134
rect 266912 153070 266964 153076
rect 267096 153128 267148 153134
rect 267096 153070 267148 153076
rect 266924 151814 266952 153070
rect 267752 151814 267780 157762
rect 268476 155168 268528 155174
rect 268476 155110 268528 155116
rect 266924 151786 267228 151814
rect 267752 151786 267872 151814
rect 267200 149954 267228 151786
rect 267844 149954 267872 151786
rect 268488 149954 268516 155110
rect 269212 155032 269264 155038
rect 269212 154974 269264 154980
rect 269224 149954 269252 154974
rect 269500 153270 269528 163200
rect 269764 159996 269816 160002
rect 269764 159938 269816 159944
rect 269488 153264 269540 153270
rect 269488 153206 269540 153212
rect 269776 149954 269804 159938
rect 270328 155650 270356 163200
rect 271248 160002 271276 163200
rect 272076 163146 272104 163200
rect 272168 163146 272196 163254
rect 272076 163118 272196 163146
rect 271236 159996 271288 160002
rect 271236 159938 271288 159944
rect 272524 159996 272576 160002
rect 272524 159938 272576 159944
rect 271972 156868 272024 156874
rect 271972 156810 272024 156816
rect 270500 155984 270552 155990
rect 270500 155926 270552 155932
rect 270316 155644 270368 155650
rect 270316 155586 270368 155592
rect 270512 149954 270540 155926
rect 271052 155100 271104 155106
rect 271052 155042 271104 155048
rect 271064 149954 271092 155042
rect 271984 149954 272012 156810
rect 272536 151978 272564 159938
rect 272432 151972 272484 151978
rect 272432 151914 272484 151920
rect 272524 151972 272576 151978
rect 272524 151914 272576 151920
rect 272444 149954 272472 151914
rect 272628 151842 272656 163254
rect 272890 163200 272946 164400
rect 273718 163200 273774 164400
rect 274546 163200 274602 164400
rect 275374 163200 275430 164400
rect 276202 163200 276258 164400
rect 277122 163200 277178 164400
rect 277950 163200 278006 164400
rect 278778 163200 278834 164400
rect 279606 163200 279662 164400
rect 279712 163254 280016 163282
rect 272904 153338 272932 163200
rect 273732 156942 273760 163200
rect 274560 159497 274588 163200
rect 275388 160002 275416 163200
rect 275376 159996 275428 160002
rect 275376 159938 275428 159944
rect 274546 159488 274602 159497
rect 274546 159423 274602 159432
rect 274822 159352 274878 159361
rect 274822 159287 274878 159296
rect 273720 156936 273772 156942
rect 273720 156878 273772 156884
rect 273536 156120 273588 156126
rect 273536 156062 273588 156068
rect 273260 156052 273312 156058
rect 273260 155994 273312 156000
rect 272892 153332 272944 153338
rect 272892 153274 272944 153280
rect 272616 151836 272668 151842
rect 272616 151778 272668 151784
rect 273272 150226 273300 155994
rect 273272 150198 273346 150226
rect 265268 149926 265696 149954
rect 265912 149926 266340 149954
rect 266556 149926 266984 149954
rect 267200 149926 267628 149954
rect 267844 149926 268272 149954
rect 268488 149926 268916 149954
rect 269224 149926 269560 149954
rect 269776 149926 270204 149954
rect 270512 149926 270848 149954
rect 271064 149926 271492 149954
rect 271984 149926 272136 149954
rect 272444 149926 272780 149954
rect 273318 149940 273346 150198
rect 273548 149954 273576 156062
rect 274272 152176 274324 152182
rect 274272 152118 274324 152124
rect 274284 149954 274312 152118
rect 274836 149954 274864 159287
rect 276112 155780 276164 155786
rect 276112 155722 276164 155728
rect 275560 154352 275612 154358
rect 275560 154294 275612 154300
rect 275572 149954 275600 154294
rect 276124 149954 276152 155722
rect 276216 154358 276244 163200
rect 276848 157072 276900 157078
rect 276848 157014 276900 157020
rect 276204 154352 276256 154358
rect 276204 154294 276256 154300
rect 276860 149954 276888 157014
rect 277136 156874 277164 163200
rect 277124 156868 277176 156874
rect 277124 156810 277176 156816
rect 277492 152516 277544 152522
rect 277492 152458 277544 152464
rect 277504 149954 277532 152458
rect 277964 152182 277992 163200
rect 278136 154488 278188 154494
rect 278136 154430 278188 154436
rect 277952 152176 278004 152182
rect 277952 152118 278004 152124
rect 278148 149954 278176 154430
rect 278792 152522 278820 163200
rect 279620 163146 279648 163200
rect 279712 163146 279740 163254
rect 279620 163118 279740 163146
rect 278872 156392 278924 156398
rect 278872 156334 278924 156340
rect 278780 152516 278832 152522
rect 278780 152458 278832 152464
rect 278884 149954 278912 156334
rect 279988 154494 280016 163254
rect 280434 163200 280490 164400
rect 281262 163200 281318 164400
rect 282090 163200 282146 164400
rect 283010 163200 283066 164400
rect 283116 163254 283420 163282
rect 280344 160064 280396 160070
rect 280344 160006 280396 160012
rect 279976 154488 280028 154494
rect 279976 154430 280028 154436
rect 279608 152516 279660 152522
rect 279608 152458 279660 152464
rect 279424 152448 279476 152454
rect 279424 152390 279476 152396
rect 279436 149954 279464 152390
rect 279620 152182 279648 152458
rect 279608 152176 279660 152182
rect 279608 152118 279660 152124
rect 280356 150226 280384 160006
rect 280448 157078 280476 163200
rect 281276 160070 281304 163200
rect 281264 160064 281316 160070
rect 281264 160006 281316 160012
rect 282104 159322 282132 163200
rect 283024 163146 283052 163200
rect 283116 163146 283144 163254
rect 283024 163118 283144 163146
rect 282000 159316 282052 159322
rect 282000 159258 282052 159264
rect 282092 159316 282144 159322
rect 282092 159258 282144 159264
rect 281632 157344 281684 157350
rect 281632 157286 281684 157292
rect 280436 157072 280488 157078
rect 280436 157014 280488 157020
rect 280710 153776 280766 153785
rect 280710 153711 280766 153720
rect 280356 150198 280430 150226
rect 273548 149926 273976 149954
rect 274284 149926 274620 149954
rect 274836 149926 275264 149954
rect 275572 149926 275908 149954
rect 276124 149926 276552 149954
rect 276860 149926 277196 149954
rect 277504 149926 277840 149954
rect 278148 149926 278484 149954
rect 278884 149926 279128 149954
rect 279436 149926 279772 149954
rect 280402 149940 280430 150198
rect 280724 149954 280752 153711
rect 281644 150226 281672 157286
rect 281644 150198 281718 150226
rect 280724 149926 281060 149954
rect 281690 149940 281718 150198
rect 282012 149954 282040 159258
rect 283012 159180 283064 159186
rect 283012 159122 283064 159128
rect 282920 152244 282972 152250
rect 282920 152186 282972 152192
rect 282932 150226 282960 152186
rect 283024 151910 283052 159122
rect 283392 153882 283420 163254
rect 283838 163200 283894 164400
rect 284666 163200 284722 164400
rect 285494 163200 285550 164400
rect 286322 163200 286378 164400
rect 287150 163200 287206 164400
rect 287978 163200 288034 164400
rect 288898 163200 288954 164400
rect 289726 163200 289782 164400
rect 290554 163200 290610 164400
rect 291382 163200 291438 164400
rect 292210 163200 292266 164400
rect 293038 163200 293094 164400
rect 293866 163200 293922 164400
rect 294786 163200 294842 164400
rect 295614 163200 295670 164400
rect 296442 163200 296498 164400
rect 297270 163200 297326 164400
rect 298098 163200 298154 164400
rect 298926 163200 298982 164400
rect 299032 163254 299428 163282
rect 283852 157010 283880 163200
rect 284680 159186 284708 163200
rect 285128 159248 285180 159254
rect 285128 159190 285180 159196
rect 284668 159180 284720 159186
rect 284668 159122 284720 159128
rect 283840 157004 283892 157010
rect 283840 156946 283892 156952
rect 283472 156324 283524 156330
rect 283472 156266 283524 156272
rect 283288 153876 283340 153882
rect 283288 153818 283340 153824
rect 283380 153876 283432 153882
rect 283380 153818 283432 153824
rect 283012 151904 283064 151910
rect 283012 151846 283064 151852
rect 282932 150198 283006 150226
rect 282012 149926 282348 149954
rect 282978 149940 283006 150198
rect 283300 149954 283328 153818
rect 283484 151814 283512 156266
rect 284576 152992 284628 152998
rect 284576 152934 284628 152940
rect 283484 151786 283880 151814
rect 283852 149954 283880 151786
rect 284588 149954 284616 152934
rect 285140 149954 285168 159190
rect 285508 152998 285536 163200
rect 285772 159180 285824 159186
rect 285772 159122 285824 159128
rect 285680 156256 285732 156262
rect 285680 156198 285732 156204
rect 285496 152992 285548 152998
rect 285496 152934 285548 152940
rect 285692 150550 285720 156198
rect 285784 152250 285812 159122
rect 286336 154562 286364 163200
rect 287164 157146 287192 163200
rect 287992 159254 288020 163200
rect 287980 159248 288032 159254
rect 287980 159190 288032 159196
rect 288912 159186 288940 163200
rect 288348 159180 288400 159186
rect 288348 159122 288400 159128
rect 288900 159180 288952 159186
rect 288900 159122 288952 159128
rect 287152 157140 287204 157146
rect 287152 157082 287204 157088
rect 286232 154556 286284 154562
rect 286232 154498 286284 154504
rect 286324 154556 286376 154562
rect 286324 154498 286376 154504
rect 285772 152244 285824 152250
rect 285772 152186 285824 152192
rect 285680 150544 285732 150550
rect 285680 150486 285732 150492
rect 286244 150226 286272 154498
rect 288360 152318 288388 159122
rect 288992 156664 289044 156670
rect 288992 156606 289044 156612
rect 288440 154012 288492 154018
rect 288440 153954 288492 153960
rect 287796 152312 287848 152318
rect 287796 152254 287848 152260
rect 288348 152312 288400 152318
rect 288348 152254 288400 152260
rect 287152 151904 287204 151910
rect 287152 151846 287204 151852
rect 286508 150544 286560 150550
rect 286508 150486 286560 150492
rect 286198 150198 286272 150226
rect 283300 149926 283636 149954
rect 283852 149926 284280 149954
rect 284588 149926 284924 149954
rect 285140 149926 285568 149954
rect 286198 149940 286226 150198
rect 286520 149954 286548 150486
rect 287164 149954 287192 151846
rect 287808 149954 287836 152254
rect 288452 149954 288480 153954
rect 289004 149954 289032 156606
rect 289740 155786 289768 163200
rect 290280 159384 290332 159390
rect 290280 159326 290332 159332
rect 289728 155780 289780 155786
rect 289728 155722 289780 155728
rect 289912 152312 289964 152318
rect 289912 152254 289964 152260
rect 289924 149954 289952 152254
rect 290292 149954 290320 159326
rect 290568 157214 290596 163200
rect 290556 157208 290608 157214
rect 290556 157150 290608 157156
rect 291200 153944 291252 153950
rect 291200 153886 291252 153892
rect 291212 149954 291240 153886
rect 291396 152182 291424 163200
rect 291568 156800 291620 156806
rect 291568 156742 291620 156748
rect 291384 152176 291436 152182
rect 291384 152118 291436 152124
rect 291580 149954 291608 156742
rect 292224 152318 292252 163200
rect 293052 155922 293080 163200
rect 293880 156670 293908 163200
rect 294800 159390 294828 163200
rect 295628 159526 295656 163200
rect 295524 159520 295576 159526
rect 295524 159462 295576 159468
rect 295616 159520 295668 159526
rect 295616 159462 295668 159468
rect 294788 159384 294840 159390
rect 294788 159326 294840 159332
rect 294788 159044 294840 159050
rect 294788 158986 294840 158992
rect 294052 156732 294104 156738
rect 294052 156674 294104 156680
rect 293868 156664 293920 156670
rect 293868 156606 293920 156612
rect 293040 155916 293092 155922
rect 293040 155858 293092 155864
rect 293592 153740 293644 153746
rect 293592 153682 293644 153688
rect 292948 152584 293000 152590
rect 292948 152526 293000 152532
rect 292578 152416 292634 152425
rect 292578 152351 292634 152360
rect 292212 152312 292264 152318
rect 292212 152254 292264 152260
rect 292592 150226 292620 152351
rect 292592 150198 292666 150226
rect 286520 149926 286856 149954
rect 287164 149926 287500 149954
rect 287808 149926 288144 149954
rect 288452 149926 288788 149954
rect 289004 149926 289432 149954
rect 289924 149926 290076 149954
rect 290292 149926 290720 149954
rect 291212 149926 291364 149954
rect 291580 149926 292008 149954
rect 292638 149940 292666 150198
rect 292960 149954 292988 152526
rect 293604 149954 293632 153682
rect 294064 151814 294092 156674
rect 294064 151786 294184 151814
rect 294156 149954 294184 151786
rect 294800 149954 294828 158986
rect 295536 149954 295564 159462
rect 296456 155854 296484 163200
rect 297284 156806 297312 163200
rect 297824 159656 297876 159662
rect 297824 159598 297876 159604
rect 297836 159118 297864 159598
rect 298008 159452 298060 159458
rect 298008 159394 298060 159400
rect 297824 159112 297876 159118
rect 297824 159054 297876 159060
rect 297272 156800 297324 156806
rect 297272 156742 297324 156748
rect 296444 155848 296496 155854
rect 296444 155790 296496 155796
rect 296812 155304 296864 155310
rect 296812 155246 296864 155252
rect 296168 153808 296220 153814
rect 296168 153750 296220 153756
rect 296180 149954 296208 153750
rect 296824 149954 296852 155246
rect 297456 152652 297508 152658
rect 297456 152594 297508 152600
rect 297468 149954 297496 152594
rect 298020 151814 298048 159394
rect 298112 159050 298140 163200
rect 298940 163146 298968 163200
rect 299032 163146 299060 163254
rect 298940 163118 299060 163146
rect 298100 159044 298152 159050
rect 298100 158986 298152 158992
rect 298744 154080 298796 154086
rect 298744 154022 298796 154028
rect 298020 151786 298140 151814
rect 298112 149954 298140 151786
rect 298756 149954 298784 154022
rect 299400 152590 299428 163254
rect 299754 163200 299810 164400
rect 300674 163200 300730 164400
rect 301502 163200 301558 164400
rect 302330 163200 302386 164400
rect 303158 163200 303214 164400
rect 303986 163200 304042 164400
rect 304814 163200 304870 164400
rect 305642 163200 305698 164400
rect 306562 163200 306618 164400
rect 307390 163200 307446 164400
rect 308218 163200 308274 164400
rect 309046 163200 309102 164400
rect 309874 163200 309930 164400
rect 310702 163200 310758 164400
rect 311530 163200 311586 164400
rect 311636 163254 311848 163282
rect 299572 158024 299624 158030
rect 299572 157966 299624 157972
rect 299388 152584 299440 152590
rect 299388 152526 299440 152532
rect 299584 149954 299612 157966
rect 299768 155310 299796 163200
rect 299940 159044 299992 159050
rect 299940 158986 299992 158992
rect 299756 155304 299808 155310
rect 299756 155246 299808 155252
rect 299952 151910 299980 158986
rect 300032 158976 300084 158982
rect 300032 158918 300084 158924
rect 299940 151904 299992 151910
rect 299940 151846 299992 151852
rect 300044 149954 300072 158918
rect 300688 156738 300716 163200
rect 301516 159458 301544 163200
rect 302344 159594 302372 163200
rect 303068 159656 303120 159662
rect 303068 159598 303120 159604
rect 302332 159588 302384 159594
rect 302332 159530 302384 159536
rect 301504 159452 301556 159458
rect 301504 159394 301556 159400
rect 300676 156732 300728 156738
rect 300676 156674 300728 156680
rect 302332 155236 302384 155242
rect 302332 155178 302384 155184
rect 301320 153672 301372 153678
rect 301320 153614 301372 153620
rect 300860 152108 300912 152114
rect 300860 152050 300912 152056
rect 300872 149954 300900 152050
rect 301332 149954 301360 153614
rect 302344 150226 302372 155178
rect 302608 152040 302660 152046
rect 302608 151982 302660 151988
rect 302298 150198 302372 150226
rect 292960 149926 293296 149954
rect 293604 149926 293940 149954
rect 294156 149926 294584 149954
rect 294800 149926 295228 149954
rect 295536 149926 295872 149954
rect 296180 149926 296516 149954
rect 296824 149926 297160 149954
rect 297468 149926 297804 149954
rect 298112 149926 298448 149954
rect 298756 149926 299092 149954
rect 299584 149926 299736 149954
rect 300044 149926 300380 149954
rect 300872 149926 301024 149954
rect 301332 149926 301668 149954
rect 302298 149940 302326 150198
rect 302620 149954 302648 151982
rect 303080 151814 303108 159598
rect 303172 155242 303200 163200
rect 303160 155236 303212 155242
rect 303160 155178 303212 155184
rect 303804 154148 303856 154154
rect 303804 154090 303856 154096
rect 303080 151786 303200 151814
rect 303172 149954 303200 151786
rect 303816 149954 303844 154090
rect 304000 152114 304028 163200
rect 304356 158092 304408 158098
rect 304356 158034 304408 158040
rect 303988 152108 304040 152114
rect 303988 152050 304040 152056
rect 304368 149954 304396 158034
rect 304828 152658 304856 163200
rect 305184 159112 305236 159118
rect 305184 159054 305236 159060
rect 304816 152652 304868 152658
rect 304816 152594 304868 152600
rect 305196 149954 305224 159054
rect 305656 158914 305684 163200
rect 305644 158908 305696 158914
rect 305644 158850 305696 158856
rect 306576 155174 306604 163200
rect 307404 159118 307432 163200
rect 307392 159112 307444 159118
rect 307392 159054 307444 159060
rect 308232 159050 308260 163200
rect 309060 159662 309088 163200
rect 309048 159656 309100 159662
rect 309048 159598 309100 159604
rect 308220 159044 308272 159050
rect 308220 158986 308272 158992
rect 307668 158908 307720 158914
rect 307668 158850 307720 158856
rect 308220 158908 308272 158914
rect 308220 158850 308272 158856
rect 306932 158160 306984 158166
rect 306932 158102 306984 158108
rect 306564 155168 306616 155174
rect 306564 155110 306616 155116
rect 306380 153604 306432 153610
rect 306380 153546 306432 153552
rect 305736 152788 305788 152794
rect 305736 152730 305788 152736
rect 305748 149954 305776 152730
rect 306392 149954 306420 153546
rect 306944 149954 306972 158102
rect 307680 152794 307708 158850
rect 307668 152788 307720 152794
rect 307668 152730 307720 152736
rect 307760 152720 307812 152726
rect 307760 152662 307812 152668
rect 307772 149954 307800 152662
rect 308232 149954 308260 158850
rect 309508 154964 309560 154970
rect 309508 154906 309560 154912
rect 309232 154216 309284 154222
rect 309232 154158 309284 154164
rect 309244 150226 309272 154158
rect 309244 150198 309318 150226
rect 302620 149926 302956 149954
rect 303172 149926 303600 149954
rect 303816 149926 304152 149954
rect 304368 149926 304796 149954
rect 305196 149926 305440 149954
rect 305748 149926 306084 149954
rect 306392 149926 306728 149954
rect 306944 149926 307372 149954
rect 307772 149926 308016 149954
rect 308232 149926 308660 149954
rect 309290 149940 309318 150198
rect 309520 149954 309548 154906
rect 309888 153950 309916 163200
rect 310612 159724 310664 159730
rect 310612 159666 310664 159672
rect 309876 153944 309928 153950
rect 309876 153886 309928 153892
rect 310624 150226 310652 159666
rect 310716 158914 310744 163200
rect 311544 163146 311572 163200
rect 311636 163146 311664 163254
rect 311544 163118 311664 163146
rect 310704 158908 310756 158914
rect 310704 158850 310756 158856
rect 311532 153468 311584 153474
rect 311532 153410 311584 153416
rect 310888 152856 310940 152862
rect 310888 152798 310940 152804
rect 310578 150198 310652 150226
rect 309520 149926 309948 149954
rect 310578 149940 310606 150198
rect 310900 149954 310928 152798
rect 311544 149954 311572 153410
rect 311820 152726 311848 163254
rect 312450 163200 312506 164400
rect 313278 163200 313334 164400
rect 314106 163200 314162 164400
rect 314934 163200 314990 164400
rect 315762 163200 315818 164400
rect 316590 163200 316646 164400
rect 317418 163200 317474 164400
rect 318338 163200 318394 164400
rect 318444 163254 318656 163282
rect 312464 158914 312492 163200
rect 311992 158908 312044 158914
rect 311992 158850 312044 158856
rect 312452 158908 312504 158914
rect 312452 158850 312504 158856
rect 312004 152862 312032 158850
rect 312084 155372 312136 155378
rect 312084 155314 312136 155320
rect 311992 152856 312044 152862
rect 311992 152798 312044 152804
rect 311808 152720 311860 152726
rect 311808 152662 311860 152668
rect 312096 149954 312124 155314
rect 313292 154018 313320 163200
rect 314120 159798 314148 163200
rect 313372 159792 313424 159798
rect 313372 159734 313424 159740
rect 314108 159792 314160 159798
rect 314108 159734 314160 159740
rect 313280 154012 313332 154018
rect 313280 153954 313332 153960
rect 312820 153196 312872 153202
rect 312820 153138 312872 153144
rect 312832 149954 312860 153138
rect 313384 149954 313412 159734
rect 314948 158982 314976 163200
rect 315776 159730 315804 163200
rect 315764 159724 315816 159730
rect 315764 159666 315816 159672
rect 314936 158976 314988 158982
rect 314936 158918 314988 158924
rect 313464 158908 313516 158914
rect 313464 158850 313516 158856
rect 313476 152425 313504 158850
rect 314752 158228 314804 158234
rect 314752 158170 314804 158176
rect 314108 154284 314160 154290
rect 314108 154226 314160 154232
rect 313462 152416 313518 152425
rect 313462 152351 313518 152360
rect 314120 149954 314148 154226
rect 314764 149954 314792 158170
rect 316604 154086 316632 163200
rect 316960 158840 317012 158846
rect 316960 158782 317012 158788
rect 316592 154080 316644 154086
rect 316592 154022 316644 154028
rect 316776 153400 316828 153406
rect 316776 153342 316828 153348
rect 315396 153060 315448 153066
rect 315396 153002 315448 153008
rect 315408 149954 315436 153002
rect 316040 152380 316092 152386
rect 316040 152322 316092 152328
rect 316052 149954 316080 152322
rect 316788 149954 316816 153342
rect 316972 153202 317000 158782
rect 316960 153196 317012 153202
rect 316960 153138 317012 153144
rect 317432 153066 317460 163200
rect 318352 163146 318380 163200
rect 318444 163146 318472 163254
rect 318352 163118 318472 163146
rect 317512 155508 317564 155514
rect 317512 155450 317564 155456
rect 317420 153060 317472 153066
rect 317420 153002 317472 153008
rect 317524 149954 317552 155450
rect 318628 153202 318656 163254
rect 319166 163200 319222 164400
rect 319994 163200 320050 164400
rect 320822 163200 320878 164400
rect 321650 163200 321706 164400
rect 322478 163200 322534 164400
rect 323306 163200 323362 164400
rect 324226 163200 324282 164400
rect 325054 163200 325110 164400
rect 325882 163200 325938 164400
rect 326710 163200 326766 164400
rect 327538 163200 327594 164400
rect 328366 163200 328422 164400
rect 329194 163200 329250 164400
rect 330114 163200 330170 164400
rect 330942 163200 330998 164400
rect 331770 163200 331826 164400
rect 332598 163200 332654 164400
rect 333426 163200 333482 164400
rect 334254 163200 334310 164400
rect 335082 163200 335138 164400
rect 336002 163200 336058 164400
rect 336830 163200 336886 164400
rect 337658 163200 337714 164400
rect 338486 163200 338542 164400
rect 339314 163200 339370 164400
rect 340142 163200 340198 164400
rect 340970 163200 341026 164400
rect 341890 163200 341946 164400
rect 342718 163200 342774 164400
rect 343546 163200 343602 164400
rect 344374 163200 344430 164400
rect 345202 163200 345258 164400
rect 346030 163200 346086 164400
rect 346858 163200 346914 164400
rect 347778 163200 347834 164400
rect 348606 163200 348662 164400
rect 348712 163254 349108 163282
rect 318984 159860 319036 159866
rect 318984 159802 319036 159808
rect 317972 153196 318024 153202
rect 317972 153138 318024 153144
rect 318616 153196 318668 153202
rect 318616 153138 318668 153144
rect 317984 149954 318012 153138
rect 318996 150226 319024 159802
rect 319180 158914 319208 163200
rect 319168 158908 319220 158914
rect 319168 158850 319220 158856
rect 320008 155378 320036 163200
rect 320836 159866 320864 163200
rect 320824 159860 320876 159866
rect 320824 159802 320876 159808
rect 321664 158778 321692 163200
rect 322492 158846 322520 163200
rect 322848 158908 322900 158914
rect 322848 158850 322900 158856
rect 322480 158840 322532 158846
rect 322480 158782 322532 158788
rect 320272 158772 320324 158778
rect 320272 158714 320324 158720
rect 321652 158772 321704 158778
rect 321652 158714 321704 158720
rect 320180 155576 320232 155582
rect 320180 155518 320232 155524
rect 319996 155372 320048 155378
rect 319996 155314 320048 155320
rect 319260 153536 319312 153542
rect 319260 153478 319312 153484
rect 318950 150198 319024 150226
rect 310900 149926 311236 149954
rect 311544 149926 311880 149954
rect 312096 149926 312524 149954
rect 312832 149926 313168 149954
rect 313384 149926 313812 149954
rect 314120 149926 314456 149954
rect 314764 149926 315100 149954
rect 315408 149926 315744 149954
rect 316052 149926 316388 149954
rect 316788 149926 317032 149954
rect 317524 149926 317676 149954
rect 317984 149926 318320 149954
rect 318950 149940 318978 150198
rect 319272 149954 319300 153478
rect 320192 150226 320220 155518
rect 320284 152386 320312 158714
rect 322112 155712 322164 155718
rect 322112 155654 322164 155660
rect 321836 154420 321888 154426
rect 321836 154362 321888 154368
rect 320640 153196 320692 153202
rect 320640 153138 320692 153144
rect 320456 153128 320508 153134
rect 320456 153070 320508 153076
rect 320272 152380 320324 152386
rect 320272 152322 320324 152328
rect 320192 150198 320266 150226
rect 319272 149926 319608 149954
rect 320238 149940 320266 150198
rect 320468 149954 320496 153070
rect 320652 153066 320680 153138
rect 320640 153060 320692 153066
rect 320640 153002 320692 153008
rect 321192 152924 321244 152930
rect 321192 152866 321244 152872
rect 321204 149954 321232 152866
rect 321848 149954 321876 154362
rect 322124 151814 322152 155654
rect 322860 152538 322888 158850
rect 323320 154154 323348 163200
rect 323676 159928 323728 159934
rect 323676 159870 323728 159876
rect 323308 154148 323360 154154
rect 323308 154090 323360 154096
rect 322860 152510 323256 152538
rect 323228 152386 323256 152510
rect 323124 152380 323176 152386
rect 323124 152322 323176 152328
rect 323216 152380 323268 152386
rect 323216 152322 323268 152328
rect 322124 151786 322428 151814
rect 322400 149954 322428 151786
rect 323136 149954 323164 152322
rect 323688 149954 323716 159870
rect 324240 152930 324268 163200
rect 324964 155644 325016 155650
rect 324964 155586 325016 155592
rect 324412 153264 324464 153270
rect 324412 153206 324464 153212
rect 324228 152924 324280 152930
rect 324228 152866 324280 152872
rect 324424 149954 324452 153206
rect 324976 149954 325004 155586
rect 325068 153134 325096 163200
rect 325056 153128 325108 153134
rect 325056 153070 325108 153076
rect 325700 152040 325752 152046
rect 325700 151982 325752 151988
rect 325712 149954 325740 151982
rect 325896 151978 325924 163200
rect 326724 154222 326752 163200
rect 327448 160064 327500 160070
rect 327448 160006 327500 160012
rect 327460 159322 327488 160006
rect 327552 159322 327580 163200
rect 328380 159934 328408 163200
rect 329208 160002 329236 163200
rect 328828 159996 328880 160002
rect 328828 159938 328880 159944
rect 329196 159996 329248 160002
rect 329196 159938 329248 159944
rect 328368 159928 328420 159934
rect 328368 159870 328420 159876
rect 328458 159488 328514 159497
rect 328458 159423 328514 159432
rect 327448 159316 327500 159322
rect 327448 159258 327500 159264
rect 327540 159316 327592 159322
rect 327540 159258 327592 159264
rect 327540 156936 327592 156942
rect 327540 156878 327592 156884
rect 326712 154216 326764 154222
rect 326712 154158 326764 154164
rect 327080 153332 327132 153338
rect 327080 153274 327132 153280
rect 325884 151972 325936 151978
rect 325884 151914 325936 151920
rect 326344 151836 326396 151842
rect 326344 151778 326396 151784
rect 326356 149954 326384 151778
rect 327092 149954 327120 153274
rect 327552 149954 327580 156878
rect 328472 149954 328500 159423
rect 328840 149954 328868 159938
rect 330024 156868 330076 156874
rect 330024 156810 330076 156816
rect 329840 154352 329892 154358
rect 329840 154294 329892 154300
rect 329852 150226 329880 154294
rect 330036 151814 330064 156810
rect 330128 155446 330156 163200
rect 330668 160132 330720 160138
rect 330668 160074 330720 160080
rect 330680 159322 330708 160074
rect 330576 159316 330628 159322
rect 330576 159258 330628 159264
rect 330668 159316 330720 159322
rect 330668 159258 330720 159264
rect 330588 158778 330616 159258
rect 330576 158772 330628 158778
rect 330576 158714 330628 158720
rect 330116 155440 330168 155446
rect 330116 155382 330168 155388
rect 330956 152522 330984 163200
rect 330852 152516 330904 152522
rect 330852 152458 330904 152464
rect 330944 152516 330996 152522
rect 330944 152458 330996 152464
rect 330484 152380 330536 152386
rect 330484 152322 330536 152328
rect 330576 152380 330628 152386
rect 330576 152322 330628 152328
rect 330496 152046 330524 152322
rect 330484 152040 330536 152046
rect 330484 151982 330536 151988
rect 330588 151978 330616 152322
rect 330576 151972 330628 151978
rect 330576 151914 330628 151920
rect 330036 151786 330156 151814
rect 329852 150198 329926 150226
rect 320468 149926 320896 149954
rect 321204 149926 321540 149954
rect 321848 149926 322184 149954
rect 322400 149926 322828 149954
rect 323136 149926 323472 149954
rect 323688 149926 324116 149954
rect 324424 149926 324760 149954
rect 324976 149926 325404 149954
rect 325712 149926 326048 149954
rect 326356 149926 326692 149954
rect 327092 149926 327336 149954
rect 327552 149926 327980 149954
rect 328472 149926 328624 149954
rect 328840 149926 329268 149954
rect 329898 149940 329926 150198
rect 330128 149954 330156 151786
rect 330864 149954 330892 152458
rect 331496 152448 331548 152454
rect 331496 152390 331548 152396
rect 331508 149954 331536 152390
rect 331784 151978 331812 163200
rect 332140 154488 332192 154494
rect 332140 154430 332192 154436
rect 331772 151972 331824 151978
rect 331772 151914 331824 151920
rect 332152 149954 332180 154430
rect 332612 152454 332640 163200
rect 333336 159316 333388 159322
rect 333336 159258 333388 159264
rect 332692 157072 332744 157078
rect 332692 157014 332744 157020
rect 332600 152448 332652 152454
rect 332600 152390 332652 152396
rect 332704 149954 332732 157014
rect 333348 149954 333376 159258
rect 333440 155514 333468 163200
rect 334268 160070 334296 163200
rect 335096 160070 335124 163200
rect 333980 160064 334032 160070
rect 333980 160006 334032 160012
rect 334256 160064 334308 160070
rect 334256 160006 334308 160012
rect 335084 160064 335136 160070
rect 335084 160006 335136 160012
rect 333520 159316 333572 159322
rect 333520 159258 333572 159264
rect 333532 159186 333560 159258
rect 333520 159180 333572 159186
rect 333520 159122 333572 159128
rect 333428 155508 333480 155514
rect 333428 155450 333480 155456
rect 333992 149954 334020 160006
rect 335912 159520 335964 159526
rect 335912 159462 335964 159468
rect 335924 159254 335952 159462
rect 335912 159248 335964 159254
rect 335912 159190 335964 159196
rect 335452 157004 335504 157010
rect 335452 156946 335504 156952
rect 334624 153876 334676 153882
rect 334624 153818 334676 153824
rect 334636 149954 334664 153818
rect 335464 149954 335492 156946
rect 335912 152244 335964 152250
rect 335912 152186 335964 152192
rect 335924 149954 335952 152186
rect 336016 151842 336044 163200
rect 336096 160132 336148 160138
rect 336096 160074 336148 160080
rect 336108 159526 336136 160074
rect 336096 159520 336148 159526
rect 336096 159462 336148 159468
rect 336844 153882 336872 163200
rect 337672 155582 337700 163200
rect 338500 160070 338528 163200
rect 338488 160064 338540 160070
rect 338488 160006 338540 160012
rect 339328 159526 339356 163200
rect 339500 160064 339552 160070
rect 339500 160006 339552 160012
rect 339132 159520 339184 159526
rect 339132 159462 339184 159468
rect 339316 159520 339368 159526
rect 339316 159462 339368 159468
rect 339144 159322 339172 159462
rect 339040 159316 339092 159322
rect 339040 159258 339092 159264
rect 339132 159316 339184 159322
rect 339132 159258 339184 159264
rect 338396 159180 338448 159186
rect 338396 159122 338448 159128
rect 338120 157140 338172 157146
rect 338120 157082 338172 157088
rect 337660 155576 337712 155582
rect 337660 155518 337712 155524
rect 337200 154556 337252 154562
rect 337200 154498 337252 154504
rect 336832 153876 336884 153882
rect 336832 153818 336884 153824
rect 336740 152992 336792 152998
rect 336740 152934 336792 152940
rect 336004 151836 336056 151842
rect 336004 151778 336056 151784
rect 336752 149954 336780 152934
rect 337212 149954 337240 154498
rect 338132 150226 338160 157082
rect 338132 150198 338206 150226
rect 330128 149926 330556 149954
rect 330864 149926 331200 149954
rect 331508 149926 331844 149954
rect 332152 149926 332488 149954
rect 332704 149926 333132 149954
rect 333348 149926 333776 149954
rect 333992 149926 334420 149954
rect 334636 149926 334972 149954
rect 335464 149926 335616 149954
rect 335924 149926 336260 149954
rect 336752 149926 336904 149954
rect 337212 149926 337548 149954
rect 338178 149940 338206 150198
rect 338408 149954 338436 159122
rect 339052 149954 339080 159258
rect 339512 152998 339540 160006
rect 339960 157208 340012 157214
rect 339960 157150 340012 157156
rect 339592 155780 339644 155786
rect 339592 155722 339644 155728
rect 339500 152992 339552 152998
rect 339500 152934 339552 152940
rect 339604 151814 339632 155722
rect 339972 151814 340000 157150
rect 340156 154358 340184 163200
rect 340984 155718 341012 163200
rect 341904 159186 341932 163200
rect 342732 159254 342760 163200
rect 343456 159384 343508 159390
rect 343456 159326 343508 159332
rect 342444 159248 342496 159254
rect 342444 159190 342496 159196
rect 342720 159248 342772 159254
rect 342720 159190 342772 159196
rect 341892 159180 341944 159186
rect 341892 159122 341944 159128
rect 342260 156664 342312 156670
rect 342260 156606 342312 156612
rect 340972 155712 341024 155718
rect 340972 155654 341024 155660
rect 340144 154352 340196 154358
rect 340144 154294 340196 154300
rect 341708 152312 341760 152318
rect 341708 152254 341760 152260
rect 341064 152244 341116 152250
rect 341064 152186 341116 152192
rect 341156 152244 341208 152250
rect 341156 152186 341208 152192
rect 340144 152176 340196 152182
rect 340144 152118 340196 152124
rect 340156 151910 340184 152118
rect 340144 151904 340196 151910
rect 340144 151846 340196 151852
rect 339604 151786 339724 151814
rect 339972 151786 340368 151814
rect 339696 149954 339724 151786
rect 340340 149954 340368 151786
rect 341076 149954 341104 152186
rect 341168 151842 341196 152186
rect 341156 151836 341208 151842
rect 341156 151778 341208 151784
rect 341720 149954 341748 152254
rect 342272 150550 342300 156606
rect 342352 155916 342404 155922
rect 342352 155858 342404 155864
rect 342260 150544 342312 150550
rect 342260 150486 342312 150492
rect 342364 149954 342392 155858
rect 342456 152318 342484 159190
rect 342444 152312 342496 152318
rect 342444 152254 342496 152260
rect 343468 151814 343496 159326
rect 343560 154290 343588 163200
rect 343824 159248 343876 159254
rect 343824 159190 343876 159196
rect 343548 154284 343600 154290
rect 343548 154226 343600 154232
rect 343836 151842 343864 159190
rect 344388 155650 344416 163200
rect 345112 155848 345164 155854
rect 345112 155790 345164 155796
rect 344376 155644 344428 155650
rect 344376 155586 344428 155592
rect 344284 152312 344336 152318
rect 344284 152254 344336 152260
rect 343824 151836 343876 151842
rect 343468 151786 343680 151814
rect 342996 150544 343048 150550
rect 342996 150486 343048 150492
rect 343008 149954 343036 150486
rect 343652 149954 343680 151786
rect 343824 151778 343876 151784
rect 344296 149954 344324 152254
rect 345124 149954 345152 155790
rect 345216 152318 345244 163200
rect 346044 159390 346072 163200
rect 346032 159384 346084 159390
rect 346032 159326 346084 159332
rect 345572 156800 345624 156806
rect 345572 156742 345624 156748
rect 345204 152312 345256 152318
rect 345204 152254 345256 152260
rect 345584 149954 345612 156742
rect 346872 154426 346900 163200
rect 347792 159594 347820 163200
rect 348620 163146 348648 163200
rect 348712 163146 348740 163254
rect 348620 163118 348740 163146
rect 347136 159588 347188 159594
rect 347136 159530 347188 159536
rect 347780 159588 347832 159594
rect 347780 159530 347832 159536
rect 347148 159254 347176 159530
rect 348792 159452 348844 159458
rect 348792 159394 348844 159400
rect 348976 159452 349028 159458
rect 348976 159394 349028 159400
rect 347136 159248 347188 159254
rect 347136 159190 347188 159196
rect 348056 156732 348108 156738
rect 348056 156674 348108 156680
rect 347780 155304 347832 155310
rect 347780 155246 347832 155252
rect 346860 154420 346912 154426
rect 346860 154362 346912 154368
rect 346860 152584 346912 152590
rect 346860 152526 346912 152532
rect 346400 152176 346452 152182
rect 346400 152118 346452 152124
rect 346412 149954 346440 152118
rect 346872 149954 346900 152526
rect 347792 150226 347820 155246
rect 347792 150198 347866 150226
rect 338408 149926 338836 149954
rect 339052 149926 339480 149954
rect 339696 149926 340124 149954
rect 340340 149926 340768 149954
rect 341076 149926 341412 149954
rect 341720 149926 342056 149954
rect 342364 149926 342700 149954
rect 343008 149926 343344 149954
rect 343652 149926 343988 149954
rect 344296 149926 344632 149954
rect 345124 149926 345276 149954
rect 345584 149926 345920 149954
rect 346412 149926 346564 149954
rect 346872 149926 347208 149954
rect 347838 149940 347866 150198
rect 348068 149954 348096 156674
rect 348804 149954 348832 159394
rect 348988 159050 349016 159394
rect 348976 159044 349028 159050
rect 348976 158986 349028 158992
rect 349080 152590 349108 163254
rect 349434 163200 349490 164400
rect 350262 163200 350318 164400
rect 351090 163200 351146 164400
rect 351918 163200 351974 164400
rect 352746 163200 352802 164400
rect 353666 163200 353722 164400
rect 354494 163200 354550 164400
rect 355322 163200 355378 164400
rect 356150 163200 356206 164400
rect 356978 163200 357034 164400
rect 357084 163254 357388 163282
rect 349344 159248 349396 159254
rect 349344 159190 349396 159196
rect 349068 152584 349120 152590
rect 349068 152526 349120 152532
rect 349356 149954 349384 159190
rect 349448 151910 349476 163200
rect 349804 159520 349856 159526
rect 349804 159462 349856 159468
rect 349816 159254 349844 159462
rect 349804 159248 349856 159254
rect 349804 159190 349856 159196
rect 350080 155236 350132 155242
rect 350080 155178 350132 155184
rect 349804 152176 349856 152182
rect 349804 152118 349856 152124
rect 349436 151904 349488 151910
rect 349436 151846 349488 151852
rect 349816 151842 349844 152118
rect 349804 151836 349856 151842
rect 349804 151778 349856 151784
rect 350092 149954 350120 155178
rect 350276 154494 350304 163200
rect 351104 159118 351132 163200
rect 351932 159594 351960 163200
rect 351920 159588 351972 159594
rect 351920 159530 351972 159536
rect 351092 159112 351144 159118
rect 351092 159054 351144 159060
rect 352472 155168 352524 155174
rect 352472 155110 352524 155116
rect 350264 154488 350316 154494
rect 350264 154430 350316 154436
rect 352012 152788 352064 152794
rect 352012 152730 352064 152736
rect 351368 152652 351420 152658
rect 351368 152594 351420 152600
rect 350724 152108 350776 152114
rect 350724 152050 350776 152056
rect 350736 149954 350764 152050
rect 351380 149954 351408 152594
rect 352024 149954 352052 152730
rect 352484 151814 352512 155110
rect 352760 152794 352788 163200
rect 353208 159044 353260 159050
rect 353208 158986 353260 158992
rect 352748 152788 352800 152794
rect 352748 152730 352800 152736
rect 353220 151814 353248 158986
rect 353680 154562 353708 163200
rect 353852 159452 353904 159458
rect 353852 159394 353904 159400
rect 353668 154556 353720 154562
rect 353668 154498 353720 154504
rect 352484 151786 352604 151814
rect 353220 151786 353340 151814
rect 352576 149954 352604 151786
rect 353312 149954 353340 151786
rect 353864 149954 353892 159394
rect 354508 152658 354536 163200
rect 354864 159656 354916 159662
rect 354864 159598 354916 159604
rect 354496 152652 354548 152658
rect 354496 152594 354548 152600
rect 354876 150226 354904 159598
rect 355232 153944 355284 153950
rect 355232 153886 355284 153892
rect 354876 150198 354950 150226
rect 348068 149926 348496 149954
rect 348804 149926 349140 149954
rect 349356 149926 349784 149954
rect 350092 149926 350428 149954
rect 350736 149926 351072 149954
rect 351380 149926 351716 149954
rect 352024 149926 352360 149954
rect 352576 149926 353004 149954
rect 353312 149926 353648 149954
rect 353864 149926 354292 149954
rect 354922 149940 354950 150198
rect 355244 149954 355272 153886
rect 355336 152114 355364 163200
rect 356060 159860 356112 159866
rect 356060 159802 356112 159808
rect 355968 159792 356020 159798
rect 355968 159734 356020 159740
rect 355980 159458 356008 159734
rect 355968 159452 356020 159458
rect 355968 159394 356020 159400
rect 356072 159050 356100 159802
rect 356164 159662 356192 163200
rect 356992 163146 357020 163200
rect 357084 163146 357112 163254
rect 356992 163118 357112 163146
rect 356152 159656 356204 159662
rect 356152 159598 356204 159604
rect 356060 159044 356112 159050
rect 356060 158986 356112 158992
rect 357360 153950 357388 163254
rect 357806 163200 357862 164400
rect 358634 163200 358690 164400
rect 359554 163200 359610 164400
rect 360382 163200 360438 164400
rect 361210 163200 361266 164400
rect 362038 163200 362094 164400
rect 362866 163200 362922 164400
rect 363694 163200 363750 164400
rect 364522 163200 364578 164400
rect 365442 163200 365498 164400
rect 366270 163200 366326 164400
rect 367098 163200 367154 164400
rect 367926 163200 367982 164400
rect 368754 163200 368810 164400
rect 369582 163200 369638 164400
rect 370410 163200 370466 164400
rect 371330 163200 371386 164400
rect 372158 163200 372214 164400
rect 372986 163200 373042 164400
rect 373814 163200 373870 164400
rect 374642 163200 374698 164400
rect 375470 163200 375526 164400
rect 376298 163200 376354 164400
rect 377218 163200 377274 164400
rect 378046 163200 378102 164400
rect 378874 163200 378930 164400
rect 379702 163200 379758 164400
rect 380530 163200 380586 164400
rect 380636 163254 380848 163282
rect 357820 159798 357848 163200
rect 357808 159792 357860 159798
rect 357808 159734 357860 159740
rect 358648 159458 358676 163200
rect 359464 159520 359516 159526
rect 359464 159462 359516 159468
rect 357992 159452 358044 159458
rect 357992 159394 358044 159400
rect 358636 159452 358688 159458
rect 358636 159394 358688 159400
rect 357808 154012 357860 154018
rect 357808 153954 357860 153960
rect 357348 153944 357400 153950
rect 357348 153886 357400 153892
rect 356060 152856 356112 152862
rect 356060 152798 356112 152804
rect 355324 152108 355376 152114
rect 355324 152050 355376 152056
rect 356072 149954 356100 152798
rect 356520 152720 356572 152726
rect 356520 152662 356572 152668
rect 356532 149954 356560 152662
rect 357438 152416 357494 152425
rect 357438 152351 357494 152360
rect 357452 150226 357480 152351
rect 357452 150198 357526 150226
rect 355244 149926 355580 149954
rect 356072 149926 356224 149954
rect 356532 149926 356868 149954
rect 357498 149940 357526 150198
rect 357820 149954 357848 153954
rect 358004 151814 358032 159394
rect 359476 159050 359504 159462
rect 359464 159044 359516 159050
rect 359464 158986 359516 158992
rect 358728 158976 358780 158982
rect 358728 158918 358780 158924
rect 358740 151814 358768 158918
rect 359568 152726 359596 163200
rect 360396 161474 360424 163200
rect 360396 161446 360516 161474
rect 359740 159860 359792 159866
rect 359740 159802 359792 159808
rect 359648 159656 359700 159662
rect 359648 159598 359700 159604
rect 359660 159458 359688 159598
rect 359648 159452 359700 159458
rect 359648 159394 359700 159400
rect 359556 152720 359608 152726
rect 359556 152662 359608 152668
rect 358004 151786 358400 151814
rect 358740 151786 359044 151814
rect 358372 149954 358400 151786
rect 359016 149954 359044 151786
rect 359752 149954 359780 159802
rect 360384 154080 360436 154086
rect 360384 154022 360436 154028
rect 360396 149954 360424 154022
rect 360488 154018 360516 161446
rect 361224 158846 361252 163200
rect 361120 158840 361172 158846
rect 361120 158782 361172 158788
rect 361212 158840 361264 158846
rect 361212 158782 361264 158788
rect 361132 158574 361160 158782
rect 361120 158568 361172 158574
rect 361120 158510 361172 158516
rect 360476 154012 360528 154018
rect 360476 153954 360528 153960
rect 361028 153196 361080 153202
rect 361028 153138 361080 153144
rect 361040 149954 361068 153138
rect 361672 153060 361724 153066
rect 361672 153002 361724 153008
rect 361684 149954 361712 153002
rect 362052 152862 362080 163200
rect 362880 159662 362908 163200
rect 362868 159656 362920 159662
rect 362868 159598 362920 159604
rect 363512 158976 363564 158982
rect 363512 158918 363564 158924
rect 362960 158568 363012 158574
rect 362960 158510 363012 158516
rect 362040 152856 362092 152862
rect 362040 152798 362092 152804
rect 362316 152040 362368 152046
rect 362316 151982 362368 151988
rect 362328 149954 362356 151982
rect 362972 151842 363000 158510
rect 363052 155372 363104 155378
rect 363052 155314 363104 155320
rect 362960 151836 363012 151842
rect 362960 151778 363012 151784
rect 363064 149954 363092 155314
rect 363524 149954 363552 158918
rect 363708 154086 363736 163200
rect 363696 154080 363748 154086
rect 363696 154022 363748 154028
rect 364536 153066 364564 163200
rect 365456 159798 365484 163200
rect 365352 159792 365404 159798
rect 365352 159734 365404 159740
rect 365444 159792 365496 159798
rect 365444 159734 365496 159740
rect 365364 158982 365392 159734
rect 364800 158976 364852 158982
rect 364800 158918 364852 158924
rect 365352 158976 365404 158982
rect 365352 158918 365404 158924
rect 364524 153060 364576 153066
rect 364524 153002 364576 153008
rect 364340 151836 364392 151842
rect 364340 151778 364392 151784
rect 364352 149954 364380 151778
rect 364812 149954 364840 158918
rect 365720 154148 365772 154154
rect 365720 154090 365772 154096
rect 365732 150226 365760 154090
rect 366284 153202 366312 163200
rect 367112 154154 367140 163200
rect 367940 158778 367968 163200
rect 367192 158772 367244 158778
rect 367192 158714 367244 158720
rect 367928 158772 367980 158778
rect 367928 158714 367980 158720
rect 367100 154148 367152 154154
rect 367100 154090 367152 154096
rect 367204 153202 367232 158714
rect 368020 154216 368072 154222
rect 368020 154158 368072 154164
rect 366272 153196 366324 153202
rect 366272 153138 366324 153144
rect 367192 153196 367244 153202
rect 367192 153138 367244 153144
rect 366732 153128 366784 153134
rect 366732 153070 366784 153076
rect 366088 152924 366140 152930
rect 366088 152866 366140 152872
rect 365732 150198 365806 150226
rect 357820 149926 358156 149954
rect 358372 149926 358800 149954
rect 359016 149926 359444 149954
rect 359752 149926 360088 149954
rect 360396 149926 360732 149954
rect 361040 149926 361376 149954
rect 361684 149926 362020 149954
rect 362328 149926 362664 149954
rect 363064 149926 363308 149954
rect 363524 149926 363952 149954
rect 364352 149926 364596 149954
rect 364812 149926 365240 149954
rect 365778 149940 365806 150198
rect 366100 149954 366128 152866
rect 366744 149954 366772 153070
rect 367376 152380 367428 152386
rect 367376 152322 367428 152328
rect 367388 149954 367416 152322
rect 368032 149954 368060 154158
rect 368664 153196 368716 153202
rect 368664 153138 368716 153144
rect 368676 149954 368704 153138
rect 368768 152930 368796 163200
rect 369216 159928 369268 159934
rect 369216 159870 369268 159876
rect 368756 152924 368808 152930
rect 368756 152866 368808 152872
rect 369228 149954 369256 159870
rect 369596 159730 369624 163200
rect 370044 159996 370096 160002
rect 370044 159938 370096 159944
rect 369584 159724 369636 159730
rect 369584 159666 369636 159672
rect 370056 149954 370084 159938
rect 370424 155242 370452 163200
rect 370596 155440 370648 155446
rect 370596 155382 370648 155388
rect 370412 155236 370464 155242
rect 370412 155178 370464 155184
rect 370608 149954 370636 155382
rect 371344 153202 371372 163200
rect 372172 160002 372200 163200
rect 372160 159996 372212 160002
rect 372160 159938 372212 159944
rect 371884 158976 371936 158982
rect 371884 158918 371936 158924
rect 371896 158846 371924 158918
rect 371884 158840 371936 158846
rect 371884 158782 371936 158788
rect 371332 153196 371384 153202
rect 371332 153138 371384 153144
rect 373000 152522 373028 163200
rect 373632 159928 373684 159934
rect 373632 159870 373684 159876
rect 373644 159186 373672 159870
rect 373632 159180 373684 159186
rect 373632 159122 373684 159128
rect 373080 155508 373132 155514
rect 373080 155450 373132 155456
rect 371240 152516 371292 152522
rect 371240 152458 371292 152464
rect 372988 152516 373040 152522
rect 372988 152458 373040 152464
rect 371252 149954 371280 152458
rect 372620 152448 372672 152454
rect 372620 152390 372672 152396
rect 371884 151972 371936 151978
rect 371884 151914 371936 151920
rect 371896 149954 371924 151914
rect 372632 149954 372660 152390
rect 373092 149954 373120 155450
rect 373828 155310 373856 163200
rect 374460 160064 374512 160070
rect 374460 160006 374512 160012
rect 374092 159316 374144 159322
rect 374092 159258 374144 159264
rect 373816 155304 373868 155310
rect 373816 155246 373868 155252
rect 374104 150226 374132 159258
rect 374104 150198 374178 150226
rect 366100 149926 366436 149954
rect 366744 149926 367080 149954
rect 367388 149926 367724 149954
rect 368032 149926 368368 149954
rect 368676 149926 369012 149954
rect 369228 149926 369656 149954
rect 370056 149926 370300 149954
rect 370608 149926 370944 149954
rect 371252 149926 371588 149954
rect 371896 149926 372232 149954
rect 372632 149926 372876 149954
rect 373092 149926 373520 149954
rect 374150 149940 374178 150198
rect 374472 149954 374500 160006
rect 374656 159916 374684 163200
rect 374656 159888 374868 159916
rect 374736 159384 374788 159390
rect 374736 159326 374788 159332
rect 374552 158976 374604 158982
rect 374552 158918 374604 158924
rect 374564 158710 374592 158918
rect 374748 158778 374776 159326
rect 374840 158846 374868 159888
rect 374828 158840 374880 158846
rect 374828 158782 374880 158788
rect 374736 158772 374788 158778
rect 374736 158714 374788 158720
rect 374552 158704 374604 158710
rect 374552 158646 374604 158652
rect 375484 152454 375512 163200
rect 376312 159866 376340 163200
rect 376300 159860 376352 159866
rect 376300 159802 376352 159808
rect 376300 155576 376352 155582
rect 376300 155518 376352 155524
rect 375748 153876 375800 153882
rect 375748 153818 375800 153824
rect 375472 152448 375524 152454
rect 375472 152390 375524 152396
rect 375380 152244 375432 152250
rect 375380 152186 375432 152192
rect 375392 150226 375420 152186
rect 375392 150198 375466 150226
rect 374472 149926 374808 149954
rect 375438 149940 375466 150198
rect 375760 149954 375788 153818
rect 376312 149954 376340 155518
rect 377232 153882 377260 163200
rect 378060 159322 378088 163200
rect 378888 160070 378916 163200
rect 378876 160064 378928 160070
rect 378876 160006 378928 160012
rect 379716 159934 379744 163200
rect 380544 163146 380572 163200
rect 380636 163146 380664 163254
rect 380544 163118 380664 163146
rect 379428 159928 379480 159934
rect 379428 159870 379480 159876
rect 379704 159928 379756 159934
rect 379704 159870 379756 159876
rect 378048 159316 378100 159322
rect 378048 159258 378100 159264
rect 377588 159180 377640 159186
rect 377588 159122 377640 159128
rect 377220 153876 377272 153882
rect 377220 153818 377272 153824
rect 377036 152992 377088 152998
rect 377036 152934 377088 152940
rect 377048 149954 377076 152934
rect 377600 149954 377628 159122
rect 378784 159044 378836 159050
rect 378784 158986 378836 158992
rect 378692 155712 378744 155718
rect 378692 155654 378744 155660
rect 378324 154352 378376 154358
rect 378324 154294 378376 154300
rect 378336 149954 378364 154294
rect 378704 151814 378732 155654
rect 378796 151978 378824 158986
rect 378784 151972 378836 151978
rect 378784 151914 378836 151920
rect 379440 151814 379468 159870
rect 380820 154222 380848 163254
rect 381358 163200 381414 164400
rect 382186 163200 382242 164400
rect 383106 163200 383162 164400
rect 383934 163200 383990 164400
rect 384762 163200 384818 164400
rect 385590 163200 385646 164400
rect 386418 163200 386474 164400
rect 387246 163200 387302 164400
rect 387352 163254 387656 163282
rect 380900 154284 380952 154290
rect 380900 154226 380952 154232
rect 380808 154216 380860 154222
rect 380808 154158 380860 154164
rect 380256 152176 380308 152182
rect 380256 152118 380308 152124
rect 378704 151786 378916 151814
rect 379440 151786 379560 151814
rect 378888 149954 378916 151786
rect 379532 149954 379560 151786
rect 380268 149954 380296 152118
rect 380912 149954 380940 154226
rect 381372 152386 381400 163200
rect 381452 155644 381504 155650
rect 381452 155586 381504 155592
rect 381360 152380 381412 152386
rect 381360 152322 381412 152328
rect 381464 149954 381492 155586
rect 382200 152998 382228 163200
rect 382740 159248 382792 159254
rect 382740 159190 382792 159196
rect 382372 159112 382424 159118
rect 382372 159054 382424 159060
rect 382188 152992 382240 152998
rect 382188 152934 382240 152940
rect 382384 152318 382412 159054
rect 382280 152312 382332 152318
rect 382280 152254 382332 152260
rect 382372 152312 382424 152318
rect 382372 152254 382424 152260
rect 382292 149954 382320 152254
rect 382752 149954 382780 159190
rect 383120 159050 383148 163200
rect 383108 159044 383160 159050
rect 383108 158986 383160 158992
rect 383660 158840 383712 158846
rect 383712 158788 383792 158794
rect 383660 158782 383792 158788
rect 383672 158766 383792 158782
rect 383660 154420 383712 154426
rect 383660 154362 383712 154368
rect 383672 149954 383700 154362
rect 383764 152182 383792 158766
rect 383948 154290 383976 163200
rect 384776 158914 384804 163200
rect 385500 159588 385552 159594
rect 385500 159530 385552 159536
rect 384764 158908 384816 158914
rect 384764 158850 384816 158856
rect 383936 154284 383988 154290
rect 383936 154226 383988 154232
rect 385040 152584 385092 152590
rect 385040 152526 385092 152532
rect 383752 152176 383804 152182
rect 383752 152118 383804 152124
rect 384120 151972 384172 151978
rect 384120 151914 384172 151920
rect 384132 149954 384160 151914
rect 385052 150226 385080 152526
rect 385512 152250 385540 159530
rect 385604 159254 385632 163200
rect 385868 159384 385920 159390
rect 385868 159326 385920 159332
rect 385592 159248 385644 159254
rect 385592 159190 385644 159196
rect 385500 152244 385552 152250
rect 385500 152186 385552 152192
rect 385880 151978 385908 159326
rect 386328 158976 386380 158982
rect 386328 158918 386380 158924
rect 386052 154488 386104 154494
rect 386052 154430 386104 154436
rect 385868 151972 385920 151978
rect 385868 151914 385920 151920
rect 385408 151836 385460 151842
rect 385408 151778 385460 151784
rect 385052 150198 385126 150226
rect 375760 149926 376096 149954
rect 376312 149926 376740 149954
rect 377048 149926 377384 149954
rect 377600 149926 378028 149954
rect 378336 149926 378672 149954
rect 378888 149926 379316 149954
rect 379532 149926 379960 149954
rect 380268 149926 380604 149954
rect 380912 149926 381248 149954
rect 381464 149926 381892 149954
rect 382292 149926 382536 149954
rect 382752 149926 383180 149954
rect 383672 149926 383824 149954
rect 384132 149926 384468 149954
rect 385098 149940 385126 150198
rect 385420 149954 385448 151778
rect 386064 149954 386092 154430
rect 386340 151910 386368 158918
rect 386432 152590 386460 163200
rect 387260 163146 387288 163200
rect 387352 163146 387380 163254
rect 387260 163118 387380 163146
rect 387628 154358 387656 163254
rect 388074 163200 388130 164400
rect 388994 163200 389050 164400
rect 389822 163200 389878 164400
rect 390650 163200 390706 164400
rect 391478 163200 391534 164400
rect 392306 163200 392362 164400
rect 393134 163200 393190 164400
rect 393962 163200 394018 164400
rect 394882 163200 394938 164400
rect 395710 163200 395766 164400
rect 396538 163200 396594 164400
rect 397366 163200 397422 164400
rect 398194 163200 398250 164400
rect 399022 163200 399078 164400
rect 399850 163200 399906 164400
rect 399956 163254 400168 163282
rect 388088 158846 388116 163200
rect 389008 159390 389036 163200
rect 389836 159594 389864 163200
rect 389824 159588 389876 159594
rect 389824 159530 389876 159536
rect 388996 159384 389048 159390
rect 388996 159326 389048 159332
rect 388352 159316 388404 159322
rect 388352 159258 388404 159264
rect 387892 158840 387944 158846
rect 387892 158782 387944 158788
rect 388076 158840 388128 158846
rect 388076 158782 388128 158788
rect 387616 154352 387668 154358
rect 387616 154294 387668 154300
rect 386420 152584 386472 152590
rect 386420 152526 386472 152532
rect 386696 152312 386748 152318
rect 386696 152254 386748 152260
rect 386328 151904 386380 151910
rect 386328 151846 386380 151852
rect 386708 149954 386736 152254
rect 387340 152244 387392 152250
rect 387340 152186 387392 152192
rect 387352 149954 387380 152186
rect 387904 152046 387932 158782
rect 387984 152788 388036 152794
rect 387984 152730 388036 152736
rect 387892 152040 387944 152046
rect 387892 151982 387944 151988
rect 387996 149954 388024 152730
rect 388364 152250 388392 159258
rect 389180 158908 389232 158914
rect 389180 158850 389232 158856
rect 388628 154556 388680 154562
rect 388628 154498 388680 154504
rect 388352 152244 388404 152250
rect 388352 152186 388404 152192
rect 388640 149954 388668 154498
rect 389192 152318 389220 158850
rect 390376 158840 390428 158846
rect 390376 158782 390428 158788
rect 390388 152794 390416 158782
rect 390664 154426 390692 163200
rect 390744 159452 390796 159458
rect 390744 159394 390796 159400
rect 390652 154420 390704 154426
rect 390652 154362 390704 154368
rect 390376 152788 390428 152794
rect 390376 152730 390428 152736
rect 389272 152652 389324 152658
rect 389272 152594 389324 152600
rect 389180 152312 389232 152318
rect 389180 152254 389232 152260
rect 389284 149954 389312 152594
rect 389916 152108 389968 152114
rect 389916 152050 389968 152056
rect 389928 149954 389956 152050
rect 390756 149954 390784 159394
rect 391492 158982 391520 163200
rect 392320 159186 392348 163200
rect 392400 159520 392452 159526
rect 392400 159462 392452 159468
rect 392308 159180 392360 159186
rect 392308 159122 392360 159128
rect 391480 158976 391532 158982
rect 391480 158918 391532 158924
rect 391204 153944 391256 153950
rect 391204 153886 391256 153892
rect 391216 149954 391244 153886
rect 391940 152176 391992 152182
rect 391940 152118 391992 152124
rect 391952 149954 391980 152118
rect 392412 149954 392440 159462
rect 393148 152658 393176 163200
rect 393780 154012 393832 154018
rect 393780 153954 393832 153960
rect 393320 152720 393372 152726
rect 393320 152662 393372 152668
rect 393136 152652 393188 152658
rect 393136 152594 393188 152600
rect 393332 149954 393360 152662
rect 393792 149954 393820 153954
rect 393976 153950 394004 163200
rect 394608 158976 394660 158982
rect 394608 158918 394660 158924
rect 393964 153944 394016 153950
rect 393964 153886 394016 153892
rect 394620 152250 394648 158918
rect 394896 152726 394924 163200
rect 395160 159792 395212 159798
rect 395160 159734 395212 159740
rect 395172 152862 395200 159734
rect 395252 159656 395304 159662
rect 395252 159598 395304 159604
rect 395068 152856 395120 152862
rect 395068 152798 395120 152804
rect 395160 152856 395212 152862
rect 395160 152798 395212 152804
rect 394884 152720 394936 152726
rect 394884 152662 394936 152668
rect 394608 152244 394660 152250
rect 394608 152186 394660 152192
rect 394700 151904 394752 151910
rect 394700 151846 394752 151852
rect 394712 150226 394740 151846
rect 394712 150198 394786 150226
rect 385420 149926 385756 149954
rect 386064 149926 386400 149954
rect 386708 149926 387044 149954
rect 387352 149926 387688 149954
rect 387996 149926 388332 149954
rect 388640 149926 388976 149954
rect 389284 149926 389620 149954
rect 389928 149926 390264 149954
rect 390756 149926 390908 149954
rect 391216 149926 391552 149954
rect 391952 149926 392196 149954
rect 392412 149926 392840 149954
rect 393332 149926 393484 149954
rect 393792 149926 394128 149954
rect 394758 149940 394786 150198
rect 395080 149954 395108 152798
rect 395264 151814 395292 159598
rect 395724 159118 395752 163200
rect 396264 159996 396316 160002
rect 396264 159938 396316 159944
rect 395712 159112 395764 159118
rect 395712 159054 395764 159060
rect 396276 151910 396304 159938
rect 396552 159798 396580 163200
rect 396540 159792 396592 159798
rect 396540 159734 396592 159740
rect 396356 154080 396408 154086
rect 396356 154022 396408 154028
rect 396264 151904 396316 151910
rect 396264 151846 396316 151852
rect 395264 151786 395660 151814
rect 395632 149954 395660 151786
rect 396368 149954 396396 154022
rect 397380 154018 397408 163200
rect 398104 160064 398156 160070
rect 398104 160006 398156 160012
rect 397368 154012 397420 154018
rect 397368 153954 397420 153960
rect 398116 153134 398144 160006
rect 398208 154086 398236 163200
rect 399036 159662 399064 163200
rect 399864 163146 399892 163200
rect 399956 163146 399984 163254
rect 399864 163118 399984 163146
rect 399024 159656 399076 159662
rect 399024 159598 399076 159604
rect 399576 159248 399628 159254
rect 399576 159190 399628 159196
rect 398840 154148 398892 154154
rect 398840 154090 398892 154096
rect 398196 154080 398248 154086
rect 398196 154022 398248 154028
rect 397920 153128 397972 153134
rect 397920 153070 397972 153076
rect 398104 153128 398156 153134
rect 398104 153070 398156 153076
rect 396908 153060 396960 153066
rect 396908 153002 396960 153008
rect 396920 149954 396948 153002
rect 397552 152856 397604 152862
rect 397552 152798 397604 152804
rect 397564 149954 397592 152798
rect 397932 151814 397960 153070
rect 397932 151786 398144 151814
rect 398116 149954 398144 151786
rect 398852 149954 398880 154090
rect 399588 151978 399616 159190
rect 400140 152862 400168 163254
rect 400770 163200 400826 164400
rect 401598 163200 401654 164400
rect 402426 163200 402482 164400
rect 403254 163200 403310 164400
rect 404082 163200 404138 164400
rect 404910 163200 404966 164400
rect 405738 163200 405794 164400
rect 406658 163200 406714 164400
rect 406764 163254 407068 163282
rect 400680 159724 400732 159730
rect 400680 159666 400732 159672
rect 400220 152924 400272 152930
rect 400220 152866 400272 152872
rect 400128 152856 400180 152862
rect 400128 152798 400180 152804
rect 399484 151972 399536 151978
rect 399484 151914 399536 151920
rect 399576 151972 399628 151978
rect 399576 151914 399628 151920
rect 399496 149954 399524 151914
rect 400232 149954 400260 152866
rect 400692 149954 400720 159666
rect 400784 159458 400812 163200
rect 400772 159452 400824 159458
rect 400772 159394 400824 159400
rect 401612 154154 401640 163200
rect 401692 155236 401744 155242
rect 401692 155178 401744 155184
rect 401600 154148 401652 154154
rect 401600 154090 401652 154096
rect 401704 150226 401732 155178
rect 402060 153196 402112 153202
rect 402060 153138 402112 153144
rect 401704 150198 401778 150226
rect 395080 149926 395416 149954
rect 395632 149926 396060 149954
rect 396368 149926 396612 149954
rect 396920 149926 397256 149954
rect 397564 149926 397900 149954
rect 398116 149926 398544 149954
rect 398852 149926 399188 149954
rect 399496 149926 399832 149954
rect 400232 149926 400476 149954
rect 400692 149926 401120 149954
rect 401750 149940 401778 150198
rect 402072 149954 402100 153138
rect 402440 152930 402468 163200
rect 403268 160002 403296 163200
rect 403256 159996 403308 160002
rect 403256 159938 403308 159944
rect 403900 159384 403952 159390
rect 403900 159326 403952 159332
rect 403532 155304 403584 155310
rect 403532 155246 403584 155252
rect 402428 152924 402480 152930
rect 402428 152866 402480 152872
rect 403348 152516 403400 152522
rect 403348 152458 403400 152464
rect 402980 151904 403032 151910
rect 402980 151846 403032 151852
rect 402992 150226 403020 151846
rect 402992 150198 403066 150226
rect 402072 149926 402408 149954
rect 403038 149940 403066 150198
rect 403360 149954 403388 152458
rect 403544 151814 403572 155246
rect 403912 151842 403940 159326
rect 404096 159322 404124 163200
rect 404084 159316 404136 159322
rect 404084 159258 404136 159264
rect 404268 159180 404320 159186
rect 404268 159122 404320 159128
rect 404280 151910 404308 159122
rect 404924 152522 404952 163200
rect 405648 159112 405700 159118
rect 405648 159054 405700 159060
rect 404912 152516 404964 152522
rect 404912 152458 404964 152464
rect 405280 152448 405332 152454
rect 405280 152390 405332 152396
rect 404636 152040 404688 152046
rect 404636 151982 404688 151988
rect 404268 151904 404320 151910
rect 404268 151846 404320 151852
rect 403900 151836 403952 151842
rect 403544 151786 403848 151814
rect 403820 150498 403848 151786
rect 403900 151778 403952 151784
rect 403820 150470 403940 150498
rect 403912 149954 403940 150470
rect 404648 149954 404676 151982
rect 405292 149954 405320 152390
rect 405660 152114 405688 159054
rect 405752 158914 405780 163200
rect 406672 163146 406700 163200
rect 406764 163146 406792 163254
rect 406672 163118 406792 163146
rect 405832 159928 405884 159934
rect 405832 159870 405884 159876
rect 405740 158908 405792 158914
rect 405740 158850 405792 158856
rect 405844 153134 405872 159870
rect 405924 159860 405976 159866
rect 405924 159802 405976 159808
rect 405832 153128 405884 153134
rect 405832 153070 405884 153076
rect 405648 152108 405700 152114
rect 405648 152050 405700 152056
rect 405936 149954 405964 159802
rect 406568 153876 406620 153882
rect 406568 153818 406620 153824
rect 406580 149954 406608 153818
rect 407040 153066 407068 163254
rect 407486 163200 407542 164400
rect 408314 163200 408370 164400
rect 409142 163200 409198 164400
rect 409970 163200 410026 164400
rect 410798 163200 410854 164400
rect 411626 163200 411682 164400
rect 412546 163200 412602 164400
rect 413374 163200 413430 164400
rect 414202 163200 414258 164400
rect 415030 163200 415086 164400
rect 415136 163254 415348 163282
rect 407500 159730 407528 163200
rect 407488 159724 407540 159730
rect 407488 159666 407540 159672
rect 407856 153196 407908 153202
rect 407856 153138 407908 153144
rect 407028 153060 407080 153066
rect 407028 153002 407080 153008
rect 407212 152176 407264 152182
rect 407212 152118 407264 152124
rect 407224 149954 407252 152118
rect 407868 149954 407896 153138
rect 408328 152425 408356 163200
rect 408592 159656 408644 159662
rect 408592 159598 408644 159604
rect 408500 153128 408552 153134
rect 408500 153070 408552 153076
rect 408314 152416 408370 152425
rect 408314 152351 408370 152360
rect 408512 149954 408540 153070
rect 408604 152454 408632 159598
rect 409156 158982 409184 163200
rect 409984 159934 410012 163200
rect 409972 159928 410024 159934
rect 409972 159870 410024 159876
rect 410812 159662 410840 163200
rect 410800 159656 410852 159662
rect 410800 159598 410852 159604
rect 411444 159044 411496 159050
rect 411444 158986 411496 158992
rect 409144 158976 409196 158982
rect 409144 158918 409196 158924
rect 410892 158976 410944 158982
rect 410892 158918 410944 158924
rect 409328 158908 409380 158914
rect 409328 158850 409380 158856
rect 409236 154216 409288 154222
rect 409236 154158 409288 154164
rect 408592 152448 408644 152454
rect 408592 152390 408644 152396
rect 409248 149954 409276 154158
rect 409340 152182 409368 158850
rect 410904 152998 410932 158918
rect 410432 152992 410484 152998
rect 410432 152934 410484 152940
rect 410892 152992 410944 152998
rect 410892 152934 410944 152940
rect 409880 152380 409932 152386
rect 409880 152322 409932 152328
rect 409328 152176 409380 152182
rect 409328 152118 409380 152124
rect 409892 149954 409920 152322
rect 410444 149954 410472 152934
rect 411456 150226 411484 158986
rect 411640 153134 411668 163200
rect 412560 159118 412588 163200
rect 412548 159112 412600 159118
rect 412548 159054 412600 159060
rect 413388 158778 413416 163200
rect 413744 159792 413796 159798
rect 413744 159734 413796 159740
rect 413376 158772 413428 158778
rect 413376 158714 413428 158720
rect 411720 154284 411772 154290
rect 411720 154226 411772 154232
rect 411628 153128 411680 153134
rect 411628 153070 411680 153076
rect 411410 150198 411484 150226
rect 403360 149926 403696 149954
rect 403912 149926 404340 149954
rect 404648 149926 404984 149954
rect 405292 149926 405628 149954
rect 405936 149926 406272 149954
rect 406580 149926 406916 149954
rect 407224 149926 407560 149954
rect 407868 149926 408204 149954
rect 408512 149926 408848 149954
rect 409248 149926 409492 149954
rect 409892 149926 410136 149954
rect 410444 149926 410780 149954
rect 411410 149940 411438 150198
rect 411732 149954 411760 154226
rect 413652 152584 413704 152590
rect 413652 152526 413704 152532
rect 412640 152312 412692 152318
rect 412640 152254 412692 152260
rect 412652 150226 412680 152254
rect 413008 152040 413060 152046
rect 413008 151982 413060 151988
rect 412652 150198 412726 150226
rect 411732 149926 412068 149954
rect 412698 149940 412726 150198
rect 413020 149954 413048 151982
rect 413664 149954 413692 152526
rect 413756 151978 413784 159734
rect 414216 159594 414244 163200
rect 415044 163146 415072 163200
rect 415136 163146 415164 163254
rect 415044 163118 415164 163146
rect 413836 159588 413888 159594
rect 413836 159530 413888 159536
rect 414204 159588 414256 159594
rect 414204 159530 414256 159536
rect 413848 152386 413876 159530
rect 413928 159112 413980 159118
rect 413928 159054 413980 159060
rect 413940 152590 413968 159054
rect 414296 154352 414348 154358
rect 414296 154294 414348 154300
rect 413928 152584 413980 152590
rect 413928 152526 413980 152532
rect 413836 152380 413888 152386
rect 413836 152322 413888 152328
rect 413744 151972 413796 151978
rect 413744 151914 413796 151920
rect 414308 149954 414336 154294
rect 415320 153202 415348 163254
rect 415858 163200 415914 164400
rect 416686 163200 416742 164400
rect 417514 163200 417570 164400
rect 418434 163200 418490 164400
rect 419262 163200 419318 164400
rect 420090 163200 420146 164400
rect 420918 163200 420974 164400
rect 421746 163200 421802 164400
rect 422574 163200 422630 164400
rect 423402 163200 423458 164400
rect 424322 163200 424378 164400
rect 425150 163200 425206 164400
rect 425978 163200 426034 164400
rect 426084 163254 426296 163282
rect 415308 153196 415360 153202
rect 415308 153138 415360 153144
rect 415872 152794 415900 163200
rect 416596 159996 416648 160002
rect 416596 159938 416648 159944
rect 414940 152788 414992 152794
rect 414940 152730 414992 152736
rect 415860 152788 415912 152794
rect 415860 152730 415912 152736
rect 414952 149954 414980 152730
rect 416608 152386 416636 159938
rect 416700 158914 416728 163200
rect 417528 159390 417556 163200
rect 417608 159928 417660 159934
rect 417608 159870 417660 159876
rect 417516 159384 417568 159390
rect 417516 159326 417568 159332
rect 416688 158908 416740 158914
rect 416688 158850 416740 158856
rect 416872 154420 416924 154426
rect 416872 154362 416924 154368
rect 416228 152380 416280 152386
rect 416228 152322 416280 152328
rect 416596 152380 416648 152386
rect 416596 152322 416648 152328
rect 415676 151836 415728 151842
rect 415676 151778 415728 151784
rect 415688 149954 415716 151778
rect 416240 149954 416268 152322
rect 416884 149954 416912 154362
rect 417424 152448 417476 152454
rect 417424 152390 417476 152396
rect 417332 152244 417384 152250
rect 417332 152186 417384 152192
rect 417344 151814 417372 152186
rect 417436 152114 417464 152390
rect 417620 152318 417648 159870
rect 418448 152454 418476 163200
rect 419276 152658 419304 163200
rect 420104 158982 420132 163200
rect 420932 159798 420960 163200
rect 420920 159792 420972 159798
rect 420920 159734 420972 159740
rect 420092 158976 420144 158982
rect 420092 158918 420144 158924
rect 419632 158908 419684 158914
rect 419632 158850 419684 158856
rect 419540 153944 419592 153950
rect 419540 153886 419592 153892
rect 418804 152652 418856 152658
rect 418804 152594 418856 152600
rect 419264 152652 419316 152658
rect 419264 152594 419316 152600
rect 418436 152448 418488 152454
rect 418436 152390 418488 152396
rect 417608 152312 417660 152318
rect 417608 152254 417660 152260
rect 417424 152108 417476 152114
rect 417424 152050 417476 152056
rect 418160 151904 418212 151910
rect 418160 151846 418212 151852
rect 417344 151786 417464 151814
rect 417436 149954 417464 151786
rect 418172 149954 418200 151846
rect 418816 149954 418844 152594
rect 419552 149954 419580 153886
rect 419644 151978 419672 158850
rect 419724 158772 419776 158778
rect 419724 158714 419776 158720
rect 419632 151972 419684 151978
rect 419632 151914 419684 151920
rect 419736 151842 419764 158714
rect 420092 152720 420144 152726
rect 420092 152662 420144 152668
rect 419724 151836 419776 151842
rect 419724 151778 419776 151784
rect 420104 149954 420132 152662
rect 421760 152386 421788 163200
rect 422300 154012 422352 154018
rect 422300 153954 422352 153960
rect 421748 152380 421800 152386
rect 421748 152322 421800 152328
rect 421472 152312 421524 152318
rect 421472 152254 421524 152260
rect 420920 152040 420972 152046
rect 420920 151982 420972 151988
rect 420932 149954 420960 151982
rect 421484 151910 421512 152254
rect 421380 151904 421432 151910
rect 421380 151846 421432 151852
rect 421472 151904 421524 151910
rect 421472 151846 421524 151852
rect 421392 149954 421420 151846
rect 422312 150226 422340 153954
rect 422588 152114 422616 163200
rect 422668 154080 422720 154086
rect 422668 154022 422720 154028
rect 422576 152108 422628 152114
rect 422576 152050 422628 152056
rect 422312 150198 422386 150226
rect 413020 149926 413356 149954
rect 413664 149926 414000 149954
rect 414308 149926 414644 149954
rect 414952 149926 415288 149954
rect 415688 149926 415932 149954
rect 416240 149926 416576 149954
rect 416884 149926 417220 149954
rect 417436 149926 417864 149954
rect 418172 149926 418508 149954
rect 418816 149926 419152 149954
rect 419552 149926 419796 149954
rect 420104 149926 420440 149954
rect 420932 149926 421084 149954
rect 421392 149926 421728 149954
rect 422358 149940 422386 150198
rect 422680 149954 422708 154022
rect 423416 152726 423444 163200
rect 424336 159526 424364 163200
rect 424324 159520 424376 159526
rect 424324 159462 424376 159468
rect 424508 159452 424560 159458
rect 424508 159394 424560 159400
rect 423588 158976 423640 158982
rect 423588 158918 423640 158924
rect 423404 152720 423456 152726
rect 423404 152662 423456 152668
rect 423600 152046 423628 158918
rect 423956 152856 424008 152862
rect 423956 152798 424008 152804
rect 423312 152040 423364 152046
rect 423312 151982 423364 151988
rect 423588 152040 423640 152046
rect 423588 151982 423640 151988
rect 423324 149954 423352 151982
rect 423968 149954 423996 152798
rect 424520 149954 424548 159394
rect 425164 152318 425192 163200
rect 425992 163146 426020 163200
rect 426084 163146 426112 163254
rect 425992 163118 426112 163146
rect 425336 154148 425388 154154
rect 425336 154090 425388 154096
rect 425152 152312 425204 152318
rect 425152 152254 425204 152260
rect 425348 149954 425376 154090
rect 425888 152924 425940 152930
rect 425888 152866 425940 152872
rect 425900 149954 425928 152866
rect 426268 152862 426296 163254
rect 426806 163200 426862 164400
rect 427634 163200 427690 164400
rect 428462 163200 428518 164400
rect 429290 163200 429346 164400
rect 430210 163200 430266 164400
rect 431038 163200 431094 164400
rect 431866 163200 431922 164400
rect 432694 163200 432750 164400
rect 433522 163200 433578 164400
rect 434350 163200 434406 164400
rect 434456 163254 434668 163282
rect 426256 152856 426308 152862
rect 426256 152798 426308 152804
rect 426716 152312 426768 152318
rect 426716 152254 426768 152260
rect 426532 152244 426584 152250
rect 426532 152186 426584 152192
rect 426544 149954 426572 152186
rect 426728 152114 426756 152254
rect 426820 152114 426848 163200
rect 427648 159458 427676 163200
rect 427636 159452 427688 159458
rect 427636 159394 427688 159400
rect 426992 159316 427044 159322
rect 426992 159258 427044 159264
rect 426716 152108 426768 152114
rect 426716 152050 426768 152056
rect 426808 152108 426860 152114
rect 426808 152050 426860 152056
rect 427004 149954 427032 159258
rect 428476 152930 428504 163200
rect 429200 153060 429252 153066
rect 429200 153002 429252 153008
rect 428464 152924 428516 152930
rect 428464 152866 428516 152872
rect 427820 152516 427872 152522
rect 427820 152458 427872 152464
rect 427832 149954 427860 152458
rect 428372 152176 428424 152182
rect 428372 152118 428424 152124
rect 428384 149954 428412 152118
rect 429212 149954 429240 153002
rect 429304 152182 429332 163200
rect 429568 159724 429620 159730
rect 429568 159666 429620 159672
rect 429292 152176 429344 152182
rect 429292 152118 429344 152124
rect 429580 149954 429608 159666
rect 430224 152522 430252 163200
rect 431052 152998 431080 163200
rect 430948 152992 431000 152998
rect 430948 152934 431000 152940
rect 431040 152992 431092 152998
rect 431040 152934 431092 152940
rect 430212 152516 430264 152522
rect 430212 152458 430264 152464
rect 430578 152416 430634 152425
rect 430578 152351 430634 152360
rect 430592 150226 430620 152351
rect 430592 150198 430666 150226
rect 422680 149926 423016 149954
rect 423324 149926 423660 149954
rect 423968 149926 424304 149954
rect 424520 149926 424948 149954
rect 425348 149926 425592 149954
rect 425900 149926 426236 149954
rect 426544 149926 426880 149954
rect 427004 149926 427432 149954
rect 427832 149926 428076 149954
rect 428384 149926 428720 149954
rect 429212 149926 429364 149954
rect 429580 149926 430008 149954
rect 430638 149940 430666 150198
rect 430960 149954 430988 152934
rect 431880 152425 431908 163200
rect 432144 159656 432196 159662
rect 432144 159598 432196 159604
rect 431866 152416 431922 152425
rect 431866 152351 431922 152360
rect 431592 151904 431644 151910
rect 431592 151846 431644 151852
rect 431604 149954 431632 151846
rect 432156 149954 432184 159598
rect 432708 153134 432736 163200
rect 432696 153128 432748 153134
rect 432696 153070 432748 153076
rect 433536 153066 433564 163200
rect 434364 163146 434392 163200
rect 434456 163146 434484 163254
rect 434364 163118 434484 163146
rect 432880 153060 432932 153066
rect 432880 153002 432932 153008
rect 433524 153060 433576 153066
rect 433524 153002 433576 153008
rect 432892 149954 432920 153002
rect 434640 152590 434668 163254
rect 435178 163200 435234 164400
rect 436098 163200 436154 164400
rect 436926 163200 436982 164400
rect 437032 163254 437336 163282
rect 434812 159588 434864 159594
rect 434812 159530 434864 159536
rect 433524 152584 433576 152590
rect 433524 152526 433576 152532
rect 434628 152584 434680 152590
rect 434628 152526 434680 152532
rect 433536 149954 433564 152526
rect 434168 151836 434220 151842
rect 434168 151778 434220 151784
rect 434180 149954 434208 151778
rect 434824 149954 434852 159530
rect 435192 153814 435220 163200
rect 436112 161474 436140 163200
rect 436940 163146 436968 163200
rect 437032 163146 437060 163254
rect 436940 163118 437060 163146
rect 436112 161446 436232 161474
rect 435180 153808 435232 153814
rect 435180 153750 435232 153756
rect 435456 153196 435508 153202
rect 435456 153138 435508 153144
rect 435468 149954 435496 153138
rect 436100 152788 436152 152794
rect 436100 152730 436152 152736
rect 436112 149954 436140 152730
rect 436204 151842 436232 161446
rect 437308 152794 437336 163254
rect 437754 163200 437810 164400
rect 438582 163200 438638 164400
rect 439410 163200 439466 164400
rect 440238 163200 440294 164400
rect 441066 163200 441122 164400
rect 441986 163200 442042 164400
rect 442814 163200 442870 164400
rect 443642 163200 443698 164400
rect 444470 163200 444526 164400
rect 445298 163200 445354 164400
rect 445404 163254 445708 163282
rect 437664 159384 437716 159390
rect 437664 159326 437716 159332
rect 437296 152788 437348 152794
rect 437296 152730 437348 152736
rect 436284 152380 436336 152386
rect 436284 152322 436336 152328
rect 436296 151910 436324 152322
rect 436744 151972 436796 151978
rect 436744 151914 436796 151920
rect 436284 151904 436336 151910
rect 436284 151846 436336 151852
rect 436192 151836 436244 151842
rect 436192 151778 436244 151784
rect 436756 149954 436784 151914
rect 437676 150226 437704 159326
rect 437768 153202 437796 163200
rect 437756 153196 437808 153202
rect 437756 153138 437808 153144
rect 438596 152454 438624 163200
rect 438860 152652 438912 152658
rect 438860 152594 438912 152600
rect 438032 152448 438084 152454
rect 438032 152390 438084 152396
rect 438584 152448 438636 152454
rect 438584 152390 438636 152396
rect 437676 150198 437750 150226
rect 430960 149926 431296 149954
rect 431604 149926 431940 149954
rect 432156 149926 432584 149954
rect 432892 149926 433228 149954
rect 433536 149926 433872 149954
rect 434180 149926 434516 149954
rect 434824 149926 435160 149954
rect 435468 149926 435804 149954
rect 436112 149926 436448 149954
rect 436756 149926 437092 149954
rect 437722 149940 437750 150198
rect 438044 149954 438072 152390
rect 438872 149954 438900 152594
rect 439424 152046 439452 163200
rect 439502 152960 439558 152969
rect 440252 152930 440280 163200
rect 440424 159792 440476 159798
rect 440424 159734 440476 159740
rect 439502 152895 439504 152904
rect 439556 152895 439558 152904
rect 440240 152924 440292 152930
rect 439504 152866 439556 152872
rect 440240 152866 440292 152872
rect 439320 152040 439372 152046
rect 439320 151982 439372 151988
rect 439412 152040 439464 152046
rect 439412 151982 439464 151988
rect 439332 149954 439360 151982
rect 440436 149954 440464 159734
rect 441080 157334 441108 163200
rect 441080 157306 441384 157334
rect 441252 152380 441304 152386
rect 441252 152322 441304 152328
rect 440608 151904 440660 151910
rect 440608 151846 440660 151852
rect 438044 149926 438380 149954
rect 438872 149926 439024 149954
rect 439332 149926 439668 149954
rect 440312 149926 440464 149954
rect 440620 149954 440648 151846
rect 441264 149954 441292 152322
rect 441356 152130 441384 157306
rect 442000 152930 442028 163200
rect 442448 159520 442500 159526
rect 442448 159462 442500 159468
rect 441528 152924 441580 152930
rect 441528 152866 441580 152872
rect 441988 152924 442040 152930
rect 441988 152866 442040 152872
rect 441540 152318 441568 152866
rect 441896 152720 441948 152726
rect 441896 152662 441948 152668
rect 441712 152380 441764 152386
rect 441712 152322 441764 152328
rect 441528 152312 441580 152318
rect 441528 152254 441580 152260
rect 441724 152130 441752 152322
rect 441356 152102 441752 152130
rect 441908 149954 441936 152662
rect 442460 149954 442488 159462
rect 442724 152924 442776 152930
rect 442724 152866 442776 152872
rect 442736 151842 442764 152866
rect 442828 152658 442856 163200
rect 442908 153808 442960 153814
rect 442908 153750 442960 153756
rect 442816 152652 442868 152658
rect 442816 152594 442868 152600
rect 442920 151910 442948 153750
rect 442998 152960 443054 152969
rect 442998 152895 443000 152904
rect 443052 152895 443054 152904
rect 443000 152866 443052 152872
rect 443656 152250 443684 163200
rect 443828 152856 443880 152862
rect 443828 152798 443880 152804
rect 443184 152244 443236 152250
rect 443184 152186 443236 152192
rect 443644 152244 443696 152250
rect 443644 152186 443696 152192
rect 442908 151904 442960 151910
rect 442908 151846 442960 151852
rect 442724 151836 442776 151842
rect 442724 151778 442776 151784
rect 443196 149954 443224 152186
rect 443840 149954 443868 152798
rect 444484 152726 444512 163200
rect 445312 163146 445340 163200
rect 445404 163146 445432 163254
rect 445312 163118 445432 163146
rect 445024 159452 445076 159458
rect 445024 159394 445076 159400
rect 444472 152720 444524 152726
rect 444472 152662 444524 152668
rect 444472 152108 444524 152114
rect 444472 152050 444524 152056
rect 444484 149954 444512 152050
rect 445036 149954 445064 159394
rect 445680 152862 445708 163254
rect 446126 163200 446182 164400
rect 446954 163200 447010 164400
rect 447874 163200 447930 164400
rect 448702 163200 448758 164400
rect 449530 163200 449586 164400
rect 450358 163200 450414 164400
rect 451186 163200 451242 164400
rect 452014 163200 452070 164400
rect 452842 163200 452898 164400
rect 453762 163200 453818 164400
rect 454590 163200 454646 164400
rect 455418 163200 455474 164400
rect 456246 163200 456302 164400
rect 457074 163200 457130 164400
rect 457902 163200 457958 164400
rect 458730 163200 458786 164400
rect 459650 163200 459706 164400
rect 460478 163200 460534 164400
rect 461306 163200 461362 164400
rect 462134 163200 462190 164400
rect 462962 163200 463018 164400
rect 463790 163200 463846 164400
rect 464618 163200 464674 164400
rect 465538 163200 465594 164400
rect 466366 163200 466422 164400
rect 467194 163200 467250 164400
rect 468022 163200 468078 164400
rect 468850 163200 468906 164400
rect 469678 163200 469734 164400
rect 470506 163200 470562 164400
rect 471426 163200 471482 164400
rect 472254 163200 472310 164400
rect 473082 163200 473138 164400
rect 473910 163200 473966 164400
rect 474738 163200 474794 164400
rect 475566 163200 475622 164400
rect 476394 163200 476450 164400
rect 477314 163200 477370 164400
rect 478142 163200 478198 164400
rect 478970 163200 479026 164400
rect 479798 163200 479854 164400
rect 480626 163200 480682 164400
rect 481454 163200 481510 164400
rect 482282 163200 482338 164400
rect 483202 163200 483258 164400
rect 484030 163200 484086 164400
rect 484136 163254 484348 163282
rect 446140 159526 446168 163200
rect 446128 159520 446180 159526
rect 446128 159462 446180 159468
rect 446968 152930 446996 163200
rect 447888 159458 447916 163200
rect 447876 159452 447928 159458
rect 447876 159394 447928 159400
rect 448716 159390 448744 163200
rect 449544 159866 449572 163200
rect 449532 159860 449584 159866
rect 449532 159802 449584 159808
rect 450372 159730 450400 163200
rect 450360 159724 450412 159730
rect 450360 159666 450412 159672
rect 451200 159662 451228 163200
rect 451188 159656 451240 159662
rect 451188 159598 451240 159604
rect 452028 159594 452056 163200
rect 452016 159588 452068 159594
rect 452016 159530 452068 159536
rect 448704 159384 448756 159390
rect 448704 159326 448756 159332
rect 452856 158914 452884 163200
rect 453776 159798 453804 163200
rect 453764 159792 453816 159798
rect 453764 159734 453816 159740
rect 454604 159322 454632 163200
rect 455432 160070 455460 163200
rect 455420 160064 455472 160070
rect 455420 160006 455472 160012
rect 454592 159316 454644 159322
rect 454592 159258 454644 159264
rect 452844 158908 452896 158914
rect 452844 158850 452896 158856
rect 456260 158846 456288 163200
rect 456800 159520 456852 159526
rect 456800 159462 456852 159468
rect 456248 158840 456300 158846
rect 456248 158782 456300 158788
rect 456812 153202 456840 159462
rect 457088 159186 457116 163200
rect 457916 159254 457944 163200
rect 458744 159526 458772 163200
rect 459560 159860 459612 159866
rect 459560 159802 459612 159808
rect 458732 159520 458784 159526
rect 458732 159462 458784 159468
rect 457904 159248 457956 159254
rect 457904 159190 457956 159196
rect 457076 159180 457128 159186
rect 457076 159122 457128 159128
rect 452844 153196 452896 153202
rect 452844 153138 452896 153144
rect 456800 153196 456852 153202
rect 456800 153138 456852 153144
rect 459192 153196 459244 153202
rect 459192 153138 459244 153144
rect 448980 153128 449032 153134
rect 448980 153070 449032 153076
rect 447692 152992 447744 152998
rect 447692 152934 447744 152940
rect 445760 152924 445812 152930
rect 445760 152866 445812 152872
rect 446956 152924 447008 152930
rect 446956 152866 447008 152872
rect 445668 152856 445720 152862
rect 445668 152798 445720 152804
rect 445772 149954 445800 152866
rect 447140 152516 447192 152522
rect 447140 152458 447192 152464
rect 446404 152176 446456 152182
rect 446404 152118 446456 152124
rect 446416 149954 446444 152118
rect 447152 149954 447180 152458
rect 447704 149954 447732 152934
rect 448518 152416 448574 152425
rect 448518 152351 448574 152360
rect 448532 149954 448560 152351
rect 448992 149954 449020 153070
rect 449900 153060 449952 153066
rect 449900 153002 449952 153008
rect 449912 150226 449940 153002
rect 452200 152788 452252 152794
rect 452200 152730 452252 152736
rect 450268 152584 450320 152590
rect 450268 152526 450320 152532
rect 449912 150198 449986 150226
rect 440620 149926 440956 149954
rect 441264 149926 441600 149954
rect 441908 149926 442244 149954
rect 442460 149926 442888 149954
rect 443196 149926 443532 149954
rect 443840 149926 444176 149954
rect 444484 149926 444820 149954
rect 445036 149926 445464 149954
rect 445772 149926 446108 149954
rect 446416 149926 446752 149954
rect 447152 149926 447396 149954
rect 447704 149926 448040 149954
rect 448532 149926 448684 149954
rect 448992 149926 449328 149954
rect 449958 149940 449986 150198
rect 450280 149954 450308 152526
rect 451556 151972 451608 151978
rect 451556 151914 451608 151920
rect 450912 151904 450964 151910
rect 450912 151846 450964 151852
rect 450924 149954 450952 151846
rect 451568 149954 451596 151914
rect 452212 149954 452240 152730
rect 452856 149954 452884 153138
rect 458548 152856 458600 152862
rect 458548 152798 458600 152804
rect 458180 152720 458232 152726
rect 458180 152662 458232 152668
rect 456800 152652 456852 152658
rect 456800 152594 456852 152600
rect 453488 152448 453540 152454
rect 453488 152390 453540 152396
rect 453500 149954 453528 152390
rect 455420 152380 455472 152386
rect 455420 152322 455472 152328
rect 454776 152312 454828 152318
rect 454776 152254 454828 152260
rect 454224 152040 454276 152046
rect 454224 151982 454276 151988
rect 454236 149954 454264 151982
rect 454788 149954 454816 152254
rect 455432 149954 455460 152322
rect 456064 151836 456116 151842
rect 456064 151778 456116 151784
rect 456076 149954 456104 151778
rect 456812 149954 456840 152594
rect 457352 152244 457404 152250
rect 457352 152186 457404 152192
rect 457364 149954 457392 152186
rect 458192 150226 458220 152662
rect 458192 150198 458266 150226
rect 450280 149926 450616 149954
rect 450924 149926 451260 149954
rect 451568 149926 451904 149954
rect 452212 149926 452548 149954
rect 452856 149926 453192 149954
rect 453500 149926 453836 149954
rect 454236 149926 454480 149954
rect 454788 149926 455124 149954
rect 455432 149926 455768 149954
rect 456076 149926 456412 149954
rect 456812 149926 457056 149954
rect 457364 149926 457700 149954
rect 458238 149940 458266 150198
rect 458560 149954 458588 152798
rect 459204 149954 459232 153138
rect 459572 152046 459600 159802
rect 459664 159118 459692 163200
rect 460112 159452 460164 159458
rect 460112 159394 460164 159400
rect 459652 159112 459704 159118
rect 459652 159054 459704 159060
rect 459836 152924 459888 152930
rect 459836 152866 459888 152872
rect 459560 152040 459612 152046
rect 459560 151982 459612 151988
rect 459848 149954 459876 152866
rect 460124 151814 460152 159394
rect 460492 158982 460520 163200
rect 461320 159866 461348 163200
rect 461308 159860 461360 159866
rect 461308 159802 461360 159808
rect 461860 159656 461912 159662
rect 461860 159598 461912 159604
rect 461124 159384 461176 159390
rect 461124 159326 461176 159332
rect 460480 158976 460532 158982
rect 460480 158918 460532 158924
rect 460124 151786 460428 151814
rect 460400 149954 460428 151786
rect 461136 149954 461164 159326
rect 461872 153202 461900 159598
rect 462148 159458 462176 163200
rect 462228 159724 462280 159730
rect 462228 159666 462280 159672
rect 462136 159452 462188 159458
rect 462136 159394 462188 159400
rect 461860 153196 461912 153202
rect 461860 153138 461912 153144
rect 461768 152040 461820 152046
rect 461768 151982 461820 151988
rect 461780 149954 461808 151982
rect 462240 151814 462268 159666
rect 462976 159050 463004 163200
rect 463608 159588 463660 159594
rect 463608 159530 463660 159536
rect 462964 159044 463016 159050
rect 462964 158986 463016 158992
rect 463056 153196 463108 153202
rect 463056 153138 463108 153144
rect 462240 151786 462360 151814
rect 462332 149954 462360 151786
rect 463068 149954 463096 153138
rect 463620 151814 463648 159530
rect 463804 159390 463832 163200
rect 463792 159384 463844 159390
rect 463792 159326 463844 159332
rect 464252 158908 464304 158914
rect 464252 158850 464304 158856
rect 463620 151786 463740 151814
rect 463712 149954 463740 151786
rect 464264 149954 464292 158850
rect 464632 158778 464660 163200
rect 464988 159792 465040 159798
rect 464988 159734 465040 159740
rect 464620 158772 464672 158778
rect 464620 158714 464672 158720
rect 465000 151814 465028 159734
rect 465080 159520 465132 159526
rect 465080 159462 465132 159468
rect 465092 153066 465120 159462
rect 465552 159322 465580 163200
rect 465448 159316 465500 159322
rect 465448 159258 465500 159264
rect 465540 159316 465592 159322
rect 465540 159258 465592 159264
rect 465080 153060 465132 153066
rect 465080 153002 465132 153008
rect 465460 151814 465488 159258
rect 466380 158914 466408 163200
rect 466644 160064 466696 160070
rect 466644 160006 466696 160012
rect 466460 159112 466512 159118
rect 466460 159054 466512 159060
rect 466368 158908 466420 158914
rect 466368 158850 466420 158856
rect 466472 153202 466500 159054
rect 466552 158976 466604 158982
rect 466552 158918 466604 158924
rect 466460 153196 466512 153202
rect 466460 153138 466512 153144
rect 466564 153134 466592 158918
rect 466552 153128 466604 153134
rect 466552 153070 466604 153076
rect 465000 151786 465120 151814
rect 465460 151786 465580 151814
rect 465092 149954 465120 151786
rect 465552 149954 465580 151786
rect 466656 150226 466684 160006
rect 467208 160002 467236 163200
rect 468036 160070 468064 163200
rect 468024 160064 468076 160070
rect 468024 160006 468076 160012
rect 467196 159996 467248 160002
rect 467196 159938 467248 159944
rect 468024 159860 468076 159866
rect 468024 159802 468076 159808
rect 467840 159452 467892 159458
rect 467840 159394 467892 159400
rect 466828 158840 466880 158846
rect 466828 158782 466880 158788
rect 466610 150198 466684 150226
rect 458560 149926 458896 149954
rect 459204 149926 459540 149954
rect 459848 149926 460184 149954
rect 460400 149926 460828 149954
rect 461136 149926 461472 149954
rect 461780 149926 462116 149954
rect 462332 149926 462760 149954
rect 463068 149926 463404 149954
rect 463712 149926 464048 149954
rect 464264 149926 464692 149954
rect 465092 149926 465336 149954
rect 465552 149926 465980 149954
rect 466610 149940 466638 150198
rect 466840 149954 466868 158782
rect 467852 151842 467880 159394
rect 467932 159180 467984 159186
rect 467932 159122 467984 159128
rect 467840 151836 467892 151842
rect 467840 151778 467892 151784
rect 467944 150226 467972 159122
rect 468036 151910 468064 159802
rect 468864 159730 468892 163200
rect 468852 159724 468904 159730
rect 468852 159666 468904 159672
rect 469692 159526 469720 163200
rect 470520 159594 470548 163200
rect 471440 159798 471468 163200
rect 471428 159792 471480 159798
rect 471428 159734 471480 159740
rect 472268 159594 472296 163200
rect 470508 159588 470560 159594
rect 470508 159530 470560 159536
rect 472256 159588 472308 159594
rect 472256 159530 472308 159536
rect 469680 159520 469732 159526
rect 469680 159462 469732 159468
rect 471704 159384 471756 159390
rect 471704 159326 471756 159332
rect 468116 159248 468168 159254
rect 468116 159190 468168 159196
rect 468024 151904 468076 151910
rect 468024 151846 468076 151852
rect 467898 150198 467972 150226
rect 466840 149926 467268 149954
rect 467898 149940 467926 150198
rect 468128 149954 468156 159190
rect 469220 159044 469272 159050
rect 469220 158986 469272 158992
rect 468852 153060 468904 153066
rect 468852 153002 468904 153008
rect 468864 149954 468892 153002
rect 469232 151978 469260 158986
rect 471244 158772 471296 158778
rect 471244 158714 471296 158720
rect 471256 153202 471284 158714
rect 469496 153196 469548 153202
rect 469496 153138 469548 153144
rect 471244 153196 471296 153202
rect 471244 153138 471296 153144
rect 469220 151972 469272 151978
rect 469220 151914 469272 151920
rect 469508 149954 469536 153138
rect 471716 153134 471744 159326
rect 472256 159316 472308 159322
rect 472256 159258 472308 159264
rect 470140 153128 470192 153134
rect 470140 153070 470192 153076
rect 471704 153128 471756 153134
rect 471704 153070 471756 153076
rect 470152 149954 470180 153070
rect 472268 153066 472296 159258
rect 472348 158908 472400 158914
rect 472348 158850 472400 158856
rect 472256 153060 472308 153066
rect 472256 153002 472308 153008
rect 472360 152998 472388 158850
rect 473096 158778 473124 163200
rect 473360 159996 473412 160002
rect 473360 159938 473412 159944
rect 473084 158772 473136 158778
rect 473084 158714 473136 158720
rect 473372 153134 473400 159938
rect 473924 159050 473952 163200
rect 473912 159044 473964 159050
rect 473912 158986 473964 158992
rect 474752 158914 474780 163200
rect 474832 159724 474884 159730
rect 474832 159666 474884 159672
rect 474740 158908 474792 158914
rect 474740 158850 474792 158856
rect 474844 153202 474872 159666
rect 475580 158982 475608 163200
rect 476028 160064 476080 160070
rect 476028 160006 476080 160012
rect 475568 158976 475620 158982
rect 475568 158918 475620 158924
rect 473544 153196 473596 153202
rect 473544 153138 473596 153144
rect 474832 153196 474884 153202
rect 474832 153138 474884 153144
rect 472716 153128 472768 153134
rect 472716 153070 472768 153076
rect 473360 153128 473412 153134
rect 473360 153070 473412 153076
rect 472348 152992 472400 152998
rect 472348 152934 472400 152940
rect 472072 151972 472124 151978
rect 472072 151914 472124 151920
rect 470784 151904 470836 151910
rect 470784 151846 470836 151852
rect 470796 149954 470824 151846
rect 471428 151836 471480 151842
rect 471428 151778 471480 151784
rect 471440 149954 471468 151778
rect 472084 149954 472112 151914
rect 472728 149954 472756 153070
rect 473556 149954 473584 153138
rect 475292 153128 475344 153134
rect 475292 153070 475344 153076
rect 474004 153060 474056 153066
rect 474004 153002 474056 153008
rect 474016 149954 474044 153002
rect 474740 152992 474792 152998
rect 474740 152934 474792 152940
rect 474752 149954 474780 152934
rect 475304 149954 475332 153070
rect 476040 151814 476068 160006
rect 476120 159656 476172 159662
rect 476120 159598 476172 159604
rect 476132 153134 476160 159598
rect 476408 158846 476436 163200
rect 477328 159458 477356 163200
rect 478156 159526 478184 163200
rect 478984 159866 479012 163200
rect 478972 159860 479024 159866
rect 478972 159802 479024 159808
rect 478420 159792 478472 159798
rect 478420 159734 478472 159740
rect 477408 159520 477460 159526
rect 477408 159462 477460 159468
rect 478144 159520 478196 159526
rect 478144 159462 478196 159468
rect 477316 159452 477368 159458
rect 477316 159394 477368 159400
rect 476396 158840 476448 158846
rect 476396 158782 476448 158788
rect 476580 153196 476632 153202
rect 476580 153138 476632 153144
rect 476120 153128 476172 153134
rect 476120 153070 476172 153076
rect 476040 151786 476160 151814
rect 476132 149954 476160 151786
rect 476592 149954 476620 153138
rect 477420 151814 477448 159462
rect 477868 153128 477920 153134
rect 477868 153070 477920 153076
rect 477420 151786 477540 151814
rect 477512 150226 477540 151786
rect 477512 150198 477586 150226
rect 468128 149926 468556 149954
rect 468864 149926 469200 149954
rect 469508 149926 469844 149954
rect 470152 149926 470488 149954
rect 470796 149926 471132 149954
rect 471440 149926 471776 149954
rect 472084 149926 472420 149954
rect 472728 149926 473064 149954
rect 473556 149926 473708 149954
rect 474016 149926 474352 149954
rect 474752 149926 474996 149954
rect 475304 149926 475640 149954
rect 476132 149926 476284 149954
rect 476592 149926 476928 149954
rect 477558 149940 477586 150198
rect 477880 149954 477908 153070
rect 478432 149954 478460 159734
rect 479812 159594 479840 163200
rect 480640 159934 480668 163200
rect 480628 159928 480680 159934
rect 480628 159870 480680 159876
rect 479064 159588 479116 159594
rect 479064 159530 479116 159536
rect 479800 159588 479852 159594
rect 479800 159530 479852 159536
rect 479076 149954 479104 159530
rect 480260 159044 480312 159050
rect 480260 158986 480312 158992
rect 479708 158772 479760 158778
rect 479708 158714 479760 158720
rect 479720 149954 479748 158714
rect 480272 151814 480300 158986
rect 480996 158908 481048 158914
rect 480996 158850 481048 158856
rect 480272 151786 480392 151814
rect 480364 149954 480392 151786
rect 481008 149954 481036 158850
rect 481468 158778 481496 163200
rect 482296 159662 482324 163200
rect 482284 159656 482336 159662
rect 482284 159598 482336 159604
rect 481732 158976 481784 158982
rect 481732 158918 481784 158924
rect 481456 158772 481508 158778
rect 481456 158714 481508 158720
rect 481744 149954 481772 158918
rect 482376 158840 482428 158846
rect 482376 158782 482428 158788
rect 482388 149954 482416 158782
rect 483216 152998 483244 163200
rect 484044 163146 484072 163200
rect 484136 163146 484164 163254
rect 484044 163118 484164 163146
rect 483664 159520 483716 159526
rect 483664 159462 483716 159468
rect 483296 159452 483348 159458
rect 483296 159394 483348 159400
rect 483204 152992 483256 152998
rect 483204 152934 483256 152940
rect 483308 150226 483336 159394
rect 483308 150198 483382 150226
rect 477880 149926 478216 149954
rect 478432 149926 478860 149954
rect 479076 149926 479504 149954
rect 479720 149926 480148 149954
rect 480364 149926 480792 149954
rect 481008 149926 481436 149954
rect 481744 149926 482080 149954
rect 482388 149926 482724 149954
rect 483354 149940 483382 150198
rect 483676 149954 483704 159462
rect 484320 153134 484348 163254
rect 484858 163200 484914 164400
rect 485686 163200 485742 164400
rect 486514 163200 486570 164400
rect 487342 163200 487398 164400
rect 488170 163200 488226 164400
rect 488276 163254 488488 163282
rect 484584 159860 484636 159866
rect 484584 159802 484636 159808
rect 484308 153128 484360 153134
rect 484308 153070 484360 153076
rect 484596 150226 484624 159802
rect 484768 159588 484820 159594
rect 484768 159530 484820 159536
rect 484780 151814 484808 159530
rect 484872 153066 484900 163200
rect 485700 153202 485728 163200
rect 485872 159928 485924 159934
rect 485872 159870 485924 159876
rect 485688 153196 485740 153202
rect 485688 153138 485740 153144
rect 484860 153060 484912 153066
rect 484860 153002 484912 153008
rect 484780 151786 484900 151814
rect 484596 150198 484670 150226
rect 483676 149926 484012 149954
rect 484642 149940 484670 150198
rect 484872 149954 484900 151786
rect 485884 150226 485912 159870
rect 486148 158772 486200 158778
rect 486148 158714 486200 158720
rect 485884 150198 485958 150226
rect 484872 149926 485300 149954
rect 485930 149940 485958 150198
rect 486160 149954 486188 158714
rect 486528 152046 486556 163200
rect 486516 152040 486568 152046
rect 486516 151982 486568 151988
rect 487356 151978 487384 163200
rect 488184 163146 488212 163200
rect 488276 163146 488304 163254
rect 488184 163118 488304 163146
rect 487436 159656 487488 159662
rect 487436 159598 487488 159604
rect 487344 151972 487396 151978
rect 487344 151914 487396 151920
rect 487448 149954 487476 159598
rect 488172 153128 488224 153134
rect 488172 153070 488224 153076
rect 487528 152992 487580 152998
rect 487528 152934 487580 152940
rect 486160 149926 486588 149954
rect 487232 149926 487476 149954
rect 487540 149954 487568 152934
rect 488184 149954 488212 153070
rect 488460 151842 488488 163254
rect 489090 163200 489146 164400
rect 489918 163200 489974 164400
rect 490746 163200 490802 164400
rect 491574 163200 491630 164400
rect 492402 163200 492458 164400
rect 493230 163200 493286 164400
rect 494058 163200 494114 164400
rect 494978 163200 495034 164400
rect 495084 163254 495296 163282
rect 488724 153060 488776 153066
rect 488724 153002 488776 153008
rect 488448 151836 488500 151842
rect 488448 151778 488500 151784
rect 488736 149954 488764 153002
rect 489104 151910 489132 163200
rect 489368 153196 489420 153202
rect 489368 153138 489420 153144
rect 489092 151904 489144 151910
rect 489092 151846 489144 151852
rect 489380 149954 489408 153138
rect 489932 153134 489960 163200
rect 489920 153128 489972 153134
rect 489920 153070 489972 153076
rect 490760 152998 490788 163200
rect 490748 152992 490800 152998
rect 490748 152934 490800 152940
rect 491588 152862 491616 163200
rect 492416 153202 492444 163200
rect 492404 153196 492456 153202
rect 492404 153138 492456 153144
rect 493244 153134 493272 163200
rect 492772 153128 492824 153134
rect 492772 153070 492824 153076
rect 493232 153128 493284 153134
rect 493232 153070 493284 153076
rect 491576 152856 491628 152862
rect 491576 152798 491628 152804
rect 490012 152040 490064 152046
rect 490012 151982 490064 151988
rect 490024 149954 490052 151982
rect 490656 151972 490708 151978
rect 490656 151914 490708 151920
rect 490668 149954 490696 151914
rect 491944 151904 491996 151910
rect 491944 151846 491996 151852
rect 491300 151836 491352 151842
rect 491300 151778 491352 151784
rect 491312 149954 491340 151778
rect 491956 149954 491984 151846
rect 492784 149954 492812 153070
rect 494072 152998 494100 163200
rect 494992 163146 495020 163200
rect 495084 163146 495112 163254
rect 494992 163118 495112 163146
rect 495268 153202 495296 163254
rect 495806 163200 495862 164400
rect 496634 163200 496690 164400
rect 497462 163200 497518 164400
rect 498290 163200 498346 164400
rect 499118 163200 499174 164400
rect 499224 163254 499528 163282
rect 494520 153196 494572 153202
rect 494520 153138 494572 153144
rect 495256 153196 495308 153202
rect 495256 153138 495308 153144
rect 493232 152992 493284 152998
rect 493232 152934 493284 152940
rect 494060 152992 494112 152998
rect 494060 152934 494112 152940
rect 493244 149954 493272 152934
rect 494060 152856 494112 152862
rect 494060 152798 494112 152804
rect 494072 149954 494100 152798
rect 494532 149954 494560 153138
rect 495820 153134 495848 163200
rect 496648 153202 496676 163200
rect 496452 153196 496504 153202
rect 496452 153138 496504 153144
rect 496636 153196 496688 153202
rect 496636 153138 496688 153144
rect 495440 153128 495492 153134
rect 495440 153070 495492 153076
rect 495808 153128 495860 153134
rect 495808 153070 495860 153076
rect 495452 150226 495480 153070
rect 495808 152992 495860 152998
rect 495808 152934 495860 152940
rect 495452 150198 495526 150226
rect 487540 149926 487876 149954
rect 488184 149926 488520 149954
rect 488736 149926 489072 149954
rect 489380 149926 489716 149954
rect 490024 149926 490360 149954
rect 490668 149926 491004 149954
rect 491312 149926 491648 149954
rect 491956 149926 492292 149954
rect 492784 149926 492936 149954
rect 493244 149926 493580 149954
rect 494072 149926 494224 149954
rect 494532 149926 494868 149954
rect 495498 149940 495526 150198
rect 495820 149954 495848 152934
rect 496464 149954 496492 153138
rect 497096 153128 497148 153134
rect 497096 153070 497148 153076
rect 497108 149954 497136 153070
rect 497476 153066 497504 163200
rect 498304 153202 498332 163200
rect 499132 163146 499160 163200
rect 499224 163146 499252 163254
rect 499132 163118 499252 163146
rect 497740 153196 497792 153202
rect 497740 153138 497792 153144
rect 498292 153196 498344 153202
rect 498292 153138 498344 153144
rect 499028 153196 499080 153202
rect 499028 153138 499080 153144
rect 497464 153060 497516 153066
rect 497464 153002 497516 153008
rect 497752 149954 497780 153138
rect 498292 153060 498344 153066
rect 498292 153002 498344 153008
rect 498304 149954 498332 153002
rect 499040 149954 499068 153138
rect 499500 151858 499528 163254
rect 499946 163200 500002 164400
rect 500052 163254 500264 163282
rect 499960 163146 499988 163200
rect 500052 163146 500080 163254
rect 499960 163118 500080 163146
rect 499500 151830 499620 151858
rect 499592 149954 499620 151830
rect 500236 149954 500264 163254
rect 500866 163200 500922 164400
rect 500972 163254 501644 163282
rect 500880 151814 500908 163200
rect 500972 153202 501000 163254
rect 501616 163146 501644 163254
rect 501694 163200 501750 164400
rect 502522 163200 502578 164400
rect 503350 163200 503406 164400
rect 503732 163254 504128 163282
rect 501708 163146 501736 163200
rect 501616 163118 501736 163146
rect 500960 153196 501012 153202
rect 500960 153138 501012 153144
rect 501604 153196 501656 153202
rect 501604 153138 501656 153144
rect 500880 151786 501000 151814
rect 500972 149954 501000 151786
rect 501616 149954 501644 153138
rect 502536 150226 502564 163200
rect 503364 152998 503392 163200
rect 502892 152992 502944 152998
rect 502892 152934 502944 152940
rect 503352 152992 503404 152998
rect 503352 152934 503404 152940
rect 502536 150198 502610 150226
rect 495820 149926 496156 149954
rect 496464 149926 496800 149954
rect 497108 149926 497444 149954
rect 497752 149926 498088 149954
rect 498304 149926 498732 149954
rect 499040 149926 499376 149954
rect 499592 149926 500020 149954
rect 500236 149926 500664 149954
rect 500972 149926 501308 149954
rect 501616 149926 501952 149954
rect 502582 149940 502610 150198
rect 502904 149954 502932 152934
rect 503732 149954 503760 163254
rect 504100 163146 504128 163254
rect 504178 163200 504234 164400
rect 505006 163200 505062 164400
rect 505112 163254 505784 163282
rect 504192 163146 504220 163200
rect 504100 163118 504220 163146
rect 505020 158778 505048 163200
rect 504088 158772 504140 158778
rect 504088 158714 504140 158720
rect 505008 158772 505060 158778
rect 505008 158714 505060 158720
rect 504100 149954 504128 158714
rect 505112 150226 505140 163254
rect 505756 163146 505784 163254
rect 505834 163200 505890 164400
rect 506754 163200 506810 164400
rect 507582 163200 507638 164400
rect 508410 163200 508466 164400
rect 509238 163200 509294 164400
rect 510066 163200 510122 164400
rect 510894 163200 510950 164400
rect 511722 163200 511778 164400
rect 512012 163254 512592 163282
rect 505848 163146 505876 163200
rect 505756 163118 505876 163146
rect 506388 158840 506440 158846
rect 506388 158782 506440 158788
rect 506204 158772 506256 158778
rect 506204 158714 506256 158720
rect 505112 150198 505186 150226
rect 502904 149926 503240 149954
rect 503732 149926 503884 149954
rect 504100 149926 504528 149954
rect 505158 149940 505186 150198
rect 506216 149954 506244 158714
rect 506400 150226 506428 158782
rect 506768 158778 506796 163200
rect 507596 158846 507624 163200
rect 507584 158840 507636 158846
rect 507584 158782 507636 158788
rect 508424 158778 508452 163200
rect 508688 158908 508740 158914
rect 508688 158850 508740 158856
rect 506756 158772 506808 158778
rect 506756 158714 506808 158720
rect 507492 158772 507544 158778
rect 507492 158714 507544 158720
rect 508412 158772 508464 158778
rect 508412 158714 508464 158720
rect 506400 150198 506474 150226
rect 505816 149926 506244 149954
rect 506446 149940 506474 150198
rect 507504 149954 507532 158714
rect 507768 151972 507820 151978
rect 507768 151914 507820 151920
rect 507780 150226 507808 151914
rect 507104 149926 507532 149954
rect 507734 150198 507808 150226
rect 507734 149940 507762 150198
rect 508700 149954 508728 158850
rect 509252 151978 509280 163200
rect 510080 158914 510108 163200
rect 510068 158908 510120 158914
rect 510068 158850 510120 158856
rect 509976 158772 510028 158778
rect 509976 158714 510028 158720
rect 509240 151972 509292 151978
rect 509240 151914 509292 151920
rect 509056 151836 509108 151842
rect 509056 151778 509108 151784
rect 509068 150226 509096 151778
rect 508392 149926 508728 149954
rect 509022 150198 509096 150226
rect 509022 149940 509050 150198
rect 509988 149954 510016 158714
rect 510436 153196 510488 153202
rect 510436 153138 510488 153144
rect 510448 149954 510476 153138
rect 510908 151842 510936 163200
rect 511736 158778 511764 163200
rect 511724 158772 511776 158778
rect 511724 158714 511776 158720
rect 512012 153202 512040 163254
rect 512564 163146 512592 163254
rect 512642 163200 512698 164400
rect 513470 163200 513526 164400
rect 514298 163200 514354 164400
rect 514864 163254 515076 163282
rect 512656 163146 512684 163200
rect 512564 163118 512684 163146
rect 512000 153196 512052 153202
rect 512000 153138 512052 153144
rect 512552 153196 512604 153202
rect 512552 153138 512604 153144
rect 511264 153128 511316 153134
rect 511264 153070 511316 153076
rect 510896 151836 510948 151842
rect 510896 151778 510948 151784
rect 511276 149954 511304 153070
rect 511724 153060 511776 153066
rect 511724 153002 511776 153008
rect 511736 149954 511764 153002
rect 512564 149954 512592 153138
rect 513484 153134 513512 163200
rect 513472 153128 513524 153134
rect 513472 153070 513524 153076
rect 514312 153066 514340 163200
rect 514864 153202 514892 163254
rect 515048 163146 515076 163254
rect 515126 163200 515182 164400
rect 515954 163200 516010 164400
rect 516152 163254 516732 163282
rect 515140 163146 515168 163200
rect 515048 163118 515168 163146
rect 515128 158772 515180 158778
rect 515128 158714 515180 158720
rect 514852 153196 514904 153202
rect 514852 153138 514904 153144
rect 514300 153060 514352 153066
rect 514300 153002 514352 153008
rect 513196 152992 513248 152998
rect 513196 152934 513248 152940
rect 513208 149954 513236 152934
rect 513840 152924 513892 152930
rect 513840 152866 513892 152872
rect 513852 149954 513880 152866
rect 514484 152448 514536 152454
rect 514484 152390 514536 152396
rect 514496 149954 514524 152390
rect 515140 149954 515168 158714
rect 515968 152998 515996 163200
rect 515956 152992 516008 152998
rect 515956 152934 516008 152940
rect 516152 152930 516180 163254
rect 516704 163146 516732 163254
rect 516782 163200 516838 164400
rect 517610 163200 517666 164400
rect 518530 163200 518586 164400
rect 518912 163254 519308 163282
rect 516796 163146 516824 163200
rect 516704 163118 516824 163146
rect 517624 161474 517652 163200
rect 517532 161446 517652 161474
rect 517532 158794 517560 161446
rect 518348 159520 518400 159526
rect 518348 159462 518400 159468
rect 517440 158766 517560 158794
rect 516140 152924 516192 152930
rect 516140 152866 516192 152872
rect 517440 152454 517468 158766
rect 517428 152448 517480 152454
rect 517428 152390 517480 152396
rect 515772 152108 515824 152114
rect 515772 152050 515824 152056
rect 515784 149954 515812 152050
rect 515956 152040 516008 152046
rect 515956 151982 516008 151988
rect 509680 149926 510016 149954
rect 510324 149926 510476 149954
rect 510968 149926 511304 149954
rect 511612 149926 511764 149954
rect 512256 149926 512592 149954
rect 512900 149926 513236 149954
rect 513544 149926 513880 149954
rect 514188 149926 514524 149954
rect 514832 149926 515168 149954
rect 515476 149926 515812 149954
rect 515968 149954 515996 151982
rect 517428 151972 517480 151978
rect 517428 151914 517480 151920
rect 517060 151836 517112 151842
rect 517060 151778 517112 151784
rect 517072 149954 517100 151778
rect 517440 150226 517468 151914
rect 515968 149926 516120 149954
rect 516764 149926 517100 149954
rect 517394 150198 517468 150226
rect 517394 149940 517422 150198
rect 518360 149954 518388 159462
rect 518544 158778 518572 163200
rect 518716 159384 518768 159390
rect 518716 159326 518768 159332
rect 518532 158772 518584 158778
rect 518532 158714 518584 158720
rect 518728 150226 518756 159326
rect 518912 152114 518940 163254
rect 519280 163146 519308 163254
rect 519358 163200 519414 164400
rect 519464 163254 520136 163282
rect 519372 163146 519400 163200
rect 519280 163118 519400 163146
rect 518900 152108 518952 152114
rect 518900 152050 518952 152056
rect 519464 152046 519492 163254
rect 519726 163160 519782 163169
rect 520108 163146 520136 163254
rect 520186 163200 520242 164400
rect 520292 163254 520964 163282
rect 520200 163146 520228 163200
rect 520108 163118 520228 163146
rect 519726 163095 519782 163104
rect 519542 161664 519598 161673
rect 519542 161599 519598 161608
rect 519452 152040 519504 152046
rect 519452 151982 519504 151988
rect 518052 149926 518388 149954
rect 518682 150198 518756 150226
rect 518682 149940 518710 150198
rect 519556 147937 519584 161599
rect 519634 160168 519690 160177
rect 519634 160103 519690 160112
rect 519542 147928 519598 147937
rect 519542 147863 519598 147872
rect 519648 146577 519676 160103
rect 519740 149297 519768 163095
rect 520186 158672 520242 158681
rect 520186 158607 520242 158616
rect 520002 157176 520058 157185
rect 520002 157111 520058 157120
rect 519818 151056 519874 151065
rect 519818 150991 519874 151000
rect 519726 149288 519782 149297
rect 519726 149223 519782 149232
rect 519726 148064 519782 148073
rect 519726 147999 519782 148008
rect 519634 146568 519690 146577
rect 519634 146503 519690 146512
rect 519542 143440 519598 143449
rect 519542 143375 519598 143384
rect 519358 141944 519414 141953
rect 519358 141879 519414 141888
rect 117240 132518 117360 132546
rect 117332 132410 117360 132518
rect 117240 132382 117360 132410
rect 117240 127945 117268 132382
rect 519372 130257 519400 141879
rect 519556 131617 519584 143375
rect 519740 135697 519768 147999
rect 519832 138417 519860 150991
rect 519910 149560 519966 149569
rect 519910 149495 519966 149504
rect 519818 138408 519874 138417
rect 519818 138343 519874 138352
rect 519924 137057 519952 149495
rect 520016 143857 520044 157111
rect 520094 154048 520150 154057
rect 520094 153983 520150 153992
rect 520002 143848 520058 143857
rect 520002 143783 520058 143792
rect 520108 141137 520136 153983
rect 520200 145217 520228 158607
rect 520292 151842 520320 163254
rect 520936 163146 520964 163254
rect 521014 163200 521070 164400
rect 521842 163200 521898 164400
rect 522670 163200 522726 164400
rect 523498 163200 523554 164400
rect 521028 163146 521056 163200
rect 520936 163118 521056 163146
rect 521856 161474 521884 163200
rect 521672 161446 521884 161474
rect 521672 158794 521700 161446
rect 522684 159526 522712 163200
rect 522672 159520 522724 159526
rect 522672 159462 522724 159468
rect 523512 159390 523540 163200
rect 523500 159384 523552 159390
rect 523500 159326 523552 159332
rect 521580 158766 521700 158794
rect 521198 155680 521254 155689
rect 521198 155615 521254 155624
rect 521106 152552 521162 152561
rect 521106 152487 521162 152496
rect 520280 151836 520332 151842
rect 520280 151778 520332 151784
rect 520922 146568 520978 146577
rect 520922 146503 520978 146512
rect 520186 145208 520242 145217
rect 520186 145143 520242 145152
rect 520094 141128 520150 141137
rect 520094 141063 520150 141072
rect 520186 140448 520242 140457
rect 520186 140383 520242 140392
rect 520002 138952 520058 138961
rect 520002 138887 520058 138896
rect 519910 137048 519966 137057
rect 519910 136983 519966 136992
rect 519910 135824 519966 135833
rect 519910 135759 519966 135768
rect 519726 135688 519782 135697
rect 519726 135623 519782 135632
rect 519818 134328 519874 134337
rect 519818 134263 519874 134272
rect 519634 132832 519690 132841
rect 519634 132767 519690 132776
rect 519542 131608 519598 131617
rect 519542 131543 519598 131552
rect 519358 130248 519414 130257
rect 519358 130183 519414 130192
rect 519542 129840 519598 129849
rect 519542 129775 519598 129784
rect 117226 127936 117282 127945
rect 117226 127871 117282 127880
rect 519450 126712 519506 126721
rect 519450 126647 519506 126656
rect 519358 120592 519414 120601
rect 519358 120527 519414 120536
rect 519372 111217 519400 120527
rect 519464 116657 519492 126647
rect 519556 119377 519584 129775
rect 519648 122097 519676 132767
rect 519726 131336 519782 131345
rect 519726 131271 519782 131280
rect 519634 122088 519690 122097
rect 519634 122023 519690 122032
rect 519740 120737 519768 131271
rect 519832 123457 519860 134263
rect 519924 124817 519952 135759
rect 520016 127537 520044 138887
rect 520094 137456 520150 137465
rect 520094 137391 520150 137400
rect 520002 127528 520058 127537
rect 520002 127463 520058 127472
rect 520108 126177 520136 137391
rect 520200 128897 520228 140383
rect 520936 134473 520964 146503
rect 521014 144936 521070 144945
rect 521014 144871 521070 144880
rect 520922 134464 520978 134473
rect 520922 134399 520978 134408
rect 521028 132977 521056 144871
rect 521120 139777 521148 152487
rect 521212 142497 521240 155615
rect 521580 151978 521608 158766
rect 521568 151972 521620 151978
rect 521568 151914 521620 151920
rect 521198 142488 521254 142497
rect 521198 142423 521254 142432
rect 521106 139768 521162 139777
rect 521106 139703 521162 139712
rect 521014 132968 521070 132977
rect 521014 132903 521070 132912
rect 520186 128888 520242 128897
rect 520186 128823 520242 128832
rect 520186 128344 520242 128353
rect 520186 128279 520242 128288
rect 520094 126168 520150 126177
rect 520094 126103 520150 126112
rect 520094 125216 520150 125225
rect 520094 125151 520150 125160
rect 519910 124808 519966 124817
rect 519910 124743 519966 124752
rect 520002 123720 520058 123729
rect 520002 123655 520058 123664
rect 519818 123448 519874 123457
rect 519818 123383 519874 123392
rect 519818 122224 519874 122233
rect 519818 122159 519874 122168
rect 519726 120728 519782 120737
rect 519726 120663 519782 120672
rect 519542 119368 519598 119377
rect 519542 119303 519598 119312
rect 519726 119232 519782 119241
rect 519726 119167 519782 119176
rect 519542 117600 519598 117609
rect 519542 117535 519598 117544
rect 519450 116648 519506 116657
rect 519450 116583 519506 116592
rect 519358 111208 519414 111217
rect 519358 111143 519414 111152
rect 519556 108497 519584 117535
rect 519634 114608 519690 114617
rect 519634 114543 519690 114552
rect 519542 108488 519598 108497
rect 519542 108423 519598 108432
rect 519648 105777 519676 114543
rect 519740 109857 519768 119167
rect 519832 112577 519860 122159
rect 519910 116104 519966 116113
rect 519910 116039 519966 116048
rect 519818 112568 519874 112577
rect 519818 112503 519874 112512
rect 519726 109848 519782 109857
rect 519726 109783 519782 109792
rect 519924 107137 519952 116039
rect 520016 113937 520044 123655
rect 520108 115297 520136 125151
rect 520200 118017 520228 128279
rect 520186 118008 520242 118017
rect 520186 117943 520242 117952
rect 520094 115288 520150 115297
rect 520094 115223 520150 115232
rect 520002 113928 520058 113937
rect 520002 113863 520058 113872
rect 520370 113112 520426 113121
rect 520370 113047 520426 113056
rect 519910 107128 519966 107137
rect 519910 107063 519966 107072
rect 519634 105768 519690 105777
rect 519634 105703 519690 105712
rect 520278 105496 520334 105505
rect 520278 105431 520334 105440
rect 117134 104816 117190 104825
rect 117134 104751 117190 104760
rect 117042 101008 117098 101017
rect 117042 100943 117098 100952
rect 519634 99376 519690 99385
rect 519634 99311 519690 99320
rect 116858 99104 116914 99113
rect 116858 99039 116914 99048
rect 116766 97200 116822 97209
rect 116766 97135 116822 97144
rect 519266 96384 519322 96393
rect 519266 96319 519322 96328
rect 116674 95296 116730 95305
rect 116674 95231 116730 95240
rect 116582 93392 116638 93401
rect 116582 93327 116638 93336
rect 116124 92472 116176 92478
rect 116124 92414 116176 92420
rect 116136 91361 116164 92414
rect 116122 91352 116178 91361
rect 116122 91287 116178 91296
rect 116124 89684 116176 89690
rect 116124 89626 116176 89632
rect 116136 89457 116164 89626
rect 519280 89457 519308 96319
rect 519648 92177 519676 99311
rect 519726 97880 519782 97889
rect 519726 97815 519782 97824
rect 519634 92168 519690 92177
rect 519634 92103 519690 92112
rect 519740 90817 519768 97815
rect 520292 97617 520320 105431
rect 520384 104417 520412 113047
rect 521566 111616 521622 111625
rect 521566 111551 521622 111560
rect 521474 110120 521530 110129
rect 521474 110055 521530 110064
rect 521106 108488 521162 108497
rect 521106 108423 521162 108432
rect 520370 104408 520426 104417
rect 520370 104343 520426 104352
rect 520922 104000 520978 104009
rect 520922 103935 520978 103944
rect 520278 97608 520334 97617
rect 520278 97543 520334 97552
rect 520936 96257 520964 103935
rect 521014 102504 521070 102513
rect 521014 102439 521070 102448
rect 520922 96248 520978 96257
rect 520922 96183 520978 96192
rect 521028 95033 521056 102439
rect 521120 100337 521148 108423
rect 521382 106992 521438 107001
rect 521382 106927 521438 106936
rect 521198 101008 521254 101017
rect 521198 100943 521254 100952
rect 521106 100328 521162 100337
rect 521106 100263 521162 100272
rect 521014 95024 521070 95033
rect 521014 94959 521070 94968
rect 520002 94888 520058 94897
rect 520002 94823 520058 94832
rect 519726 90808 519782 90817
rect 519726 90743 519782 90752
rect 116122 89448 116178 89457
rect 116122 89383 116178 89392
rect 519266 89448 519322 89457
rect 519266 89383 519322 89392
rect 116032 88324 116084 88330
rect 116032 88266 116084 88272
rect 116044 87553 116072 88266
rect 520016 88097 520044 94823
rect 521212 93537 521240 100943
rect 521396 98977 521424 106927
rect 521488 101697 521516 110055
rect 521580 103057 521608 111551
rect 521566 103048 521622 103057
rect 521566 102983 521622 102992
rect 521474 101688 521530 101697
rect 521474 101623 521530 101632
rect 521382 98968 521438 98977
rect 521382 98903 521438 98912
rect 521198 93528 521254 93537
rect 521198 93463 521254 93472
rect 520186 93392 520242 93401
rect 520186 93327 520242 93336
rect 520002 88088 520058 88097
rect 520002 88023 520058 88032
rect 116030 87544 116086 87553
rect 116030 87479 116086 87488
rect 520200 86737 520228 93327
rect 521290 91896 521346 91905
rect 521290 91831 521346 91840
rect 520922 90264 520978 90273
rect 520922 90199 520978 90208
rect 520186 86728 520242 86737
rect 520186 86663 520242 86672
rect 520278 85776 520334 85785
rect 520278 85711 520334 85720
rect 115202 85640 115258 85649
rect 115202 85575 115258 85584
rect 116584 83972 116636 83978
rect 116584 83914 116636 83920
rect 116596 83745 116624 83914
rect 116582 83736 116638 83745
rect 116582 83671 116638 83680
rect 116216 82816 116268 82822
rect 116216 82758 116268 82764
rect 520002 82784 520058 82793
rect 116228 81841 116256 82758
rect 520002 82719 520058 82728
rect 116214 81832 116270 81841
rect 116214 81767 116270 81776
rect 115940 80028 115992 80034
rect 115940 79970 115992 79976
rect 115952 79937 115980 79970
rect 115938 79928 115994 79937
rect 115938 79863 115994 79872
rect 519634 79656 519690 79665
rect 519634 79591 519690 79600
rect 114192 78668 114244 78674
rect 114192 78610 114244 78616
rect 116124 78668 116176 78674
rect 116124 78610 116176 78616
rect 116136 78033 116164 78610
rect 116122 78024 116178 78033
rect 116122 77959 116178 77968
rect 116674 74080 116730 74089
rect 116674 74015 116730 74024
rect 116582 72176 116638 72185
rect 116582 72111 116638 72120
rect 116596 71806 116624 72111
rect 114192 71800 114244 71806
rect 114192 71742 114244 71748
rect 116584 71800 116636 71806
rect 116584 71742 116636 71748
rect 114100 69080 114152 69086
rect 114100 69022 114152 69028
rect 114008 67652 114060 67658
rect 114008 67594 114060 67600
rect 113916 66292 113968 66298
rect 113916 66234 113968 66240
rect 113364 64728 113416 64734
rect 113364 64670 113416 64676
rect 113376 64569 113404 64670
rect 113362 64560 113418 64569
rect 113362 64495 113418 64504
rect 113824 63572 113876 63578
rect 113824 63514 113876 63520
rect 112444 62144 112496 62150
rect 112444 62086 112496 62092
rect 110326 58032 110382 58041
rect 109696 57990 110326 58018
rect 109696 41154 109724 57990
rect 110326 57967 110382 57976
rect 110326 56808 110382 56817
rect 110326 56743 110382 56752
rect 110340 55214 110368 56743
rect 109788 55186 110368 55214
rect 109788 41290 109816 55186
rect 110326 53952 110382 53961
rect 109880 53910 110326 53938
rect 109880 42106 109908 53910
rect 110326 53887 110382 53896
rect 110326 52592 110382 52601
rect 110326 52527 110382 52536
rect 110340 51218 110368 52527
rect 110340 51190 110460 51218
rect 110326 51096 110382 51105
rect 109972 51054 110326 51082
rect 109972 42378 110000 51054
rect 110326 51031 110382 51040
rect 110432 50946 110460 51190
rect 110064 50918 110460 50946
rect 110064 42650 110092 50918
rect 110326 48376 110382 48385
rect 110156 48334 110326 48362
rect 110156 42922 110184 48334
rect 110326 48311 110382 48320
rect 110326 47152 110382 47161
rect 110326 47087 110382 47096
rect 110340 45554 110368 47087
rect 110340 45526 110828 45554
rect 110326 42936 110382 42945
rect 110156 42894 110326 42922
rect 110326 42871 110382 42880
rect 110064 42622 110552 42650
rect 110326 42392 110382 42401
rect 109972 42350 110326 42378
rect 110326 42327 110382 42336
rect 109880 42078 110460 42106
rect 109788 41262 110000 41290
rect 109696 41126 109908 41154
rect 109880 40610 109908 41126
rect 109420 40582 109908 40610
rect 109420 40034 109448 40582
rect 109972 40474 110000 41262
rect 109788 40446 110000 40474
rect 109788 40034 109816 40446
rect 109420 40006 109632 40034
rect 109788 40006 110368 40034
rect 109604 34762 109632 40006
rect 110340 34898 110368 40006
rect 110432 35057 110460 42078
rect 110418 35048 110474 35057
rect 110418 34983 110474 34992
rect 110340 34870 110460 34898
rect 110326 34776 110382 34785
rect 109604 34734 110326 34762
rect 110326 34711 110382 34720
rect 110326 34640 110382 34649
rect 109604 34598 110326 34626
rect 109604 28994 109632 34598
rect 110326 34575 110382 34584
rect 110432 34514 110460 34870
rect 110340 34486 110460 34514
rect 110340 29481 110368 34486
rect 110524 29730 110552 42622
rect 110694 42392 110750 42401
rect 110694 42327 110750 42336
rect 110602 41440 110658 41449
rect 110602 41375 110658 41384
rect 110616 34649 110644 41375
rect 110602 34640 110658 34649
rect 110602 34575 110658 34584
rect 110708 29889 110736 42327
rect 110694 29880 110750 29889
rect 110694 29815 110750 29824
rect 110800 29730 110828 45526
rect 111062 44296 111118 44305
rect 111062 44231 111118 44240
rect 110878 42936 110934 42945
rect 110878 42871 110934 42880
rect 110432 29702 110552 29730
rect 110616 29702 110828 29730
rect 110326 29472 110382 29481
rect 110326 29407 110382 29416
rect 110326 29336 110382 29345
rect 109880 29294 110326 29322
rect 109880 28994 109908 29294
rect 110326 29271 110382 29280
rect 110326 29200 110382 29209
rect 109512 28966 109632 28994
rect 109696 28966 109908 28994
rect 110156 29158 110326 29186
rect 110156 28994 110184 29158
rect 110326 29135 110382 29144
rect 110156 28966 110276 28994
rect 109512 28642 109540 28966
rect 109696 28914 109724 28966
rect 109696 28886 110000 28914
rect 109972 28642 110000 28886
rect 109512 28614 109908 28642
rect 109972 28614 110184 28642
rect 109880 23474 109908 28614
rect 109604 23446 109908 23474
rect 109604 22094 109632 23446
rect 110156 22094 110184 28614
rect 109420 22066 109632 22094
rect 109788 22066 110184 22094
rect 109420 12434 109448 22066
rect 109788 20714 109816 22066
rect 110248 20714 110276 28966
rect 109696 20686 109816 20714
rect 109880 20686 110276 20714
rect 109420 12406 109632 12434
rect 33046 2680 33102 2689
rect 33046 2615 33102 2624
rect 42062 2680 42118 2689
rect 42706 2680 42762 2689
rect 42642 2638 42706 2666
rect 42062 2615 42118 2624
rect 42706 2615 42762 2624
rect 44730 2680 44786 2689
rect 44730 2615 44786 2624
rect 58990 2680 59046 2689
rect 58990 2615 59046 2624
rect 59174 2680 59230 2689
rect 62762 2680 62818 2689
rect 62698 2638 62762 2666
rect 59174 2615 59230 2624
rect 62762 2615 62818 2624
rect 63038 2680 63094 2689
rect 63038 2615 63094 2624
rect 64602 2680 64658 2689
rect 64602 2615 64658 2624
rect 66994 2680 67050 2689
rect 66994 2615 67050 2624
rect 76562 2680 76618 2689
rect 76562 2615 76618 2624
rect 89166 2680 89222 2689
rect 89166 2615 89222 2624
rect 89718 2680 89774 2689
rect 89718 2615 89774 2624
rect 89902 2680 89958 2689
rect 89902 2615 89958 2624
rect 90362 2680 90418 2689
rect 90362 2615 90418 2624
rect 92478 2680 92534 2689
rect 92754 2680 92810 2689
rect 92690 2638 92754 2666
rect 92478 2615 92534 2624
rect 92754 2615 92810 2624
rect 95146 2680 95202 2689
rect 95146 2615 95202 2624
rect 95330 2680 95386 2689
rect 95330 2615 95386 2624
rect 96434 2680 96490 2689
rect 96434 2615 96490 2624
rect 99930 2680 99986 2689
rect 99930 2615 99986 2624
rect 100850 2680 100906 2689
rect 100850 2615 100906 2624
rect 101770 2680 101826 2689
rect 101770 2615 101826 2624
rect 101954 2680 102010 2689
rect 101954 2615 102010 2624
rect 102782 2680 102838 2689
rect 102782 2615 102838 2624
rect 29550 2544 29606 2553
rect 29302 2502 29550 2530
rect 29550 2479 29606 2488
rect 26054 2408 26110 2417
rect 25990 2366 26054 2394
rect 26054 2343 26110 2352
rect 22926 2272 22982 2281
rect 22678 2230 22926 2258
rect 22926 2207 22982 2216
rect 19614 2136 19670 2145
rect 2700 1358 2728 2108
rect 6012 1873 6040 2108
rect 5998 1864 6054 1873
rect 5998 1799 6054 1808
rect 9324 1601 9352 2108
rect 12636 1737 12664 2108
rect 15962 2094 16252 2122
rect 19366 2094 19614 2122
rect 16224 2009 16252 2094
rect 19614 2071 19670 2080
rect 16210 2000 16266 2009
rect 16210 1935 16266 1944
rect 12622 1728 12678 1737
rect 12622 1663 12678 1672
rect 9310 1592 9366 1601
rect 9310 1527 9366 1536
rect 32692 1426 32720 2108
rect 32680 1420 32732 1426
rect 32680 1362 32732 1368
rect 2688 1352 2740 1358
rect 2688 1294 2740 1300
rect 32784 870 32904 898
rect 32784 800 32812 870
rect 32770 -400 32826 800
rect 32876 762 32904 870
rect 33060 762 33088 2615
rect 36004 1290 36032 2108
rect 35992 1284 36044 1290
rect 35992 1226 36044 1232
rect 39316 1222 39344 2108
rect 42076 1902 42104 2615
rect 44744 1902 44772 2615
rect 42064 1896 42116 1902
rect 42064 1838 42116 1844
rect 44732 1896 44784 1902
rect 44732 1838 44784 1844
rect 46032 1494 46060 2108
rect 46020 1488 46072 1494
rect 46020 1430 46072 1436
rect 39304 1216 39356 1222
rect 39304 1158 39356 1164
rect 49344 1154 49372 2108
rect 49332 1148 49384 1154
rect 49332 1090 49384 1096
rect 52656 1086 52684 2108
rect 55968 1465 55996 2108
rect 59004 1902 59032 2615
rect 58992 1896 59044 1902
rect 58992 1838 59044 1844
rect 59188 1834 59216 2615
rect 59176 1828 59228 1834
rect 59176 1770 59228 1776
rect 59372 1766 59400 2108
rect 63052 1834 63080 2615
rect 63040 1828 63092 1834
rect 63040 1770 63092 1776
rect 59360 1760 59412 1766
rect 59360 1702 59412 1708
rect 64616 1494 64644 2615
rect 64604 1488 64656 1494
rect 55954 1456 56010 1465
rect 64604 1430 64656 1436
rect 55954 1391 56010 1400
rect 52644 1080 52696 1086
rect 52644 1022 52696 1028
rect 65996 1018 66024 2108
rect 67008 1902 67036 2615
rect 66996 1896 67048 1902
rect 66996 1838 67048 1844
rect 69308 1630 69336 2108
rect 69296 1624 69348 1630
rect 69296 1566 69348 1572
rect 72712 1494 72740 2108
rect 72700 1488 72752 1494
rect 72700 1430 72752 1436
rect 65984 1012 66036 1018
rect 65984 954 66036 960
rect 76024 950 76052 2108
rect 76576 1766 76604 2615
rect 76564 1760 76616 1766
rect 76564 1702 76616 1708
rect 79336 1562 79364 2108
rect 82648 1698 82676 2108
rect 86052 1766 86080 2108
rect 86040 1760 86092 1766
rect 86040 1702 86092 1708
rect 82636 1692 82688 1698
rect 82636 1634 82688 1640
rect 79324 1556 79376 1562
rect 79324 1498 79376 1504
rect 89180 1193 89208 2615
rect 89364 1834 89392 2108
rect 89352 1828 89404 1834
rect 89352 1770 89404 1776
rect 89166 1184 89222 1193
rect 89166 1119 89222 1128
rect 76012 944 76064 950
rect 76012 886 76064 892
rect 89732 882 89760 2615
rect 89916 1329 89944 2615
rect 90376 1902 90404 2615
rect 90364 1896 90416 1902
rect 92492 1884 92520 2615
rect 92572 1896 92624 1902
rect 92492 1856 92572 1884
rect 90364 1838 90416 1844
rect 92572 1838 92624 1844
rect 89902 1320 89958 1329
rect 89902 1255 89958 1264
rect 95160 1193 95188 2615
rect 95344 1902 95372 2615
rect 95332 1896 95384 1902
rect 95332 1838 95384 1844
rect 95146 1184 95202 1193
rect 95146 1119 95202 1128
rect 95988 882 96016 2108
rect 96448 1329 96476 2615
rect 99406 2094 99880 2122
rect 99852 1714 99880 2094
rect 99944 1902 99972 2615
rect 99932 1896 99984 1902
rect 99932 1838 99984 1844
rect 100024 1896 100076 1902
rect 100024 1838 100076 1844
rect 100036 1714 100064 1838
rect 99852 1686 100064 1714
rect 96434 1320 96490 1329
rect 96434 1255 96490 1264
rect 98274 1320 98330 1329
rect 98274 1255 98330 1264
rect 89720 876 89772 882
rect 89720 818 89772 824
rect 95976 876 96028 882
rect 95976 818 96028 824
rect 98288 800 98316 1255
rect 100864 882 100892 2615
rect 101784 1630 101812 2615
rect 101772 1624 101824 1630
rect 101772 1566 101824 1572
rect 101968 1329 101996 2615
rect 102704 1902 102732 2108
rect 102692 1896 102744 1902
rect 102692 1838 102744 1844
rect 101954 1320 102010 1329
rect 101954 1255 102010 1264
rect 101404 1012 101456 1018
rect 101404 954 101456 960
rect 101416 882 101444 954
rect 100852 876 100904 882
rect 100852 818 100904 824
rect 101404 876 101456 882
rect 101404 818 101456 824
rect 102796 814 102824 2615
rect 105912 1896 105964 1902
rect 105912 1838 105964 1844
rect 103980 1692 104032 1698
rect 103980 1634 104032 1640
rect 103992 1562 104020 1634
rect 105924 1630 105952 1838
rect 106016 1630 106044 2108
rect 109132 1896 109184 1902
rect 109184 1844 109264 1850
rect 109132 1838 109264 1844
rect 109144 1822 109264 1838
rect 109328 1834 109356 2108
rect 109236 1698 109264 1822
rect 109316 1828 109368 1834
rect 109316 1770 109368 1776
rect 109224 1692 109276 1698
rect 109224 1634 109276 1640
rect 105912 1624 105964 1630
rect 105912 1566 105964 1572
rect 106004 1624 106056 1630
rect 106004 1566 106056 1572
rect 109040 1624 109092 1630
rect 109092 1572 109264 1578
rect 109040 1566 109264 1572
rect 103980 1556 104032 1562
rect 109052 1550 109264 1566
rect 103980 1498 104032 1504
rect 109236 1426 109264 1550
rect 109604 1494 109632 12406
rect 109696 11914 109724 20686
rect 109880 19334 109908 20686
rect 110326 20224 110382 20233
rect 110326 20159 110382 20168
rect 110340 19334 110368 20159
rect 109788 19306 109908 19334
rect 109972 19306 110368 19334
rect 109788 12186 109816 19306
rect 109972 16574 110000 19306
rect 109880 16546 110000 16574
rect 109880 12458 109908 16546
rect 110326 12472 110382 12481
rect 109880 12430 110326 12458
rect 110326 12407 110382 12416
rect 110326 12200 110382 12209
rect 109788 12158 110326 12186
rect 110326 12135 110382 12144
rect 109696 11886 110368 11914
rect 110340 9194 110368 11886
rect 110432 9602 110460 29702
rect 110510 29608 110566 29617
rect 110510 29543 110566 29552
rect 110524 9761 110552 29543
rect 110616 20097 110644 29702
rect 110892 29594 110920 42871
rect 110970 35048 111026 35057
rect 110970 34983 111026 34992
rect 110708 29566 110920 29594
rect 110602 20088 110658 20097
rect 110602 20023 110658 20032
rect 110602 12200 110658 12209
rect 110602 12135 110658 12144
rect 110510 9752 110566 9761
rect 110510 9687 110566 9696
rect 110432 9574 110552 9602
rect 110340 9166 110460 9194
rect 110326 9072 110382 9081
rect 110326 9007 110382 9016
rect 110340 8922 110368 9007
rect 109696 8894 110368 8922
rect 109696 1902 109724 8894
rect 110326 8800 110382 8809
rect 110248 8758 110326 8786
rect 110248 8650 110276 8758
rect 110326 8735 110382 8744
rect 109788 8622 110276 8650
rect 109788 1902 109816 8622
rect 110326 8528 110382 8537
rect 110248 8486 110326 8514
rect 110248 8106 110276 8486
rect 110326 8463 110382 8472
rect 110326 8392 110382 8401
rect 110326 8327 110382 8336
rect 109880 8078 110276 8106
rect 109880 3233 109908 8078
rect 110340 7698 110368 8327
rect 110432 7857 110460 9166
rect 110418 7848 110474 7857
rect 110418 7783 110474 7792
rect 109972 7670 110368 7698
rect 109866 3224 109922 3233
rect 109866 3159 109922 3168
rect 109866 2952 109922 2961
rect 109866 2887 109922 2896
rect 109880 1902 109908 2887
rect 109684 1896 109736 1902
rect 109684 1838 109736 1844
rect 109776 1896 109828 1902
rect 109776 1838 109828 1844
rect 109868 1896 109920 1902
rect 109868 1838 109920 1844
rect 109972 1766 110000 7670
rect 110524 7562 110552 9574
rect 110616 9081 110644 12135
rect 110602 9072 110658 9081
rect 110602 9007 110658 9016
rect 110248 7534 110552 7562
rect 110248 7290 110276 7534
rect 110064 7262 110276 7290
rect 110064 3913 110092 7262
rect 110708 7018 110736 29566
rect 110786 29472 110842 29481
rect 110786 29407 110842 29416
rect 110800 20233 110828 29407
rect 110984 24854 111012 34983
rect 111076 29617 111104 44231
rect 111246 34776 111302 34785
rect 111246 34711 111302 34720
rect 111154 34640 111210 34649
rect 111154 34575 111210 34584
rect 111062 29608 111118 29617
rect 111062 29543 111118 29552
rect 111168 29345 111196 34575
rect 111154 29336 111210 29345
rect 111154 29271 111210 29280
rect 111260 29209 111288 34711
rect 111338 29880 111394 29889
rect 111338 29815 111394 29824
rect 111246 29200 111302 29209
rect 111246 29135 111302 29144
rect 110892 24826 111012 24854
rect 110786 20224 110842 20233
rect 110786 20159 110842 20168
rect 110786 20088 110842 20097
rect 110786 20023 110842 20032
rect 110156 6990 110736 7018
rect 110050 3904 110106 3913
rect 110050 3839 110106 3848
rect 109960 1760 110012 1766
rect 109960 1702 110012 1708
rect 110052 1760 110104 1766
rect 110052 1702 110104 1708
rect 109592 1488 109644 1494
rect 109592 1430 109644 1436
rect 110064 1426 110092 1702
rect 110156 1630 110184 6990
rect 110800 6882 110828 20023
rect 110892 15194 110920 24826
rect 110892 15166 111104 15194
rect 110970 12472 111026 12481
rect 110970 12407 111026 12416
rect 110878 9752 110934 9761
rect 110878 9687 110934 9696
rect 110248 6854 110828 6882
rect 110144 1624 110196 1630
rect 110144 1566 110196 1572
rect 110248 1562 110276 6854
rect 110892 5681 110920 9687
rect 110984 8809 111012 12407
rect 110970 8800 111026 8809
rect 110970 8735 111026 8744
rect 111076 8537 111104 15166
rect 111062 8528 111118 8537
rect 111062 8463 111118 8472
rect 111352 8401 111380 29815
rect 111338 8392 111394 8401
rect 111338 8327 111394 8336
rect 110970 7848 111026 7857
rect 110970 7783 111026 7792
rect 110878 5672 110934 5681
rect 110878 5607 110934 5616
rect 110326 5548 110382 5557
rect 110326 5483 110382 5492
rect 110340 3074 110368 5483
rect 110694 4176 110750 4185
rect 110694 4111 110750 4120
rect 110340 3046 110644 3074
rect 110326 2952 110382 2961
rect 110326 2887 110382 2896
rect 110340 1873 110368 2887
rect 110326 1864 110382 1873
rect 110326 1799 110382 1808
rect 110616 1698 110644 3046
rect 110708 2961 110736 4111
rect 110984 3641 111012 7783
rect 110970 3632 111026 3641
rect 110970 3567 111026 3576
rect 110694 2952 110750 2961
rect 110694 2887 110750 2896
rect 111708 2848 111760 2854
rect 111706 2816 111708 2825
rect 111760 2816 111762 2825
rect 111706 2751 111762 2760
rect 112456 1834 112484 62086
rect 112536 42832 112588 42838
rect 112536 42774 112588 42780
rect 112444 1828 112496 1834
rect 112444 1770 112496 1776
rect 110604 1692 110656 1698
rect 110604 1634 110656 1640
rect 110236 1556 110288 1562
rect 110236 1498 110288 1504
rect 109132 1420 109184 1426
rect 109132 1362 109184 1368
rect 109224 1420 109276 1426
rect 109224 1362 109276 1368
rect 110052 1420 110104 1426
rect 110052 1362 110104 1368
rect 109144 1306 109172 1362
rect 109408 1352 109460 1358
rect 109144 1300 109408 1306
rect 109144 1294 109460 1300
rect 109144 1278 109448 1294
rect 109040 1216 109092 1222
rect 109040 1158 109092 1164
rect 109052 814 109080 1158
rect 112548 950 112576 42774
rect 113836 7721 113864 63514
rect 113928 19009 113956 66234
rect 114020 30433 114048 67594
rect 114112 41857 114140 69022
rect 114204 53145 114232 71742
rect 116306 70272 116362 70281
rect 116306 70207 116362 70216
rect 116320 69086 116348 70207
rect 116308 69080 116360 69086
rect 116308 69022 116360 69028
rect 116122 68368 116178 68377
rect 116122 68303 116178 68312
rect 116136 67658 116164 68303
rect 116124 67652 116176 67658
rect 116124 67594 116176 67600
rect 116582 66464 116638 66473
rect 116582 66399 116638 66408
rect 116596 66298 116624 66399
rect 116584 66292 116636 66298
rect 116584 66234 116636 66240
rect 116688 64874 116716 74015
rect 519266 73672 519322 73681
rect 519266 73607 519322 73616
rect 519280 67833 519308 73607
rect 519648 73273 519676 79591
rect 519726 78160 519782 78169
rect 519726 78095 519782 78104
rect 519634 73264 519690 73273
rect 519634 73199 519690 73208
rect 519740 72457 519768 78095
rect 520016 75993 520044 82719
rect 520186 81152 520242 81161
rect 520186 81087 520242 81096
rect 520094 76664 520150 76673
rect 520094 76599 520150 76608
rect 520002 75984 520058 75993
rect 520002 75919 520058 75928
rect 520002 75168 520058 75177
rect 520002 75103 520058 75112
rect 519726 72448 519782 72457
rect 519726 72383 519782 72392
rect 519450 72040 519506 72049
rect 519450 71975 519506 71984
rect 519266 67824 519322 67833
rect 519266 67759 519322 67768
rect 519266 67552 519322 67561
rect 519266 67487 519322 67496
rect 116596 64846 116716 64874
rect 116596 64734 116624 64846
rect 116584 64728 116636 64734
rect 116584 64670 116636 64676
rect 116214 64560 116270 64569
rect 116214 64495 116270 64504
rect 116228 63578 116256 64495
rect 116216 63572 116268 63578
rect 116216 63514 116268 63520
rect 116122 62656 116178 62665
rect 116122 62591 116178 62600
rect 116136 62150 116164 62591
rect 116124 62144 116176 62150
rect 116124 62086 116176 62092
rect 519280 61033 519308 67487
rect 519464 66473 519492 71975
rect 520016 69193 520044 75103
rect 520108 70553 520136 76599
rect 520200 74633 520228 81087
rect 520292 78577 520320 85711
rect 520936 82657 520964 90199
rect 521014 87272 521070 87281
rect 521014 87207 521070 87216
rect 520922 82648 520978 82657
rect 520922 82583 520978 82592
rect 521028 79937 521056 87207
rect 521198 84280 521254 84289
rect 521198 84215 521254 84224
rect 521014 79928 521070 79937
rect 521014 79863 521070 79872
rect 520278 78568 520334 78577
rect 520278 78503 520334 78512
rect 521212 77217 521240 84215
rect 521304 84017 521332 91831
rect 521382 88768 521438 88777
rect 521382 88703 521438 88712
rect 521290 84008 521346 84017
rect 521290 83943 521346 83952
rect 521396 81297 521424 88703
rect 521382 81288 521438 81297
rect 521382 81223 521438 81232
rect 521198 77208 521254 77217
rect 521198 77143 521254 77152
rect 520186 74624 520242 74633
rect 520186 74559 520242 74568
rect 520094 70544 520150 70553
rect 520094 70479 520150 70488
rect 520186 70408 520242 70417
rect 520186 70343 520242 70352
rect 520002 69184 520058 69193
rect 520002 69119 520058 69128
rect 519634 69048 519690 69057
rect 519634 68983 519690 68992
rect 519450 66464 519506 66473
rect 519450 66399 519506 66408
rect 519648 63753 519676 68983
rect 519818 66056 519874 66065
rect 519818 65991 519874 66000
rect 519634 63744 519690 63753
rect 519634 63679 519690 63688
rect 519266 61024 519322 61033
rect 519266 60959 519322 60968
rect 116582 60616 116638 60625
rect 116582 60551 116638 60560
rect 114190 53136 114246 53145
rect 114190 53071 114246 53080
rect 116122 43344 116178 43353
rect 116122 43279 116178 43288
rect 116136 42838 116164 43279
rect 116124 42832 116176 42838
rect 116124 42774 116176 42780
rect 114098 41848 114154 41857
rect 114098 41783 114154 41792
rect 114006 30424 114062 30433
rect 114006 30359 114062 30368
rect 116398 26072 116454 26081
rect 116398 26007 116454 26016
rect 116306 20360 116362 20369
rect 116306 20295 116362 20304
rect 113914 19000 113970 19009
rect 113914 18935 113970 18944
rect 116214 18456 116270 18465
rect 116214 18391 116270 18400
rect 116030 16416 116086 16425
rect 116030 16351 116086 16360
rect 115938 12608 115994 12617
rect 115938 12543 115994 12552
rect 113822 7712 113878 7721
rect 113822 7647 113878 7656
rect 115952 2145 115980 12543
rect 116044 2417 116072 16351
rect 116122 14512 116178 14521
rect 116122 14447 116178 14456
rect 116030 2408 116086 2417
rect 116030 2343 116086 2352
rect 116136 2281 116164 14447
rect 116228 2553 116256 18391
rect 116320 7562 116348 20295
rect 116412 7682 116440 26007
rect 116490 22264 116546 22273
rect 116490 22199 116546 22208
rect 116400 7676 116452 7682
rect 116400 7618 116452 7624
rect 116320 7534 116440 7562
rect 116308 7472 116360 7478
rect 116308 7414 116360 7420
rect 116320 3369 116348 7414
rect 116306 3360 116362 3369
rect 116306 3295 116362 3304
rect 116306 3088 116362 3097
rect 116306 3023 116362 3032
rect 116214 2544 116270 2553
rect 116214 2479 116270 2488
rect 116122 2272 116178 2281
rect 116122 2207 116178 2216
rect 115938 2136 115994 2145
rect 115938 2071 115994 2080
rect 116320 1290 116348 3023
rect 116412 1426 116440 7534
rect 116400 1420 116452 1426
rect 116400 1362 116452 1368
rect 116308 1284 116360 1290
rect 116308 1226 116360 1232
rect 116504 1222 116532 22199
rect 116596 1766 116624 60551
rect 519832 59673 519860 65991
rect 520200 65113 520228 70343
rect 520186 65104 520242 65113
rect 520186 65039 520242 65048
rect 521106 64560 521162 64569
rect 521106 64495 521162 64504
rect 520738 62928 520794 62937
rect 520738 62863 520794 62872
rect 520278 61432 520334 61441
rect 520278 61367 520334 61376
rect 519818 59664 519874 59673
rect 519818 59599 519874 59608
rect 520186 56944 520242 56953
rect 520292 56930 520320 61367
rect 520752 58313 520780 62863
rect 521120 62393 521148 64495
rect 521106 62384 521162 62393
rect 521106 62319 521162 62328
rect 521014 59936 521070 59945
rect 521014 59871 521070 59880
rect 520738 58304 520794 58313
rect 520738 58239 520794 58248
rect 520242 56902 520320 56930
rect 520370 56944 520426 56953
rect 520186 56879 520242 56888
rect 520370 56879 520426 56888
rect 520278 55448 520334 55457
rect 520278 55383 520334 55392
rect 519266 53816 519322 53825
rect 519266 53751 519322 53760
rect 519280 50153 519308 53751
rect 520094 52320 520150 52329
rect 520094 52255 520150 52264
rect 520002 50824 520058 50833
rect 520002 50759 520058 50768
rect 519266 50144 519322 50153
rect 519266 50079 519322 50088
rect 519450 47832 519506 47841
rect 519450 47767 519506 47776
rect 519464 44713 519492 47767
rect 520016 47433 520044 50759
rect 520108 48793 520136 52255
rect 520292 51513 520320 55383
rect 520384 52873 520412 56879
rect 521028 55593 521056 59871
rect 521106 58440 521162 58449
rect 521106 58375 521162 58384
rect 521014 55584 521070 55593
rect 521014 55519 521070 55528
rect 521120 54233 521148 58375
rect 521106 54224 521162 54233
rect 521106 54159 521162 54168
rect 520370 52864 520426 52873
rect 520370 52799 520426 52808
rect 520278 51504 520334 51513
rect 520278 51439 520334 51448
rect 520186 49328 520242 49337
rect 520186 49263 520242 49272
rect 520094 48784 520150 48793
rect 520094 48719 520150 48728
rect 520002 47424 520058 47433
rect 520002 47359 520058 47368
rect 519910 46336 519966 46345
rect 519910 46271 519966 46280
rect 519450 44704 519506 44713
rect 519450 44639 519506 44648
rect 519818 44704 519874 44713
rect 519818 44639 519874 44648
rect 519832 41993 519860 44639
rect 519924 43353 519952 46271
rect 520200 46073 520228 49263
rect 520186 46064 520242 46073
rect 520186 45999 520242 46008
rect 519910 43344 519966 43353
rect 519910 43279 519966 43288
rect 520186 43208 520242 43217
rect 520186 43143 520242 43152
rect 519818 41984 519874 41993
rect 519818 41919 519874 41928
rect 520094 41712 520150 41721
rect 520094 41647 520150 41656
rect 116766 39536 116822 39545
rect 116766 39471 116822 39480
rect 116674 37632 116730 37641
rect 116674 37567 116730 37576
rect 116584 1760 116636 1766
rect 116584 1702 116636 1708
rect 116492 1216 116544 1222
rect 116492 1158 116544 1164
rect 112536 944 112588 950
rect 112536 886 112588 892
rect 116688 882 116716 37567
rect 116780 3233 116808 39471
rect 520108 39273 520136 41647
rect 520200 40633 520228 43143
rect 520186 40624 520242 40633
rect 520186 40559 520242 40568
rect 520186 40216 520242 40225
rect 520186 40151 520242 40160
rect 520094 39264 520150 39273
rect 520094 39199 520150 39208
rect 519818 38720 519874 38729
rect 519818 38655 519874 38664
rect 519832 36553 519860 38655
rect 520200 37913 520228 40151
rect 520186 37904 520242 37913
rect 520186 37839 520242 37848
rect 521566 37224 521622 37233
rect 521566 37159 521622 37168
rect 519818 36544 519874 36553
rect 519818 36479 519874 36488
rect 521580 36009 521608 37159
rect 521566 36000 521622 36009
rect 521566 35935 521622 35944
rect 521106 35592 521162 35601
rect 521106 35527 521162 35536
rect 521120 34513 521148 35527
rect 521106 34504 521162 34513
rect 521106 34439 521162 34448
rect 520922 34096 520978 34105
rect 520922 34031 520978 34040
rect 116950 33824 117006 33833
rect 116950 33759 117006 33768
rect 116858 31784 116914 31793
rect 116858 31719 116914 31728
rect 116766 3224 116822 3233
rect 116766 3159 116822 3168
rect 116872 1018 116900 31719
rect 116964 3777 116992 33759
rect 520936 33153 520964 34031
rect 520922 33144 520978 33153
rect 520922 33079 520978 33088
rect 520922 32600 520978 32609
rect 520922 32535 520978 32544
rect 520936 31657 520964 32535
rect 520922 31648 520978 31657
rect 520922 31583 520978 31592
rect 520922 31104 520978 31113
rect 520922 31039 520978 31048
rect 520936 30297 520964 31039
rect 520922 30288 520978 30297
rect 520922 30223 520978 30232
rect 117042 29880 117098 29889
rect 117042 29815 117098 29824
rect 116950 3768 117006 3777
rect 116950 3703 117006 3712
rect 117056 1154 117084 29815
rect 521106 29608 521162 29617
rect 521106 29543 521162 29552
rect 521120 28393 521148 29543
rect 521106 28384 521162 28393
rect 521106 28319 521162 28328
rect 117134 27976 117190 27985
rect 117134 27911 117190 27920
rect 117148 3505 117176 27911
rect 117226 24168 117282 24177
rect 117226 24103 117282 24112
rect 117134 3496 117190 3505
rect 117134 3431 117190 3440
rect 117044 1148 117096 1154
rect 117044 1090 117096 1096
rect 116860 1012 116912 1018
rect 116860 954 116912 960
rect 116676 876 116728 882
rect 116676 818 116728 824
rect 117240 814 117268 24103
rect 521106 21992 521162 22001
rect 521106 21927 521162 21936
rect 521120 20913 521148 21927
rect 521106 20904 521162 20913
rect 521106 20839 521162 20848
rect 520738 20496 520794 20505
rect 520738 20431 520794 20440
rect 520752 19553 520780 20431
rect 520738 19544 520794 19553
rect 520738 19479 520794 19488
rect 520922 19000 520978 19009
rect 520922 18935 520978 18944
rect 520936 18193 520964 18935
rect 520922 18184 520978 18193
rect 520922 18119 520978 18128
rect 521106 9344 521162 9353
rect 521106 9279 521162 9288
rect 521120 8265 521148 9279
rect 521106 8256 521162 8265
rect 521106 8191 521162 8200
rect 520370 7984 520426 7993
rect 520370 7919 520426 7928
rect 520384 6769 520412 7919
rect 520370 6760 520426 6769
rect 520370 6695 520426 6704
rect 521106 6624 521162 6633
rect 521106 6559 521162 6568
rect 521120 5273 521148 6559
rect 520922 5264 520978 5273
rect 520922 5199 520978 5208
rect 521106 5264 521162 5273
rect 521106 5199 521162 5208
rect 520936 3777 520964 5199
rect 521014 3904 521070 3913
rect 521014 3839 521070 3848
rect 520922 3768 520978 3777
rect 520922 3703 520978 3712
rect 143644 2514 143980 2530
rect 443656 2514 443992 2530
rect 143632 2508 143980 2514
rect 143684 2502 143980 2508
rect 425796 2508 425848 2514
rect 143632 2450 143684 2456
rect 425796 2450 425848 2456
rect 443644 2508 443992 2514
rect 443696 2502 443992 2508
rect 443644 2450 443696 2456
rect 193600 2094 193936 2122
rect 243648 2094 243984 2122
rect 293604 2094 293940 2122
rect 343652 2094 343988 2122
rect 393608 2094 393944 2122
rect 163778 1592 163834 1601
rect 163778 1527 163834 1536
rect 102784 808 102836 814
rect 32876 734 33088 762
rect 98274 -400 98330 800
rect 102784 750 102836 756
rect 109040 808 109092 814
rect 109040 750 109092 756
rect 117228 808 117280 814
rect 163792 800 163820 1527
rect 193600 1494 193628 2094
rect 229282 1728 229338 1737
rect 229282 1663 229338 1672
rect 193588 1488 193640 1494
rect 193588 1430 193640 1436
rect 229296 800 229324 1663
rect 243648 1601 243676 2094
rect 293604 1737 293632 2094
rect 293590 1728 293646 1737
rect 293590 1663 293646 1672
rect 243634 1592 243690 1601
rect 243634 1527 243690 1536
rect 294786 1456 294842 1465
rect 343652 1426 343680 2094
rect 393608 1465 393636 2094
rect 360290 1456 360346 1465
rect 294786 1391 294788 1400
rect 294840 1391 294842 1400
rect 343640 1420 343692 1426
rect 294788 1362 294840 1368
rect 360290 1391 360346 1400
rect 393594 1456 393650 1465
rect 393594 1391 393650 1400
rect 343640 1362 343692 1368
rect 294800 800 294828 1362
rect 360304 800 360332 1391
rect 425808 800 425836 2450
rect 521028 2281 521056 3839
rect 521106 2680 521162 2689
rect 521106 2615 521162 2624
rect 521014 2272 521070 2281
rect 521014 2207 521070 2216
rect 493612 2094 493948 2122
rect 493612 1426 493640 2094
rect 491300 1420 491352 1426
rect 491300 1362 491352 1368
rect 493600 1420 493652 1426
rect 493600 1362 493652 1368
rect 491312 800 491340 1362
rect 117228 750 117280 756
rect 163778 -400 163834 800
rect 229282 -400 229338 800
rect 294786 -400 294842 800
rect 360290 -400 360346 800
rect 425794 -400 425850 800
rect 491298 -400 491354 800
rect 521120 785 521148 2615
rect 521106 776 521162 785
rect 521106 711 521162 720
<< via2 >>
rect 3974 153720 4030 153776
rect 16302 159296 16358 159352
rect 17130 153992 17186 154048
rect 20534 153856 20590 153912
rect 23018 159432 23074 159488
rect 28078 156576 28134 156632
rect 29826 159568 29882 159624
rect 31482 156712 31538 156768
rect 30654 154128 30710 154184
rect 12990 152496 13046 152552
rect 9586 152360 9642 152416
rect 6090 150592 6146 150648
rect 2686 150456 2742 150512
rect 33966 157936 34022 157992
rect 40682 158072 40738 158128
rect 44086 158208 44142 158264
rect 57518 158344 57574 158400
rect 55862 156848 55918 156904
rect 55034 154264 55090 154320
rect 62578 155488 62634 155544
rect 65982 155216 66038 155272
rect 72698 156984 72754 157040
rect 76010 155760 76066 155816
rect 78586 155624 78642 155680
rect 68466 155352 68522 155408
rect 85302 155896 85358 155952
rect 86130 154400 86186 154456
rect 104622 158480 104678 158536
rect 82818 149640 82874 149696
rect 109590 148008 109646 148064
rect 115570 157120 115626 157176
rect 111062 150456 111118 150512
rect 110970 147328 111026 147384
rect 110326 146376 110382 146432
rect 110326 106256 110382 106312
rect 111338 150592 111394 150648
rect 111706 147328 111762 147384
rect 113822 144200 113878 144256
rect 116122 145152 116178 145208
rect 116030 143248 116086 143304
rect 115294 141344 115350 141400
rect 116122 139440 116178 139496
rect 116122 137536 116178 137592
rect 115202 135496 115258 135552
rect 116030 133592 116086 133648
rect 114190 132776 114246 132832
rect 113914 121352 113970 121408
rect 114006 110064 114062 110120
rect 114098 98640 114154 98696
rect 114190 87216 114246 87272
rect 116122 131688 116178 131744
rect 116582 149640 116638 149696
rect 116490 129784 116546 129840
rect 116122 125976 116178 126032
rect 116122 124108 116124 124128
rect 116124 124108 116176 124128
rect 116176 124108 116178 124128
rect 116122 124072 116178 124108
rect 115938 122168 115994 122224
rect 116122 120128 116178 120184
rect 116122 118224 116178 118280
rect 116122 116320 116178 116376
rect 116122 114452 116124 114472
rect 116124 114452 116176 114472
rect 116176 114452 116178 114472
rect 116122 114416 116178 114452
rect 115938 112512 115994 112568
rect 116122 110608 116178 110664
rect 116122 108704 116178 108760
rect 116950 102856 117006 102912
rect 121458 153720 121514 153776
rect 121642 153720 121698 153776
rect 125966 152360 126022 152416
rect 126886 152360 126942 152416
rect 128634 152496 128690 152552
rect 131026 159296 131082 159352
rect 133786 159432 133842 159488
rect 131762 153992 131818 154048
rect 132406 153992 132462 154048
rect 133234 153992 133290 154048
rect 134338 153856 134394 153912
rect 133786 151816 133842 151872
rect 136270 151816 136326 151872
rect 138018 159568 138074 159624
rect 140134 156576 140190 156632
rect 142710 156712 142766 156768
rect 142158 154128 142214 154184
rect 142342 153992 142398 154048
rect 143078 154012 143134 154048
rect 143078 153992 143080 154012
rect 143080 153992 143132 154012
rect 143132 153992 143134 154012
rect 144918 157936 144974 157992
rect 143538 152360 143594 152416
rect 147402 159452 147458 159488
rect 147402 159432 147404 159452
rect 147404 159432 147456 159452
rect 147456 159432 147458 159452
rect 147678 159432 147734 159488
rect 147494 153992 147550 154048
rect 147862 153992 147918 154048
rect 149610 158072 149666 158128
rect 152186 158208 152242 158264
rect 161570 156848 161626 156904
rect 160650 154264 160706 154320
rect 162858 158344 162914 158400
rect 166354 155488 166410 155544
rect 168930 155216 168986 155272
rect 171230 155352 171286 155408
rect 174082 156984 174138 157040
rect 176842 155760 176898 155816
rect 178682 155624 178738 155680
rect 181074 154300 181076 154320
rect 181076 154300 181128 154320
rect 181128 154300 181130 154320
rect 181074 154264 181130 154300
rect 181442 154264 181498 154320
rect 183742 155896 183798 155952
rect 184386 154400 184442 154456
rect 186318 155080 186374 155136
rect 189170 155116 189172 155136
rect 189172 155116 189224 155136
rect 189224 155116 189226 155136
rect 189170 155080 189226 155116
rect 192114 153720 192170 153776
rect 195886 153584 195942 153640
rect 196070 153620 196072 153640
rect 196072 153620 196124 153640
rect 196124 153620 196126 153640
rect 196070 153584 196126 153620
rect 198738 158480 198794 158536
rect 204718 159296 204774 159352
rect 207018 157120 207074 157176
rect 212354 153720 212410 153776
rect 227442 152360 227498 152416
rect 274546 159432 274602 159488
rect 274822 159296 274878 159352
rect 280710 153720 280766 153776
rect 292578 152360 292634 152416
rect 313462 152360 313518 152416
rect 328458 159432 328514 159488
rect 357438 152360 357494 152416
rect 408314 152360 408370 152416
rect 430578 152360 430634 152416
rect 431866 152360 431922 152416
rect 439502 152924 439558 152960
rect 439502 152904 439504 152924
rect 439504 152904 439556 152924
rect 439556 152904 439558 152924
rect 442998 152924 443054 152960
rect 442998 152904 443000 152924
rect 443000 152904 443052 152924
rect 443052 152904 443054 152924
rect 448518 152360 448574 152416
rect 519726 163104 519782 163160
rect 519542 161608 519598 161664
rect 519634 160112 519690 160168
rect 519542 147872 519598 147928
rect 520186 158616 520242 158672
rect 520002 157120 520058 157176
rect 519818 151000 519874 151056
rect 519726 149232 519782 149288
rect 519726 148008 519782 148064
rect 519634 146512 519690 146568
rect 519542 143384 519598 143440
rect 519358 141888 519414 141944
rect 519910 149504 519966 149560
rect 519818 138352 519874 138408
rect 520094 153992 520150 154048
rect 520002 143792 520058 143848
rect 521198 155624 521254 155680
rect 521106 152496 521162 152552
rect 520922 146512 520978 146568
rect 520186 145152 520242 145208
rect 520094 141072 520150 141128
rect 520186 140392 520242 140448
rect 520002 138896 520058 138952
rect 519910 136992 519966 137048
rect 519910 135768 519966 135824
rect 519726 135632 519782 135688
rect 519818 134272 519874 134328
rect 519634 132776 519690 132832
rect 519542 131552 519598 131608
rect 519358 130192 519414 130248
rect 519542 129784 519598 129840
rect 117226 127880 117282 127936
rect 519450 126656 519506 126712
rect 519358 120536 519414 120592
rect 519726 131280 519782 131336
rect 519634 122032 519690 122088
rect 520094 137400 520150 137456
rect 520002 127472 520058 127528
rect 521014 144880 521070 144936
rect 520922 134408 520978 134464
rect 521198 142432 521254 142488
rect 521106 139712 521162 139768
rect 521014 132912 521070 132968
rect 520186 128832 520242 128888
rect 520186 128288 520242 128344
rect 520094 126112 520150 126168
rect 520094 125160 520150 125216
rect 519910 124752 519966 124808
rect 520002 123664 520058 123720
rect 519818 123392 519874 123448
rect 519818 122168 519874 122224
rect 519726 120672 519782 120728
rect 519542 119312 519598 119368
rect 519726 119176 519782 119232
rect 519542 117544 519598 117600
rect 519450 116592 519506 116648
rect 519358 111152 519414 111208
rect 519634 114552 519690 114608
rect 519542 108432 519598 108488
rect 519910 116048 519966 116104
rect 519818 112512 519874 112568
rect 519726 109792 519782 109848
rect 520186 117952 520242 118008
rect 520094 115232 520150 115288
rect 520002 113872 520058 113928
rect 520370 113056 520426 113112
rect 519910 107072 519966 107128
rect 519634 105712 519690 105768
rect 520278 105440 520334 105496
rect 117134 104760 117190 104816
rect 117042 100952 117098 101008
rect 519634 99320 519690 99376
rect 116858 99048 116914 99104
rect 116766 97144 116822 97200
rect 519266 96328 519322 96384
rect 116674 95240 116730 95296
rect 116582 93336 116638 93392
rect 116122 91296 116178 91352
rect 519726 97824 519782 97880
rect 519634 92112 519690 92168
rect 521566 111560 521622 111616
rect 521474 110064 521530 110120
rect 521106 108432 521162 108488
rect 520370 104352 520426 104408
rect 520922 103944 520978 104000
rect 520278 97552 520334 97608
rect 521014 102448 521070 102504
rect 520922 96192 520978 96248
rect 521382 106936 521438 106992
rect 521198 100952 521254 101008
rect 521106 100272 521162 100328
rect 521014 94968 521070 95024
rect 520002 94832 520058 94888
rect 519726 90752 519782 90808
rect 116122 89392 116178 89448
rect 519266 89392 519322 89448
rect 521566 102992 521622 103048
rect 521474 101632 521530 101688
rect 521382 98912 521438 98968
rect 521198 93472 521254 93528
rect 520186 93336 520242 93392
rect 520002 88032 520058 88088
rect 116030 87488 116086 87544
rect 521290 91840 521346 91896
rect 520922 90208 520978 90264
rect 520186 86672 520242 86728
rect 520278 85720 520334 85776
rect 115202 85584 115258 85640
rect 116582 83680 116638 83736
rect 520002 82728 520058 82784
rect 116214 81776 116270 81832
rect 115938 79872 115994 79928
rect 519634 79600 519690 79656
rect 116122 77968 116178 78024
rect 116674 74024 116730 74080
rect 116582 72120 116638 72176
rect 113362 64504 113418 64560
rect 110326 57976 110382 58032
rect 110326 56752 110382 56808
rect 110326 53896 110382 53952
rect 110326 52536 110382 52592
rect 110326 51040 110382 51096
rect 110326 48320 110382 48376
rect 110326 47096 110382 47152
rect 110326 42880 110382 42936
rect 110326 42336 110382 42392
rect 110418 34992 110474 35048
rect 110326 34720 110382 34776
rect 110326 34584 110382 34640
rect 110694 42336 110750 42392
rect 110602 41384 110658 41440
rect 110602 34584 110658 34640
rect 110694 29824 110750 29880
rect 111062 44240 111118 44296
rect 110878 42880 110934 42936
rect 110326 29416 110382 29472
rect 110326 29280 110382 29336
rect 110326 29144 110382 29200
rect 33046 2624 33102 2680
rect 42062 2624 42118 2680
rect 42706 2624 42762 2680
rect 44730 2624 44786 2680
rect 58990 2624 59046 2680
rect 59174 2624 59230 2680
rect 62762 2624 62818 2680
rect 63038 2624 63094 2680
rect 64602 2624 64658 2680
rect 66994 2624 67050 2680
rect 76562 2624 76618 2680
rect 89166 2624 89222 2680
rect 89718 2624 89774 2680
rect 89902 2624 89958 2680
rect 90362 2624 90418 2680
rect 92478 2624 92534 2680
rect 92754 2624 92810 2680
rect 95146 2624 95202 2680
rect 95330 2624 95386 2680
rect 96434 2624 96490 2680
rect 99930 2624 99986 2680
rect 100850 2624 100906 2680
rect 101770 2624 101826 2680
rect 101954 2624 102010 2680
rect 102782 2624 102838 2680
rect 29550 2488 29606 2544
rect 26054 2352 26110 2408
rect 22926 2216 22982 2272
rect 5998 1808 6054 1864
rect 19614 2080 19670 2136
rect 16210 1944 16266 2000
rect 12622 1672 12678 1728
rect 9310 1536 9366 1592
rect 55954 1400 56010 1456
rect 89166 1128 89222 1184
rect 89902 1264 89958 1320
rect 95146 1128 95202 1184
rect 96434 1264 96490 1320
rect 98274 1264 98330 1320
rect 101954 1264 102010 1320
rect 110326 20168 110382 20224
rect 110326 12416 110382 12472
rect 110326 12144 110382 12200
rect 110510 29552 110566 29608
rect 110970 34992 111026 35048
rect 110602 20032 110658 20088
rect 110602 12144 110658 12200
rect 110510 9696 110566 9752
rect 110326 9016 110382 9072
rect 110326 8744 110382 8800
rect 110326 8472 110382 8528
rect 110326 8336 110382 8392
rect 110418 7792 110474 7848
rect 109866 3168 109922 3224
rect 109866 2896 109922 2952
rect 110602 9016 110658 9072
rect 110786 29416 110842 29472
rect 111246 34720 111302 34776
rect 111154 34584 111210 34640
rect 111062 29552 111118 29608
rect 111154 29280 111210 29336
rect 111338 29824 111394 29880
rect 111246 29144 111302 29200
rect 110786 20168 110842 20224
rect 110786 20032 110842 20088
rect 110050 3848 110106 3904
rect 110970 12416 111026 12472
rect 110878 9696 110934 9752
rect 110970 8744 111026 8800
rect 111062 8472 111118 8528
rect 111338 8336 111394 8392
rect 110970 7792 111026 7848
rect 110878 5616 110934 5672
rect 110326 5492 110382 5548
rect 110694 4120 110750 4176
rect 110326 2896 110382 2952
rect 110326 1808 110382 1864
rect 110970 3576 111026 3632
rect 110694 2896 110750 2952
rect 111706 2796 111708 2816
rect 111708 2796 111760 2816
rect 111760 2796 111762 2816
rect 111706 2760 111762 2796
rect 116306 70216 116362 70272
rect 116122 68312 116178 68368
rect 116582 66408 116638 66464
rect 519266 73616 519322 73672
rect 519726 78104 519782 78160
rect 519634 73208 519690 73264
rect 520186 81096 520242 81152
rect 520094 76608 520150 76664
rect 520002 75928 520058 75984
rect 520002 75112 520058 75168
rect 519726 72392 519782 72448
rect 519450 71984 519506 72040
rect 519266 67768 519322 67824
rect 519266 67496 519322 67552
rect 116214 64504 116270 64560
rect 116122 62600 116178 62656
rect 521014 87216 521070 87272
rect 520922 82592 520978 82648
rect 521198 84224 521254 84280
rect 521014 79872 521070 79928
rect 520278 78512 520334 78568
rect 521382 88712 521438 88768
rect 521290 83952 521346 84008
rect 521382 81232 521438 81288
rect 521198 77152 521254 77208
rect 520186 74568 520242 74624
rect 520094 70488 520150 70544
rect 520186 70352 520242 70408
rect 520002 69128 520058 69184
rect 519634 68992 519690 69048
rect 519450 66408 519506 66464
rect 519818 66000 519874 66056
rect 519634 63688 519690 63744
rect 519266 60968 519322 61024
rect 116582 60560 116638 60616
rect 114190 53080 114246 53136
rect 116122 43288 116178 43344
rect 114098 41792 114154 41848
rect 114006 30368 114062 30424
rect 116398 26016 116454 26072
rect 116306 20304 116362 20360
rect 113914 18944 113970 19000
rect 116214 18400 116270 18456
rect 116030 16360 116086 16416
rect 115938 12552 115994 12608
rect 113822 7656 113878 7712
rect 116122 14456 116178 14512
rect 116030 2352 116086 2408
rect 116490 22208 116546 22264
rect 116306 3304 116362 3360
rect 116306 3032 116362 3088
rect 116214 2488 116270 2544
rect 116122 2216 116178 2272
rect 115938 2080 115994 2136
rect 520186 65048 520242 65104
rect 521106 64504 521162 64560
rect 520738 62872 520794 62928
rect 520278 61376 520334 61432
rect 519818 59608 519874 59664
rect 520186 56888 520242 56944
rect 521106 62328 521162 62384
rect 521014 59880 521070 59936
rect 520738 58248 520794 58304
rect 520370 56888 520426 56944
rect 520278 55392 520334 55448
rect 519266 53760 519322 53816
rect 520094 52264 520150 52320
rect 520002 50768 520058 50824
rect 519266 50088 519322 50144
rect 519450 47776 519506 47832
rect 521106 58384 521162 58440
rect 521014 55528 521070 55584
rect 521106 54168 521162 54224
rect 520370 52808 520426 52864
rect 520278 51448 520334 51504
rect 520186 49272 520242 49328
rect 520094 48728 520150 48784
rect 520002 47368 520058 47424
rect 519910 46280 519966 46336
rect 519450 44648 519506 44704
rect 519818 44648 519874 44704
rect 520186 46008 520242 46064
rect 519910 43288 519966 43344
rect 520186 43152 520242 43208
rect 519818 41928 519874 41984
rect 520094 41656 520150 41712
rect 116766 39480 116822 39536
rect 116674 37576 116730 37632
rect 520186 40568 520242 40624
rect 520186 40160 520242 40216
rect 520094 39208 520150 39264
rect 519818 38664 519874 38720
rect 520186 37848 520242 37904
rect 521566 37168 521622 37224
rect 519818 36488 519874 36544
rect 521566 35944 521622 36000
rect 521106 35536 521162 35592
rect 521106 34448 521162 34504
rect 520922 34040 520978 34096
rect 116950 33768 117006 33824
rect 116858 31728 116914 31784
rect 116766 3168 116822 3224
rect 520922 33088 520978 33144
rect 520922 32544 520978 32600
rect 520922 31592 520978 31648
rect 520922 31048 520978 31104
rect 520922 30232 520978 30288
rect 117042 29824 117098 29880
rect 116950 3712 117006 3768
rect 521106 29552 521162 29608
rect 521106 28328 521162 28384
rect 117134 27920 117190 27976
rect 117226 24112 117282 24168
rect 117134 3440 117190 3496
rect 521106 21936 521162 21992
rect 521106 20848 521162 20904
rect 520738 20440 520794 20496
rect 520738 19488 520794 19544
rect 520922 18944 520978 19000
rect 520922 18128 520978 18184
rect 521106 9288 521162 9344
rect 521106 8200 521162 8256
rect 520370 7928 520426 7984
rect 520370 6704 520426 6760
rect 521106 6568 521162 6624
rect 520922 5208 520978 5264
rect 521106 5208 521162 5264
rect 521014 3848 521070 3904
rect 520922 3712 520978 3768
rect 163778 1536 163834 1592
rect 229282 1672 229338 1728
rect 293590 1672 293646 1728
rect 243634 1536 243690 1592
rect 294786 1420 294842 1456
rect 294786 1400 294788 1420
rect 294788 1400 294840 1420
rect 294840 1400 294842 1420
rect 360290 1400 360346 1456
rect 393594 1400 393650 1456
rect 521106 2624 521162 2680
rect 521014 2216 521070 2272
rect 521106 720 521162 776
<< metal3 >>
rect 519721 163162 519787 163165
rect 523200 163162 524400 163192
rect 519721 163160 524400 163162
rect 519721 163104 519726 163160
rect 519782 163104 524400 163160
rect 519721 163102 524400 163104
rect 519721 163099 519787 163102
rect 523200 163072 524400 163102
rect 519537 161666 519603 161669
rect 523200 161666 524400 161696
rect 519537 161664 524400 161666
rect 519537 161608 519542 161664
rect 519598 161608 524400 161664
rect 519537 161606 524400 161608
rect 519537 161603 519603 161606
rect 523200 161576 524400 161606
rect 519629 160170 519695 160173
rect 523200 160170 524400 160200
rect 519629 160168 524400 160170
rect 519629 160112 519634 160168
rect 519690 160112 524400 160168
rect 519629 160110 524400 160112
rect 519629 160107 519695 160110
rect 523200 160080 524400 160110
rect 29821 159626 29887 159629
rect 138013 159626 138079 159629
rect 29821 159624 138079 159626
rect 29821 159568 29826 159624
rect 29882 159568 138018 159624
rect 138074 159568 138079 159624
rect 29821 159566 138079 159568
rect 29821 159563 29887 159566
rect 138013 159563 138079 159566
rect 23013 159490 23079 159493
rect 133781 159490 133847 159493
rect 23013 159488 133847 159490
rect 23013 159432 23018 159488
rect 23074 159432 133786 159488
rect 133842 159432 133847 159488
rect 23013 159430 133847 159432
rect 23013 159427 23079 159430
rect 133781 159427 133847 159430
rect 147397 159490 147463 159493
rect 147673 159490 147739 159493
rect 147397 159488 147739 159490
rect 147397 159432 147402 159488
rect 147458 159432 147678 159488
rect 147734 159432 147739 159488
rect 147397 159430 147739 159432
rect 147397 159427 147463 159430
rect 147673 159427 147739 159430
rect 274541 159490 274607 159493
rect 328453 159490 328519 159493
rect 274541 159488 328519 159490
rect 274541 159432 274546 159488
rect 274602 159432 328458 159488
rect 328514 159432 328519 159488
rect 274541 159430 328519 159432
rect 274541 159427 274607 159430
rect 328453 159427 328519 159430
rect 16297 159354 16363 159357
rect 131021 159354 131087 159357
rect 16297 159352 131087 159354
rect 16297 159296 16302 159352
rect 16358 159296 131026 159352
rect 131082 159296 131087 159352
rect 16297 159294 131087 159296
rect 16297 159291 16363 159294
rect 131021 159291 131087 159294
rect 204713 159354 204779 159357
rect 274817 159354 274883 159357
rect 204713 159352 274883 159354
rect 204713 159296 204718 159352
rect 204774 159296 274822 159352
rect 274878 159296 274883 159352
rect 204713 159294 274883 159296
rect 204713 159291 204779 159294
rect 274817 159291 274883 159294
rect 520181 158674 520247 158677
rect 523200 158674 524400 158704
rect 520181 158672 524400 158674
rect 520181 158616 520186 158672
rect 520242 158616 524400 158672
rect 520181 158614 524400 158616
rect 520181 158611 520247 158614
rect 523200 158584 524400 158614
rect 104617 158538 104683 158541
rect 198733 158538 198799 158541
rect 104617 158536 198799 158538
rect 104617 158480 104622 158536
rect 104678 158480 198738 158536
rect 198794 158480 198799 158536
rect 104617 158478 198799 158480
rect 104617 158475 104683 158478
rect 198733 158475 198799 158478
rect 57513 158402 57579 158405
rect 162853 158402 162919 158405
rect 57513 158400 162919 158402
rect 57513 158344 57518 158400
rect 57574 158344 162858 158400
rect 162914 158344 162919 158400
rect 57513 158342 162919 158344
rect 57513 158339 57579 158342
rect 162853 158339 162919 158342
rect 44081 158266 44147 158269
rect 152181 158266 152247 158269
rect 44081 158264 152247 158266
rect 44081 158208 44086 158264
rect 44142 158208 152186 158264
rect 152242 158208 152247 158264
rect 44081 158206 152247 158208
rect 44081 158203 44147 158206
rect 152181 158203 152247 158206
rect 40677 158130 40743 158133
rect 149605 158130 149671 158133
rect 40677 158128 149671 158130
rect 40677 158072 40682 158128
rect 40738 158072 149610 158128
rect 149666 158072 149671 158128
rect 40677 158070 149671 158072
rect 40677 158067 40743 158070
rect 149605 158067 149671 158070
rect 33961 157994 34027 157997
rect 144913 157994 144979 157997
rect 33961 157992 144979 157994
rect 33961 157936 33966 157992
rect 34022 157936 144918 157992
rect 144974 157936 144979 157992
rect 33961 157934 144979 157936
rect 33961 157931 34027 157934
rect 144913 157931 144979 157934
rect 115565 157178 115631 157181
rect 207013 157178 207079 157181
rect 115565 157176 207079 157178
rect 115565 157120 115570 157176
rect 115626 157120 207018 157176
rect 207074 157120 207079 157176
rect 115565 157118 207079 157120
rect 115565 157115 115631 157118
rect 207013 157115 207079 157118
rect 519997 157178 520063 157181
rect 523200 157178 524400 157208
rect 519997 157176 524400 157178
rect 519997 157120 520002 157176
rect 520058 157120 524400 157176
rect 519997 157118 524400 157120
rect 519997 157115 520063 157118
rect 523200 157088 524400 157118
rect 72693 157042 72759 157045
rect 174077 157042 174143 157045
rect 72693 157040 174143 157042
rect 72693 156984 72698 157040
rect 72754 156984 174082 157040
rect 174138 156984 174143 157040
rect 72693 156982 174143 156984
rect 72693 156979 72759 156982
rect 174077 156979 174143 156982
rect 55857 156906 55923 156909
rect 161565 156906 161631 156909
rect 55857 156904 161631 156906
rect 55857 156848 55862 156904
rect 55918 156848 161570 156904
rect 161626 156848 161631 156904
rect 55857 156846 161631 156848
rect 55857 156843 55923 156846
rect 161565 156843 161631 156846
rect 31477 156770 31543 156773
rect 142705 156770 142771 156773
rect 31477 156768 142771 156770
rect 31477 156712 31482 156768
rect 31538 156712 142710 156768
rect 142766 156712 142771 156768
rect 31477 156710 142771 156712
rect 31477 156707 31543 156710
rect 142705 156707 142771 156710
rect 28073 156634 28139 156637
rect 140129 156634 140195 156637
rect 28073 156632 140195 156634
rect 28073 156576 28078 156632
rect 28134 156576 140134 156632
rect 140190 156576 140195 156632
rect 28073 156574 140195 156576
rect 28073 156571 28139 156574
rect 140129 156571 140195 156574
rect 85297 155954 85363 155957
rect 183737 155954 183803 155957
rect 85297 155952 183803 155954
rect 85297 155896 85302 155952
rect 85358 155896 183742 155952
rect 183798 155896 183803 155952
rect 85297 155894 183803 155896
rect 85297 155891 85363 155894
rect 183737 155891 183803 155894
rect 76005 155818 76071 155821
rect 176837 155818 176903 155821
rect 76005 155816 176903 155818
rect 76005 155760 76010 155816
rect 76066 155760 176842 155816
rect 176898 155760 176903 155816
rect 76005 155758 176903 155760
rect 76005 155755 76071 155758
rect 176837 155755 176903 155758
rect 78581 155682 78647 155685
rect 178677 155682 178743 155685
rect 78581 155680 178743 155682
rect 78581 155624 78586 155680
rect 78642 155624 178682 155680
rect 178738 155624 178743 155680
rect 78581 155622 178743 155624
rect 78581 155619 78647 155622
rect 178677 155619 178743 155622
rect 521193 155682 521259 155685
rect 523200 155682 524400 155712
rect 521193 155680 524400 155682
rect 521193 155624 521198 155680
rect 521254 155624 524400 155680
rect 521193 155622 524400 155624
rect 521193 155619 521259 155622
rect 523200 155592 524400 155622
rect 62573 155546 62639 155549
rect 166349 155546 166415 155549
rect 62573 155544 166415 155546
rect 62573 155488 62578 155544
rect 62634 155488 166354 155544
rect 166410 155488 166415 155544
rect 62573 155486 166415 155488
rect 62573 155483 62639 155486
rect 166349 155483 166415 155486
rect 68461 155410 68527 155413
rect 171225 155410 171291 155413
rect 68461 155408 171291 155410
rect 68461 155352 68466 155408
rect 68522 155352 171230 155408
rect 171286 155352 171291 155408
rect 68461 155350 171291 155352
rect 68461 155347 68527 155350
rect 171225 155347 171291 155350
rect 65977 155274 66043 155277
rect 168925 155274 168991 155277
rect 65977 155272 168991 155274
rect 65977 155216 65982 155272
rect 66038 155216 168930 155272
rect 168986 155216 168991 155272
rect 65977 155214 168991 155216
rect 65977 155211 66043 155214
rect 168925 155211 168991 155214
rect 186313 155138 186379 155141
rect 189165 155138 189231 155141
rect 186313 155136 189231 155138
rect 186313 155080 186318 155136
rect 186374 155080 189170 155136
rect 189226 155080 189231 155136
rect 186313 155078 189231 155080
rect 186313 155075 186379 155078
rect 189165 155075 189231 155078
rect 86125 154458 86191 154461
rect 184381 154458 184447 154461
rect 86125 154456 184447 154458
rect 86125 154400 86130 154456
rect 86186 154400 184386 154456
rect 184442 154400 184447 154456
rect 86125 154398 184447 154400
rect 86125 154395 86191 154398
rect 184381 154395 184447 154398
rect 55029 154322 55095 154325
rect 160645 154322 160711 154325
rect 55029 154320 160711 154322
rect 55029 154264 55034 154320
rect 55090 154264 160650 154320
rect 160706 154264 160711 154320
rect 55029 154262 160711 154264
rect 55029 154259 55095 154262
rect 160645 154259 160711 154262
rect 181069 154322 181135 154325
rect 181437 154322 181503 154325
rect 181069 154320 181503 154322
rect 181069 154264 181074 154320
rect 181130 154264 181442 154320
rect 181498 154264 181503 154320
rect 181069 154262 181503 154264
rect 181069 154259 181135 154262
rect 181437 154259 181503 154262
rect 30649 154186 30715 154189
rect 142153 154186 142219 154189
rect 30649 154184 142219 154186
rect 30649 154128 30654 154184
rect 30710 154128 142158 154184
rect 142214 154128 142219 154184
rect 30649 154126 142219 154128
rect 30649 154123 30715 154126
rect 142153 154123 142219 154126
rect 17125 154050 17191 154053
rect 131757 154050 131823 154053
rect 17125 154048 131823 154050
rect 17125 153992 17130 154048
rect 17186 153992 131762 154048
rect 131818 153992 131823 154048
rect 17125 153990 131823 153992
rect 17125 153987 17191 153990
rect 131757 153987 131823 153990
rect 132401 154050 132467 154053
rect 133229 154050 133295 154053
rect 132401 154048 133295 154050
rect 132401 153992 132406 154048
rect 132462 153992 133234 154048
rect 133290 153992 133295 154048
rect 132401 153990 133295 153992
rect 132401 153987 132467 153990
rect 133229 153987 133295 153990
rect 142337 154050 142403 154053
rect 143073 154050 143139 154053
rect 142337 154048 143139 154050
rect 142337 153992 142342 154048
rect 142398 153992 143078 154048
rect 143134 153992 143139 154048
rect 142337 153990 143139 153992
rect 142337 153987 142403 153990
rect 143073 153987 143139 153990
rect 147489 154050 147555 154053
rect 147857 154050 147923 154053
rect 147489 154048 147923 154050
rect 147489 153992 147494 154048
rect 147550 153992 147862 154048
rect 147918 153992 147923 154048
rect 147489 153990 147923 153992
rect 147489 153987 147555 153990
rect 147857 153987 147923 153990
rect 520089 154050 520155 154053
rect 523200 154050 524400 154080
rect 520089 154048 524400 154050
rect 520089 153992 520094 154048
rect 520150 153992 524400 154048
rect 520089 153990 524400 153992
rect 520089 153987 520155 153990
rect 523200 153960 524400 153990
rect 20529 153914 20595 153917
rect 134333 153914 134399 153917
rect 20529 153912 134399 153914
rect 20529 153856 20534 153912
rect 20590 153856 134338 153912
rect 134394 153856 134399 153912
rect 20529 153854 134399 153856
rect 20529 153851 20595 153854
rect 134333 153851 134399 153854
rect 3969 153778 4035 153781
rect 121453 153778 121519 153781
rect 3969 153776 121519 153778
rect 3969 153720 3974 153776
rect 4030 153720 121458 153776
rect 121514 153720 121519 153776
rect 3969 153718 121519 153720
rect 3969 153715 4035 153718
rect 121453 153715 121519 153718
rect 121637 153778 121703 153781
rect 192109 153778 192175 153781
rect 121637 153776 192175 153778
rect 121637 153720 121642 153776
rect 121698 153720 192114 153776
rect 192170 153720 192175 153776
rect 121637 153718 192175 153720
rect 121637 153715 121703 153718
rect 192109 153715 192175 153718
rect 212349 153778 212415 153781
rect 280705 153778 280771 153781
rect 212349 153776 280771 153778
rect 212349 153720 212354 153776
rect 212410 153720 280710 153776
rect 280766 153720 280771 153776
rect 212349 153718 280771 153720
rect 212349 153715 212415 153718
rect 280705 153715 280771 153718
rect 195881 153642 195947 153645
rect 196065 153642 196131 153645
rect 195881 153640 196131 153642
rect 195881 153584 195886 153640
rect 195942 153584 196070 153640
rect 196126 153584 196131 153640
rect 195881 153582 196131 153584
rect 195881 153579 195947 153582
rect 196065 153579 196131 153582
rect 439497 152962 439563 152965
rect 442993 152962 443059 152965
rect 439497 152960 443059 152962
rect 439497 152904 439502 152960
rect 439558 152904 442998 152960
rect 443054 152904 443059 152960
rect 439497 152902 443059 152904
rect 439497 152899 439563 152902
rect 442993 152899 443059 152902
rect 12985 152554 13051 152557
rect 128629 152554 128695 152557
rect 12985 152552 128695 152554
rect 12985 152496 12990 152552
rect 13046 152496 128634 152552
rect 128690 152496 128695 152552
rect 12985 152494 128695 152496
rect 12985 152491 13051 152494
rect 128629 152491 128695 152494
rect 521101 152554 521167 152557
rect 523200 152554 524400 152584
rect 521101 152552 524400 152554
rect 521101 152496 521106 152552
rect 521162 152496 524400 152552
rect 521101 152494 524400 152496
rect 521101 152491 521167 152494
rect 523200 152464 524400 152494
rect 9581 152418 9647 152421
rect 125961 152418 126027 152421
rect 9581 152416 126027 152418
rect 9581 152360 9586 152416
rect 9642 152360 125966 152416
rect 126022 152360 126027 152416
rect 9581 152358 126027 152360
rect 9581 152355 9647 152358
rect 125961 152355 126027 152358
rect 126881 152418 126947 152421
rect 143533 152418 143599 152421
rect 126881 152416 143599 152418
rect 126881 152360 126886 152416
rect 126942 152360 143538 152416
rect 143594 152360 143599 152416
rect 126881 152358 143599 152360
rect 126881 152355 126947 152358
rect 143533 152355 143599 152358
rect 227437 152418 227503 152421
rect 292573 152418 292639 152421
rect 227437 152416 292639 152418
rect 227437 152360 227442 152416
rect 227498 152360 292578 152416
rect 292634 152360 292639 152416
rect 227437 152358 292639 152360
rect 227437 152355 227503 152358
rect 292573 152355 292639 152358
rect 313457 152418 313523 152421
rect 357433 152418 357499 152421
rect 313457 152416 357499 152418
rect 313457 152360 313462 152416
rect 313518 152360 357438 152416
rect 357494 152360 357499 152416
rect 313457 152358 357499 152360
rect 313457 152355 313523 152358
rect 357433 152355 357499 152358
rect 408309 152418 408375 152421
rect 430573 152418 430639 152421
rect 408309 152416 430639 152418
rect 408309 152360 408314 152416
rect 408370 152360 430578 152416
rect 430634 152360 430639 152416
rect 408309 152358 430639 152360
rect 408309 152355 408375 152358
rect 430573 152355 430639 152358
rect 431861 152418 431927 152421
rect 448513 152418 448579 152421
rect 431861 152416 448579 152418
rect 431861 152360 431866 152416
rect 431922 152360 448518 152416
rect 448574 152360 448579 152416
rect 431861 152358 448579 152360
rect 431861 152355 431927 152358
rect 448513 152355 448579 152358
rect 133781 151874 133847 151877
rect 136265 151874 136331 151877
rect 133781 151872 136331 151874
rect 133781 151816 133786 151872
rect 133842 151816 136270 151872
rect 136326 151816 136331 151872
rect 133781 151814 136331 151816
rect 133781 151811 133847 151814
rect 136265 151811 136331 151814
rect 519813 151058 519879 151061
rect 523200 151058 524400 151088
rect 519813 151056 524400 151058
rect 519813 151000 519818 151056
rect 519874 151000 524400 151056
rect 519813 150998 524400 151000
rect 519813 150995 519879 150998
rect 523200 150968 524400 150998
rect 6085 150650 6151 150653
rect 111333 150650 111399 150653
rect 6085 150648 111399 150650
rect 6085 150592 6090 150648
rect 6146 150592 111338 150648
rect 111394 150592 111399 150648
rect 6085 150590 111399 150592
rect 6085 150587 6151 150590
rect 111333 150587 111399 150590
rect 2681 150514 2747 150517
rect 111057 150514 111123 150517
rect 2681 150512 111123 150514
rect 2681 150456 2686 150512
rect 2742 150456 111062 150512
rect 111118 150456 111123 150512
rect 2681 150454 111123 150456
rect 2681 150451 2747 150454
rect 111057 150451 111123 150454
rect 82813 149698 82879 149701
rect 116577 149698 116643 149701
rect 82813 149696 116643 149698
rect 82813 149640 82818 149696
rect 82874 149640 116582 149696
rect 116638 149640 116643 149696
rect 82813 149638 116643 149640
rect 82813 149635 82879 149638
rect 116577 149635 116643 149638
rect 519905 149562 519971 149565
rect 523200 149562 524400 149592
rect 519905 149560 524400 149562
rect 519905 149504 519910 149560
rect 519966 149504 524400 149560
rect 519905 149502 524400 149504
rect 519905 149499 519971 149502
rect 523200 149472 524400 149502
rect 519721 149290 519787 149293
rect 518788 149288 519787 149290
rect 518788 149232 519726 149288
rect 519782 149232 519787 149288
rect 518788 149230 519787 149232
rect 519721 149227 519787 149230
rect 109585 148066 109651 148069
rect 119110 148066 119170 148988
rect 109585 148064 119170 148066
rect 109585 148008 109590 148064
rect 109646 148008 119170 148064
rect 109585 148006 119170 148008
rect 519721 148066 519787 148069
rect 523200 148066 524400 148096
rect 519721 148064 524400 148066
rect 519721 148008 519726 148064
rect 519782 148008 524400 148064
rect 519721 148006 524400 148008
rect 109585 148003 109651 148006
rect 519721 148003 519787 148006
rect 523200 147976 524400 148006
rect 519537 147930 519603 147933
rect 518788 147928 519603 147930
rect 518788 147872 519542 147928
rect 519598 147872 519603 147928
rect 518788 147870 519603 147872
rect 519537 147867 519603 147870
rect 110965 147386 111031 147389
rect 111701 147386 111767 147389
rect 110965 147384 111767 147386
rect 110965 147328 110970 147384
rect 111026 147328 111706 147384
rect 111762 147328 111767 147384
rect 110965 147326 111767 147328
rect 110965 147323 111031 147326
rect 111701 147323 111767 147326
rect 110321 146434 110387 146437
rect 119110 146434 119170 147084
rect 519629 146570 519695 146573
rect 518788 146568 519695 146570
rect 518788 146512 519634 146568
rect 519690 146512 519695 146568
rect 518788 146510 519695 146512
rect 519629 146507 519695 146510
rect 520917 146570 520983 146573
rect 523200 146570 524400 146600
rect 520917 146568 524400 146570
rect 520917 146512 520922 146568
rect 520978 146512 524400 146568
rect 520917 146510 524400 146512
rect 520917 146507 520983 146510
rect 523200 146480 524400 146510
rect 110321 146432 119170 146434
rect 110321 146376 110326 146432
rect 110382 146376 119170 146432
rect 110321 146374 119170 146376
rect 110321 146371 110387 146374
rect 116117 145210 116183 145213
rect 520181 145210 520247 145213
rect 116117 145208 119140 145210
rect 116117 145152 116122 145208
rect 116178 145152 119140 145208
rect 116117 145150 119140 145152
rect 518788 145208 520247 145210
rect 518788 145152 520186 145208
rect 520242 145152 520247 145208
rect 518788 145150 520247 145152
rect 116117 145147 116183 145150
rect 520181 145147 520247 145150
rect 521009 144938 521075 144941
rect 523200 144938 524400 144968
rect 521009 144936 524400 144938
rect 521009 144880 521014 144936
rect 521070 144880 524400 144936
rect 521009 144878 524400 144880
rect 521009 144875 521075 144878
rect 523200 144848 524400 144878
rect 113817 144258 113883 144261
rect 110860 144256 113883 144258
rect 110860 144200 113822 144256
rect 113878 144200 113883 144256
rect 110860 144198 113883 144200
rect 113817 144195 113883 144198
rect 519997 143850 520063 143853
rect 518788 143848 520063 143850
rect 518788 143792 520002 143848
rect 520058 143792 520063 143848
rect 518788 143790 520063 143792
rect 519997 143787 520063 143790
rect 519537 143442 519603 143445
rect 523200 143442 524400 143472
rect 519537 143440 524400 143442
rect 519537 143384 519542 143440
rect 519598 143384 524400 143440
rect 519537 143382 524400 143384
rect 519537 143379 519603 143382
rect 523200 143352 524400 143382
rect 116025 143306 116091 143309
rect 116025 143304 119140 143306
rect 116025 143248 116030 143304
rect 116086 143248 119140 143304
rect 116025 143246 119140 143248
rect 116025 143243 116091 143246
rect 521193 142490 521259 142493
rect 518788 142488 521259 142490
rect 518788 142432 521198 142488
rect 521254 142432 521259 142488
rect 518788 142430 521259 142432
rect 521193 142427 521259 142430
rect 519353 141946 519419 141949
rect 523200 141946 524400 141976
rect 519353 141944 524400 141946
rect 519353 141888 519358 141944
rect 519414 141888 524400 141944
rect 519353 141886 524400 141888
rect 519353 141883 519419 141886
rect 523200 141856 524400 141886
rect 115289 141402 115355 141405
rect 115289 141400 119140 141402
rect 115289 141344 115294 141400
rect 115350 141344 119140 141400
rect 115289 141342 119140 141344
rect 115289 141339 115355 141342
rect 520089 141130 520155 141133
rect 518788 141128 520155 141130
rect 518788 141072 520094 141128
rect 520150 141072 520155 141128
rect 518788 141070 520155 141072
rect 520089 141067 520155 141070
rect 520181 140450 520247 140453
rect 523200 140450 524400 140480
rect 520181 140448 524400 140450
rect 520181 140392 520186 140448
rect 520242 140392 524400 140448
rect 520181 140390 524400 140392
rect 520181 140387 520247 140390
rect 523200 140360 524400 140390
rect 521101 139770 521167 139773
rect 518788 139768 521167 139770
rect 518788 139712 521106 139768
rect 521162 139712 521167 139768
rect 518788 139710 521167 139712
rect 521101 139707 521167 139710
rect 116117 139498 116183 139501
rect 116117 139496 119140 139498
rect 116117 139440 116122 139496
rect 116178 139440 119140 139496
rect 116117 139438 119140 139440
rect 116117 139435 116183 139438
rect 519997 138954 520063 138957
rect 523200 138954 524400 138984
rect 519997 138952 524400 138954
rect 519997 138896 520002 138952
rect 520058 138896 524400 138952
rect 519997 138894 524400 138896
rect 519997 138891 520063 138894
rect 523200 138864 524400 138894
rect 519813 138410 519879 138413
rect 518788 138408 519879 138410
rect 518788 138352 519818 138408
rect 519874 138352 519879 138408
rect 518788 138350 519879 138352
rect 519813 138347 519879 138350
rect 116117 137594 116183 137597
rect 116117 137592 119140 137594
rect 116117 137536 116122 137592
rect 116178 137536 119140 137592
rect 116117 137534 119140 137536
rect 116117 137531 116183 137534
rect 520089 137458 520155 137461
rect 523200 137458 524400 137488
rect 520089 137456 524400 137458
rect 520089 137400 520094 137456
rect 520150 137400 524400 137456
rect 520089 137398 524400 137400
rect 520089 137395 520155 137398
rect 523200 137368 524400 137398
rect 519905 137050 519971 137053
rect 518788 137048 519971 137050
rect 518788 136992 519910 137048
rect 519966 136992 519971 137048
rect 518788 136990 519971 136992
rect 519905 136987 519971 136990
rect 519905 135826 519971 135829
rect 523200 135826 524400 135856
rect 519905 135824 524400 135826
rect 519905 135768 519910 135824
rect 519966 135768 524400 135824
rect 519905 135766 524400 135768
rect 519905 135763 519971 135766
rect 523200 135736 524400 135766
rect 519721 135690 519787 135693
rect 518788 135688 519787 135690
rect 518788 135632 519726 135688
rect 519782 135632 519787 135688
rect 518788 135630 519787 135632
rect 519721 135627 519787 135630
rect 115197 135554 115263 135557
rect 115197 135552 119140 135554
rect 115197 135496 115202 135552
rect 115258 135496 119140 135552
rect 115197 135494 119140 135496
rect 115197 135491 115263 135494
rect 520917 134466 520983 134469
rect 518758 134464 520983 134466
rect 518758 134408 520922 134464
rect 520978 134408 520983 134464
rect 518758 134406 520983 134408
rect 518758 134300 518818 134406
rect 520917 134403 520983 134406
rect 519813 134330 519879 134333
rect 523200 134330 524400 134360
rect 519813 134328 524400 134330
rect 519813 134272 519818 134328
rect 519874 134272 524400 134328
rect 519813 134270 524400 134272
rect 519813 134267 519879 134270
rect 523200 134240 524400 134270
rect 116025 133650 116091 133653
rect 116025 133648 119140 133650
rect 116025 133592 116030 133648
rect 116086 133592 119140 133648
rect 116025 133590 119140 133592
rect 116025 133587 116091 133590
rect 521009 132970 521075 132973
rect 518788 132968 521075 132970
rect 518788 132912 521014 132968
rect 521070 132912 521075 132968
rect 518788 132910 521075 132912
rect 521009 132907 521075 132910
rect 114185 132834 114251 132837
rect 110860 132832 114251 132834
rect 110860 132776 114190 132832
rect 114246 132776 114251 132832
rect 110860 132774 114251 132776
rect 114185 132771 114251 132774
rect 519629 132834 519695 132837
rect 523200 132834 524400 132864
rect 519629 132832 524400 132834
rect 519629 132776 519634 132832
rect 519690 132776 524400 132832
rect 519629 132774 524400 132776
rect 519629 132771 519695 132774
rect 523200 132744 524400 132774
rect 116117 131746 116183 131749
rect 116117 131744 119140 131746
rect 116117 131688 116122 131744
rect 116178 131688 119140 131744
rect 116117 131686 119140 131688
rect 116117 131683 116183 131686
rect 519537 131610 519603 131613
rect 518788 131608 519603 131610
rect 518788 131552 519542 131608
rect 519598 131552 519603 131608
rect 518788 131550 519603 131552
rect 519537 131547 519603 131550
rect 519721 131338 519787 131341
rect 523200 131338 524400 131368
rect 519721 131336 524400 131338
rect 519721 131280 519726 131336
rect 519782 131280 524400 131336
rect 519721 131278 524400 131280
rect 519721 131275 519787 131278
rect 523200 131248 524400 131278
rect 519353 130250 519419 130253
rect 518788 130248 519419 130250
rect 518788 130192 519358 130248
rect 519414 130192 519419 130248
rect 518788 130190 519419 130192
rect 519353 130187 519419 130190
rect 116485 129842 116551 129845
rect 519537 129842 519603 129845
rect 523200 129842 524400 129872
rect 116485 129840 119140 129842
rect 116485 129784 116490 129840
rect 116546 129784 119140 129840
rect 116485 129782 119140 129784
rect 519537 129840 524400 129842
rect 519537 129784 519542 129840
rect 519598 129784 524400 129840
rect 519537 129782 524400 129784
rect 116485 129779 116551 129782
rect 519537 129779 519603 129782
rect 523200 129752 524400 129782
rect 520181 128890 520247 128893
rect 518788 128888 520247 128890
rect 518788 128832 520186 128888
rect 520242 128832 520247 128888
rect 518788 128830 520247 128832
rect 520181 128827 520247 128830
rect 520181 128346 520247 128349
rect 523200 128346 524400 128376
rect 520181 128344 524400 128346
rect 520181 128288 520186 128344
rect 520242 128288 524400 128344
rect 520181 128286 524400 128288
rect 520181 128283 520247 128286
rect 523200 128256 524400 128286
rect 117221 127938 117287 127941
rect 117221 127936 119140 127938
rect 117221 127880 117226 127936
rect 117282 127880 119140 127936
rect 117221 127878 119140 127880
rect 117221 127875 117287 127878
rect 519997 127530 520063 127533
rect 518788 127528 520063 127530
rect 518788 127472 520002 127528
rect 520058 127472 520063 127528
rect 518788 127470 520063 127472
rect 519997 127467 520063 127470
rect 519445 126714 519511 126717
rect 523200 126714 524400 126744
rect 519445 126712 524400 126714
rect 519445 126656 519450 126712
rect 519506 126656 524400 126712
rect 519445 126654 524400 126656
rect 519445 126651 519511 126654
rect 523200 126624 524400 126654
rect 520089 126170 520155 126173
rect 518788 126168 520155 126170
rect 518788 126112 520094 126168
rect 520150 126112 520155 126168
rect 518788 126110 520155 126112
rect 520089 126107 520155 126110
rect 116117 126034 116183 126037
rect 116117 126032 119140 126034
rect 116117 125976 116122 126032
rect 116178 125976 119140 126032
rect 116117 125974 119140 125976
rect 116117 125971 116183 125974
rect 520089 125218 520155 125221
rect 523200 125218 524400 125248
rect 520089 125216 524400 125218
rect 520089 125160 520094 125216
rect 520150 125160 524400 125216
rect 520089 125158 524400 125160
rect 520089 125155 520155 125158
rect 523200 125128 524400 125158
rect 519905 124810 519971 124813
rect 518788 124808 519971 124810
rect 518788 124752 519910 124808
rect 519966 124752 519971 124808
rect 518788 124750 519971 124752
rect 519905 124747 519971 124750
rect 116117 124130 116183 124133
rect 116117 124128 119140 124130
rect 116117 124072 116122 124128
rect 116178 124072 119140 124128
rect 116117 124070 119140 124072
rect 116117 124067 116183 124070
rect 519997 123722 520063 123725
rect 523200 123722 524400 123752
rect 519997 123720 524400 123722
rect 519997 123664 520002 123720
rect 520058 123664 524400 123720
rect 519997 123662 524400 123664
rect 519997 123659 520063 123662
rect 523200 123632 524400 123662
rect 519813 123450 519879 123453
rect 518788 123448 519879 123450
rect 518788 123392 519818 123448
rect 519874 123392 519879 123448
rect 518788 123390 519879 123392
rect 519813 123387 519879 123390
rect 115933 122226 115999 122229
rect 519813 122226 519879 122229
rect 523200 122226 524400 122256
rect 115933 122224 119140 122226
rect 115933 122168 115938 122224
rect 115994 122168 119140 122224
rect 115933 122166 119140 122168
rect 519813 122224 524400 122226
rect 519813 122168 519818 122224
rect 519874 122168 524400 122224
rect 519813 122166 524400 122168
rect 115933 122163 115999 122166
rect 519813 122163 519879 122166
rect 523200 122136 524400 122166
rect 519629 122090 519695 122093
rect 518788 122088 519695 122090
rect 518788 122032 519634 122088
rect 519690 122032 519695 122088
rect 518788 122030 519695 122032
rect 519629 122027 519695 122030
rect 113909 121410 113975 121413
rect 110860 121408 113975 121410
rect 110860 121352 113914 121408
rect 113970 121352 113975 121408
rect 110860 121350 113975 121352
rect 113909 121347 113975 121350
rect 519721 120730 519787 120733
rect 523200 120730 524400 120760
rect 518788 120728 519787 120730
rect 518788 120672 519726 120728
rect 519782 120672 519787 120728
rect 518788 120670 519787 120672
rect 519721 120667 519787 120670
rect 519862 120670 524400 120730
rect 519353 120594 519419 120597
rect 519862 120594 519922 120670
rect 523200 120640 524400 120670
rect 519353 120592 519922 120594
rect 519353 120536 519358 120592
rect 519414 120536 519922 120592
rect 519353 120534 519922 120536
rect 519353 120531 519419 120534
rect 116117 120186 116183 120189
rect 116117 120184 119140 120186
rect 116117 120128 116122 120184
rect 116178 120128 119140 120184
rect 116117 120126 119140 120128
rect 116117 120123 116183 120126
rect 519537 119370 519603 119373
rect 518788 119368 519603 119370
rect 518788 119312 519542 119368
rect 519598 119312 519603 119368
rect 518788 119310 519603 119312
rect 519537 119307 519603 119310
rect 519721 119234 519787 119237
rect 523200 119234 524400 119264
rect 519721 119232 524400 119234
rect 519721 119176 519726 119232
rect 519782 119176 524400 119232
rect 519721 119174 524400 119176
rect 519721 119171 519787 119174
rect 523200 119144 524400 119174
rect 116117 118282 116183 118285
rect 116117 118280 119140 118282
rect 116117 118224 116122 118280
rect 116178 118224 119140 118280
rect 116117 118222 119140 118224
rect 116117 118219 116183 118222
rect 520181 118010 520247 118013
rect 518788 118008 520247 118010
rect 518788 117952 520186 118008
rect 520242 117952 520247 118008
rect 518788 117950 520247 117952
rect 520181 117947 520247 117950
rect 519537 117602 519603 117605
rect 523200 117602 524400 117632
rect 519537 117600 524400 117602
rect 519537 117544 519542 117600
rect 519598 117544 524400 117600
rect 519537 117542 524400 117544
rect 519537 117539 519603 117542
rect 523200 117512 524400 117542
rect 519445 116650 519511 116653
rect 518788 116648 519511 116650
rect 518788 116592 519450 116648
rect 519506 116592 519511 116648
rect 518788 116590 519511 116592
rect 519445 116587 519511 116590
rect 116117 116378 116183 116381
rect 116117 116376 119140 116378
rect 116117 116320 116122 116376
rect 116178 116320 119140 116376
rect 116117 116318 119140 116320
rect 116117 116315 116183 116318
rect 519905 116106 519971 116109
rect 523200 116106 524400 116136
rect 519905 116104 524400 116106
rect 519905 116048 519910 116104
rect 519966 116048 524400 116104
rect 519905 116046 524400 116048
rect 519905 116043 519971 116046
rect 523200 116016 524400 116046
rect 520089 115290 520155 115293
rect 518788 115288 520155 115290
rect 518788 115232 520094 115288
rect 520150 115232 520155 115288
rect 518788 115230 520155 115232
rect 520089 115227 520155 115230
rect 519629 114610 519695 114613
rect 523200 114610 524400 114640
rect 519629 114608 524400 114610
rect 519629 114552 519634 114608
rect 519690 114552 524400 114608
rect 519629 114550 524400 114552
rect 519629 114547 519695 114550
rect 523200 114520 524400 114550
rect 116117 114474 116183 114477
rect 116117 114472 119140 114474
rect 116117 114416 116122 114472
rect 116178 114416 119140 114472
rect 116117 114414 119140 114416
rect 116117 114411 116183 114414
rect 519997 113930 520063 113933
rect 518788 113928 520063 113930
rect 518788 113872 520002 113928
rect 520058 113872 520063 113928
rect 518788 113870 520063 113872
rect 519997 113867 520063 113870
rect 520365 113114 520431 113117
rect 523200 113114 524400 113144
rect 520365 113112 524400 113114
rect 520365 113056 520370 113112
rect 520426 113056 524400 113112
rect 520365 113054 524400 113056
rect 520365 113051 520431 113054
rect 523200 113024 524400 113054
rect 115933 112570 115999 112573
rect 519813 112570 519879 112573
rect 115933 112568 119140 112570
rect 115933 112512 115938 112568
rect 115994 112512 119140 112568
rect 115933 112510 119140 112512
rect 518788 112568 519879 112570
rect 518788 112512 519818 112568
rect 519874 112512 519879 112568
rect 518788 112510 519879 112512
rect 115933 112507 115999 112510
rect 519813 112507 519879 112510
rect 521561 111618 521627 111621
rect 523200 111618 524400 111648
rect 521561 111616 524400 111618
rect 521561 111560 521566 111616
rect 521622 111560 524400 111616
rect 521561 111558 524400 111560
rect 521561 111555 521627 111558
rect 523200 111528 524400 111558
rect 519353 111210 519419 111213
rect 518788 111208 519419 111210
rect 518788 111152 519358 111208
rect 519414 111152 519419 111208
rect 518788 111150 519419 111152
rect 519353 111147 519419 111150
rect 116117 110666 116183 110669
rect 116117 110664 119140 110666
rect 116117 110608 116122 110664
rect 116178 110608 119140 110664
rect 116117 110606 119140 110608
rect 116117 110603 116183 110606
rect 114001 110122 114067 110125
rect 110860 110120 114067 110122
rect 110860 110064 114006 110120
rect 114062 110064 114067 110120
rect 110860 110062 114067 110064
rect 114001 110059 114067 110062
rect 521469 110122 521535 110125
rect 523200 110122 524400 110152
rect 521469 110120 524400 110122
rect 521469 110064 521474 110120
rect 521530 110064 524400 110120
rect 521469 110062 524400 110064
rect 521469 110059 521535 110062
rect 523200 110032 524400 110062
rect 519721 109850 519787 109853
rect 518788 109848 519787 109850
rect 518788 109792 519726 109848
rect 519782 109792 519787 109848
rect 518788 109790 519787 109792
rect 519721 109787 519787 109790
rect 116117 108762 116183 108765
rect 116117 108760 119140 108762
rect 116117 108704 116122 108760
rect 116178 108704 119140 108760
rect 116117 108702 119140 108704
rect 116117 108699 116183 108702
rect 519537 108490 519603 108493
rect 518788 108488 519603 108490
rect 518788 108432 519542 108488
rect 519598 108432 519603 108488
rect 518788 108430 519603 108432
rect 519537 108427 519603 108430
rect 521101 108490 521167 108493
rect 523200 108490 524400 108520
rect 521101 108488 524400 108490
rect 521101 108432 521106 108488
rect 521162 108432 524400 108488
rect 521101 108430 524400 108432
rect 521101 108427 521167 108430
rect 523200 108400 524400 108430
rect 519905 107130 519971 107133
rect 518788 107128 519971 107130
rect 518788 107072 519910 107128
rect 519966 107072 519971 107128
rect 518788 107070 519971 107072
rect 519905 107067 519971 107070
rect 521377 106994 521443 106997
rect 523200 106994 524400 107024
rect 521377 106992 524400 106994
rect 521377 106936 521382 106992
rect 521438 106936 524400 106992
rect 521377 106934 524400 106936
rect 521377 106931 521443 106934
rect 523200 106904 524400 106934
rect 110321 106314 110387 106317
rect 119110 106314 119170 106828
rect 110321 106312 119170 106314
rect 110321 106256 110326 106312
rect 110382 106256 119170 106312
rect 110321 106254 119170 106256
rect 110321 106251 110387 106254
rect 519629 105770 519695 105773
rect 518788 105768 519695 105770
rect 518788 105712 519634 105768
rect 519690 105712 519695 105768
rect 518788 105710 519695 105712
rect 519629 105707 519695 105710
rect 520273 105498 520339 105501
rect 523200 105498 524400 105528
rect 520273 105496 524400 105498
rect 520273 105440 520278 105496
rect 520334 105440 524400 105496
rect 520273 105438 524400 105440
rect 520273 105435 520339 105438
rect 523200 105408 524400 105438
rect 117129 104818 117195 104821
rect 117129 104816 119140 104818
rect 117129 104760 117134 104816
rect 117190 104760 119140 104816
rect 117129 104758 119140 104760
rect 117129 104755 117195 104758
rect 520365 104410 520431 104413
rect 518788 104408 520431 104410
rect 518788 104352 520370 104408
rect 520426 104352 520431 104408
rect 518788 104350 520431 104352
rect 520365 104347 520431 104350
rect 520917 104002 520983 104005
rect 523200 104002 524400 104032
rect 520917 104000 524400 104002
rect 520917 103944 520922 104000
rect 520978 103944 524400 104000
rect 520917 103942 524400 103944
rect 520917 103939 520983 103942
rect 523200 103912 524400 103942
rect 521561 103050 521627 103053
rect 518788 103048 521627 103050
rect 518788 102992 521566 103048
rect 521622 102992 521627 103048
rect 518788 102990 521627 102992
rect 521561 102987 521627 102990
rect 116945 102914 117011 102917
rect 116945 102912 119140 102914
rect 116945 102856 116950 102912
rect 117006 102856 119140 102912
rect 116945 102854 119140 102856
rect 116945 102851 117011 102854
rect 521009 102506 521075 102509
rect 523200 102506 524400 102536
rect 521009 102504 524400 102506
rect 521009 102448 521014 102504
rect 521070 102448 524400 102504
rect 521009 102446 524400 102448
rect 521009 102443 521075 102446
rect 523200 102416 524400 102446
rect 521469 101690 521535 101693
rect 518788 101688 521535 101690
rect 518788 101632 521474 101688
rect 521530 101632 521535 101688
rect 518788 101630 521535 101632
rect 521469 101627 521535 101630
rect 117037 101010 117103 101013
rect 521193 101010 521259 101013
rect 523200 101010 524400 101040
rect 117037 101008 119140 101010
rect 117037 100952 117042 101008
rect 117098 100952 119140 101008
rect 117037 100950 119140 100952
rect 521193 101008 524400 101010
rect 521193 100952 521198 101008
rect 521254 100952 524400 101008
rect 521193 100950 524400 100952
rect 117037 100947 117103 100950
rect 521193 100947 521259 100950
rect 523200 100920 524400 100950
rect 521101 100330 521167 100333
rect 518788 100328 521167 100330
rect 518788 100272 521106 100328
rect 521162 100272 521167 100328
rect 518788 100270 521167 100272
rect 521101 100267 521167 100270
rect 519629 99378 519695 99381
rect 523200 99378 524400 99408
rect 519629 99376 524400 99378
rect 519629 99320 519634 99376
rect 519690 99320 524400 99376
rect 519629 99318 524400 99320
rect 519629 99315 519695 99318
rect 523200 99288 524400 99318
rect 116853 99106 116919 99109
rect 116853 99104 119140 99106
rect 116853 99048 116858 99104
rect 116914 99048 119140 99104
rect 116853 99046 119140 99048
rect 116853 99043 116919 99046
rect 521377 98970 521443 98973
rect 518788 98968 521443 98970
rect 518788 98912 521382 98968
rect 521438 98912 521443 98968
rect 518788 98910 521443 98912
rect 521377 98907 521443 98910
rect 114093 98698 114159 98701
rect 110860 98696 114159 98698
rect 110860 98640 114098 98696
rect 114154 98640 114159 98696
rect 110860 98638 114159 98640
rect 114093 98635 114159 98638
rect 519721 97882 519787 97885
rect 523200 97882 524400 97912
rect 519721 97880 524400 97882
rect 519721 97824 519726 97880
rect 519782 97824 524400 97880
rect 519721 97822 524400 97824
rect 519721 97819 519787 97822
rect 523200 97792 524400 97822
rect 520273 97610 520339 97613
rect 518788 97608 520339 97610
rect 518788 97552 520278 97608
rect 520334 97552 520339 97608
rect 518788 97550 520339 97552
rect 520273 97547 520339 97550
rect 116761 97202 116827 97205
rect 116761 97200 119140 97202
rect 116761 97144 116766 97200
rect 116822 97144 119140 97200
rect 116761 97142 119140 97144
rect 116761 97139 116827 97142
rect 519261 96386 519327 96389
rect 523200 96386 524400 96416
rect 519261 96384 524400 96386
rect 519261 96328 519266 96384
rect 519322 96328 524400 96384
rect 519261 96326 524400 96328
rect 519261 96323 519327 96326
rect 523200 96296 524400 96326
rect 520917 96250 520983 96253
rect 518788 96248 520983 96250
rect 518788 96192 520922 96248
rect 520978 96192 520983 96248
rect 518788 96190 520983 96192
rect 520917 96187 520983 96190
rect 116669 95298 116735 95301
rect 116669 95296 119140 95298
rect 116669 95240 116674 95296
rect 116730 95240 119140 95296
rect 116669 95238 119140 95240
rect 116669 95235 116735 95238
rect 521009 95026 521075 95029
rect 518758 95024 521075 95026
rect 518758 94968 521014 95024
rect 521070 94968 521075 95024
rect 518758 94966 521075 94968
rect 518758 94860 518818 94966
rect 521009 94963 521075 94966
rect 519997 94890 520063 94893
rect 523200 94890 524400 94920
rect 519997 94888 524400 94890
rect 519997 94832 520002 94888
rect 520058 94832 524400 94888
rect 519997 94830 524400 94832
rect 519997 94827 520063 94830
rect 523200 94800 524400 94830
rect 521193 93530 521259 93533
rect 518788 93528 521259 93530
rect 518788 93472 521198 93528
rect 521254 93472 521259 93528
rect 518788 93470 521259 93472
rect 521193 93467 521259 93470
rect 116577 93394 116643 93397
rect 520181 93394 520247 93397
rect 523200 93394 524400 93424
rect 116577 93392 119140 93394
rect 116577 93336 116582 93392
rect 116638 93336 119140 93392
rect 116577 93334 119140 93336
rect 520181 93392 524400 93394
rect 520181 93336 520186 93392
rect 520242 93336 524400 93392
rect 520181 93334 524400 93336
rect 116577 93331 116643 93334
rect 520181 93331 520247 93334
rect 523200 93304 524400 93334
rect 519629 92170 519695 92173
rect 518788 92168 519695 92170
rect 518788 92112 519634 92168
rect 519690 92112 519695 92168
rect 518788 92110 519695 92112
rect 519629 92107 519695 92110
rect 521285 91898 521351 91901
rect 523200 91898 524400 91928
rect 521285 91896 524400 91898
rect 521285 91840 521290 91896
rect 521346 91840 524400 91896
rect 521285 91838 524400 91840
rect 521285 91835 521351 91838
rect 523200 91808 524400 91838
rect 116117 91354 116183 91357
rect 116117 91352 119140 91354
rect 116117 91296 116122 91352
rect 116178 91296 119140 91352
rect 116117 91294 119140 91296
rect 116117 91291 116183 91294
rect 519721 90810 519787 90813
rect 518788 90808 519787 90810
rect 518788 90752 519726 90808
rect 519782 90752 519787 90808
rect 518788 90750 519787 90752
rect 519721 90747 519787 90750
rect 520917 90266 520983 90269
rect 523200 90266 524400 90296
rect 520917 90264 524400 90266
rect 520917 90208 520922 90264
rect 520978 90208 524400 90264
rect 520917 90206 524400 90208
rect 520917 90203 520983 90206
rect 523200 90176 524400 90206
rect 116117 89450 116183 89453
rect 519261 89450 519327 89453
rect 116117 89448 119140 89450
rect 116117 89392 116122 89448
rect 116178 89392 119140 89448
rect 116117 89390 119140 89392
rect 518788 89448 519327 89450
rect 518788 89392 519266 89448
rect 519322 89392 519327 89448
rect 518788 89390 519327 89392
rect 116117 89387 116183 89390
rect 519261 89387 519327 89390
rect 521377 88770 521443 88773
rect 523200 88770 524400 88800
rect 521377 88768 524400 88770
rect 521377 88712 521382 88768
rect 521438 88712 524400 88768
rect 521377 88710 524400 88712
rect 521377 88707 521443 88710
rect 523200 88680 524400 88710
rect 519997 88090 520063 88093
rect 518788 88088 520063 88090
rect 518788 88032 520002 88088
rect 520058 88032 520063 88088
rect 518788 88030 520063 88032
rect 519997 88027 520063 88030
rect 116025 87546 116091 87549
rect 116025 87544 119140 87546
rect 116025 87488 116030 87544
rect 116086 87488 119140 87544
rect 116025 87486 119140 87488
rect 116025 87483 116091 87486
rect 114185 87274 114251 87277
rect 110860 87272 114251 87274
rect 110860 87216 114190 87272
rect 114246 87216 114251 87272
rect 110860 87214 114251 87216
rect 114185 87211 114251 87214
rect 521009 87274 521075 87277
rect 523200 87274 524400 87304
rect 521009 87272 524400 87274
rect 521009 87216 521014 87272
rect 521070 87216 524400 87272
rect 521009 87214 524400 87216
rect 521009 87211 521075 87214
rect 523200 87184 524400 87214
rect 520181 86730 520247 86733
rect 518788 86728 520247 86730
rect 518788 86672 520186 86728
rect 520242 86672 520247 86728
rect 518788 86670 520247 86672
rect 520181 86667 520247 86670
rect 520273 85778 520339 85781
rect 523200 85778 524400 85808
rect 520273 85776 524400 85778
rect 520273 85720 520278 85776
rect 520334 85720 524400 85776
rect 520273 85718 524400 85720
rect 520273 85715 520339 85718
rect 523200 85688 524400 85718
rect 115197 85642 115263 85645
rect 115197 85640 119140 85642
rect 115197 85584 115202 85640
rect 115258 85584 119140 85640
rect 115197 85582 119140 85584
rect 115197 85579 115263 85582
rect 521193 84282 521259 84285
rect 523200 84282 524400 84312
rect 521193 84280 524400 84282
rect 521193 84224 521198 84280
rect 521254 84224 524400 84280
rect 521193 84222 524400 84224
rect 521193 84219 521259 84222
rect 523200 84192 524400 84222
rect 521285 84010 521351 84013
rect 518788 84008 521351 84010
rect 518788 83952 521290 84008
rect 521346 83952 521351 84008
rect 518788 83950 521351 83952
rect 521285 83947 521351 83950
rect 116577 83738 116643 83741
rect 116577 83736 119140 83738
rect 116577 83680 116582 83736
rect 116638 83680 119140 83736
rect 116577 83678 119140 83680
rect 116577 83675 116643 83678
rect 519997 82786 520063 82789
rect 523200 82786 524400 82816
rect 519997 82784 524400 82786
rect 519997 82728 520002 82784
rect 520058 82728 524400 82784
rect 519997 82726 524400 82728
rect 519997 82723 520063 82726
rect 523200 82696 524400 82726
rect 520917 82650 520983 82653
rect 518788 82648 520983 82650
rect 518788 82592 520922 82648
rect 520978 82592 520983 82648
rect 518788 82590 520983 82592
rect 520917 82587 520983 82590
rect 116209 81834 116275 81837
rect 116209 81832 119140 81834
rect 116209 81776 116214 81832
rect 116270 81776 119140 81832
rect 116209 81774 119140 81776
rect 116209 81771 116275 81774
rect 521377 81290 521443 81293
rect 518788 81288 521443 81290
rect 518788 81232 521382 81288
rect 521438 81232 521443 81288
rect 518788 81230 521443 81232
rect 521377 81227 521443 81230
rect 520181 81154 520247 81157
rect 523200 81154 524400 81184
rect 520181 81152 524400 81154
rect 520181 81096 520186 81152
rect 520242 81096 524400 81152
rect 520181 81094 524400 81096
rect 520181 81091 520247 81094
rect 523200 81064 524400 81094
rect 115933 79930 115999 79933
rect 521009 79930 521075 79933
rect 115933 79928 119140 79930
rect 115933 79872 115938 79928
rect 115994 79872 119140 79928
rect 115933 79870 119140 79872
rect 518788 79928 521075 79930
rect 518788 79872 521014 79928
rect 521070 79872 521075 79928
rect 518788 79870 521075 79872
rect 115933 79867 115999 79870
rect 521009 79867 521075 79870
rect 519629 79658 519695 79661
rect 523200 79658 524400 79688
rect 519629 79656 524400 79658
rect 519629 79600 519634 79656
rect 519690 79600 524400 79656
rect 519629 79598 524400 79600
rect 519629 79595 519695 79598
rect 523200 79568 524400 79598
rect 520273 78570 520339 78573
rect 518788 78568 520339 78570
rect 518788 78512 520278 78568
rect 520334 78512 520339 78568
rect 518788 78510 520339 78512
rect 520273 78507 520339 78510
rect 519721 78162 519787 78165
rect 523200 78162 524400 78192
rect 519721 78160 524400 78162
rect 519721 78104 519726 78160
rect 519782 78104 524400 78160
rect 519721 78102 524400 78104
rect 519721 78099 519787 78102
rect 523200 78072 524400 78102
rect 116117 78026 116183 78029
rect 116117 78024 119140 78026
rect 116117 77968 116122 78024
rect 116178 77968 119140 78024
rect 116117 77966 119140 77968
rect 116117 77963 116183 77966
rect 521193 77210 521259 77213
rect 518788 77208 521259 77210
rect 518788 77152 521198 77208
rect 521254 77152 521259 77208
rect 518788 77150 521259 77152
rect 521193 77147 521259 77150
rect 520089 76666 520155 76669
rect 523200 76666 524400 76696
rect 520089 76664 524400 76666
rect 520089 76608 520094 76664
rect 520150 76608 524400 76664
rect 520089 76606 524400 76608
rect 520089 76603 520155 76606
rect 523200 76576 524400 76606
rect 519997 75986 520063 75989
rect 110860 75926 119140 75986
rect 518788 75984 520063 75986
rect 518788 75928 520002 75984
rect 520058 75928 520063 75984
rect 518788 75926 520063 75928
rect 519997 75923 520063 75926
rect 519997 75170 520063 75173
rect 523200 75170 524400 75200
rect 519997 75168 524400 75170
rect 519997 75112 520002 75168
rect 520058 75112 524400 75168
rect 519997 75110 524400 75112
rect 519997 75107 520063 75110
rect 523200 75080 524400 75110
rect 520181 74626 520247 74629
rect 518788 74624 520247 74626
rect 518788 74568 520186 74624
rect 520242 74568 520247 74624
rect 518788 74566 520247 74568
rect 520181 74563 520247 74566
rect 116669 74082 116735 74085
rect 116669 74080 119140 74082
rect 116669 74024 116674 74080
rect 116730 74024 119140 74080
rect 116669 74022 119140 74024
rect 116669 74019 116735 74022
rect 519261 73674 519327 73677
rect 523200 73674 524400 73704
rect 519261 73672 524400 73674
rect 519261 73616 519266 73672
rect 519322 73616 524400 73672
rect 519261 73614 524400 73616
rect 519261 73611 519327 73614
rect 523200 73584 524400 73614
rect 519629 73266 519695 73269
rect 518788 73264 519695 73266
rect 518788 73208 519634 73264
rect 519690 73208 519695 73264
rect 518788 73206 519695 73208
rect 519629 73203 519695 73206
rect 519721 72450 519787 72453
rect 518758 72448 519787 72450
rect 518758 72392 519726 72448
rect 519782 72392 519787 72448
rect 518758 72390 519787 72392
rect 116577 72178 116643 72181
rect 116577 72176 119140 72178
rect 116577 72120 116582 72176
rect 116638 72120 119140 72176
rect 116577 72118 119140 72120
rect 116577 72115 116643 72118
rect 518758 71876 518818 72390
rect 519721 72387 519787 72390
rect 519445 72042 519511 72045
rect 523200 72042 524400 72072
rect 519445 72040 524400 72042
rect 519445 71984 519450 72040
rect 519506 71984 524400 72040
rect 519445 71982 524400 71984
rect 519445 71979 519511 71982
rect 523200 71952 524400 71982
rect 520089 70546 520155 70549
rect 523200 70546 524400 70576
rect 518788 70544 520155 70546
rect 518788 70488 520094 70544
rect 520150 70488 520155 70544
rect 518788 70486 520155 70488
rect 520089 70483 520155 70486
rect 520230 70486 524400 70546
rect 520230 70413 520290 70486
rect 523200 70456 524400 70486
rect 520181 70408 520290 70413
rect 520181 70352 520186 70408
rect 520242 70352 520290 70408
rect 520181 70350 520290 70352
rect 520181 70347 520247 70350
rect 116301 70274 116367 70277
rect 116301 70272 119140 70274
rect 116301 70216 116306 70272
rect 116362 70216 119140 70272
rect 116301 70214 119140 70216
rect 116301 70211 116367 70214
rect 519997 69186 520063 69189
rect 518788 69184 520063 69186
rect 518788 69128 520002 69184
rect 520058 69128 520063 69184
rect 518788 69126 520063 69128
rect 519997 69123 520063 69126
rect 519629 69050 519695 69053
rect 523200 69050 524400 69080
rect 519629 69048 524400 69050
rect 519629 68992 519634 69048
rect 519690 68992 524400 69048
rect 519629 68990 524400 68992
rect 519629 68987 519695 68990
rect 523200 68960 524400 68990
rect 116117 68370 116183 68373
rect 116117 68368 119140 68370
rect 116117 68312 116122 68368
rect 116178 68312 119140 68368
rect 116117 68310 119140 68312
rect 116117 68307 116183 68310
rect 519261 67826 519327 67829
rect 518788 67824 519327 67826
rect 518788 67768 519266 67824
rect 519322 67768 519327 67824
rect 518788 67766 519327 67768
rect 519261 67763 519327 67766
rect 519261 67554 519327 67557
rect 523200 67554 524400 67584
rect 519261 67552 524400 67554
rect 519261 67496 519266 67552
rect 519322 67496 524400 67552
rect 519261 67494 524400 67496
rect 519261 67491 519327 67494
rect 523200 67464 524400 67494
rect 116577 66466 116643 66469
rect 519445 66466 519511 66469
rect 116577 66464 119140 66466
rect 116577 66408 116582 66464
rect 116638 66408 119140 66464
rect 116577 66406 119140 66408
rect 518788 66464 519511 66466
rect 518788 66408 519450 66464
rect 519506 66408 519511 66464
rect 518788 66406 519511 66408
rect 116577 66403 116643 66406
rect 519445 66403 519511 66406
rect 519813 66058 519879 66061
rect 523200 66058 524400 66088
rect 519813 66056 524400 66058
rect 519813 66000 519818 66056
rect 519874 66000 524400 66056
rect 519813 65998 524400 66000
rect 519813 65995 519879 65998
rect 523200 65968 524400 65998
rect 520181 65106 520247 65109
rect 518788 65104 520247 65106
rect 518788 65048 520186 65104
rect 520242 65048 520247 65104
rect 518788 65046 520247 65048
rect 520181 65043 520247 65046
rect 113357 64562 113423 64565
rect 110860 64560 113423 64562
rect 110860 64504 113362 64560
rect 113418 64504 113423 64560
rect 110860 64502 113423 64504
rect 113357 64499 113423 64502
rect 116209 64562 116275 64565
rect 521101 64562 521167 64565
rect 523200 64562 524400 64592
rect 116209 64560 119140 64562
rect 116209 64504 116214 64560
rect 116270 64504 119140 64560
rect 116209 64502 119140 64504
rect 521101 64560 524400 64562
rect 521101 64504 521106 64560
rect 521162 64504 524400 64560
rect 521101 64502 524400 64504
rect 116209 64499 116275 64502
rect 521101 64499 521167 64502
rect 523200 64472 524400 64502
rect 519629 63746 519695 63749
rect 518788 63744 519695 63746
rect 518788 63688 519634 63744
rect 519690 63688 519695 63744
rect 518788 63686 519695 63688
rect 519629 63683 519695 63686
rect 520733 62930 520799 62933
rect 523200 62930 524400 62960
rect 520733 62928 524400 62930
rect 520733 62872 520738 62928
rect 520794 62872 524400 62928
rect 520733 62870 524400 62872
rect 520733 62867 520799 62870
rect 523200 62840 524400 62870
rect 116117 62658 116183 62661
rect 116117 62656 119140 62658
rect 116117 62600 116122 62656
rect 116178 62600 119140 62656
rect 116117 62598 119140 62600
rect 116117 62595 116183 62598
rect 521101 62386 521167 62389
rect 518788 62384 521167 62386
rect 518788 62328 521106 62384
rect 521162 62328 521167 62384
rect 518788 62326 521167 62328
rect 521101 62323 521167 62326
rect 520273 61434 520339 61437
rect 523200 61434 524400 61464
rect 520273 61432 524400 61434
rect 520273 61376 520278 61432
rect 520334 61376 524400 61432
rect 520273 61374 524400 61376
rect 520273 61371 520339 61374
rect 523200 61344 524400 61374
rect 519261 61026 519327 61029
rect 518788 61024 519327 61026
rect 518788 60968 519266 61024
rect 519322 60968 519327 61024
rect 518788 60966 519327 60968
rect 519261 60963 519327 60966
rect 116577 60618 116643 60621
rect 116577 60616 119140 60618
rect 116577 60560 116582 60616
rect 116638 60560 119140 60616
rect 116577 60558 119140 60560
rect 116577 60555 116643 60558
rect 521009 59938 521075 59941
rect 523200 59938 524400 59968
rect 521009 59936 524400 59938
rect 521009 59880 521014 59936
rect 521070 59880 524400 59936
rect 521009 59878 524400 59880
rect 521009 59875 521075 59878
rect 523200 59848 524400 59878
rect 519813 59666 519879 59669
rect 518788 59664 519879 59666
rect 518788 59608 519818 59664
rect 519874 59608 519879 59664
rect 518788 59606 519879 59608
rect 519813 59603 519879 59606
rect 110321 58034 110387 58037
rect 119110 58034 119170 58684
rect 521101 58442 521167 58445
rect 523200 58442 524400 58472
rect 521101 58440 524400 58442
rect 521101 58384 521106 58440
rect 521162 58384 524400 58440
rect 521101 58382 524400 58384
rect 521101 58379 521167 58382
rect 523200 58352 524400 58382
rect 520733 58306 520799 58309
rect 518788 58304 520799 58306
rect 518788 58248 520738 58304
rect 520794 58248 520799 58304
rect 518788 58246 520799 58248
rect 520733 58243 520799 58246
rect 110321 58032 119170 58034
rect 110321 57976 110326 58032
rect 110382 57976 119170 58032
rect 110321 57974 119170 57976
rect 110321 57971 110387 57974
rect 520181 56946 520247 56949
rect 518788 56944 520247 56946
rect 518788 56888 520186 56944
rect 520242 56888 520247 56944
rect 518788 56886 520247 56888
rect 520181 56883 520247 56886
rect 520365 56946 520431 56949
rect 523200 56946 524400 56976
rect 520365 56944 524400 56946
rect 520365 56888 520370 56944
rect 520426 56888 524400 56944
rect 520365 56886 524400 56888
rect 520365 56883 520431 56886
rect 523200 56856 524400 56886
rect 110321 56810 110387 56813
rect 110321 56808 119140 56810
rect 110321 56752 110326 56808
rect 110382 56752 119140 56808
rect 110321 56750 119140 56752
rect 110321 56747 110387 56750
rect 521009 55586 521075 55589
rect 518788 55584 521075 55586
rect 518788 55528 521014 55584
rect 521070 55528 521075 55584
rect 518788 55526 521075 55528
rect 521009 55523 521075 55526
rect 520273 55450 520339 55453
rect 523200 55450 524400 55480
rect 520273 55448 524400 55450
rect 520273 55392 520278 55448
rect 520334 55392 524400 55448
rect 520273 55390 524400 55392
rect 520273 55387 520339 55390
rect 523200 55360 524400 55390
rect 110321 53954 110387 53957
rect 119110 53954 119170 54876
rect 521101 54226 521167 54229
rect 518788 54224 521167 54226
rect 518788 54168 521106 54224
rect 521162 54168 521167 54224
rect 518788 54166 521167 54168
rect 521101 54163 521167 54166
rect 110321 53952 119170 53954
rect 110321 53896 110326 53952
rect 110382 53896 119170 53952
rect 110321 53894 119170 53896
rect 110321 53891 110387 53894
rect 519261 53818 519327 53821
rect 523200 53818 524400 53848
rect 519261 53816 524400 53818
rect 519261 53760 519266 53816
rect 519322 53760 524400 53816
rect 519261 53758 524400 53760
rect 519261 53755 519327 53758
rect 523200 53728 524400 53758
rect 114185 53138 114251 53141
rect 110860 53136 114251 53138
rect 110860 53080 114190 53136
rect 114246 53080 114251 53136
rect 110860 53078 114251 53080
rect 114185 53075 114251 53078
rect 110321 52594 110387 52597
rect 119110 52594 119170 52972
rect 520365 52866 520431 52869
rect 518788 52864 520431 52866
rect 518788 52808 520370 52864
rect 520426 52808 520431 52864
rect 518788 52806 520431 52808
rect 520365 52803 520431 52806
rect 110321 52592 119170 52594
rect 110321 52536 110326 52592
rect 110382 52536 119170 52592
rect 110321 52534 119170 52536
rect 110321 52531 110387 52534
rect 520089 52322 520155 52325
rect 523200 52322 524400 52352
rect 520089 52320 524400 52322
rect 520089 52264 520094 52320
rect 520150 52264 524400 52320
rect 520089 52262 524400 52264
rect 520089 52259 520155 52262
rect 523200 52232 524400 52262
rect 520273 51506 520339 51509
rect 518788 51504 520339 51506
rect 518788 51448 520278 51504
rect 520334 51448 520339 51504
rect 518788 51446 520339 51448
rect 520273 51443 520339 51446
rect 110321 51098 110387 51101
rect 110321 51096 119140 51098
rect 110321 51040 110326 51096
rect 110382 51040 119140 51096
rect 110321 51038 119140 51040
rect 110321 51035 110387 51038
rect 519997 50826 520063 50829
rect 523200 50826 524400 50856
rect 519997 50824 524400 50826
rect 519997 50768 520002 50824
rect 520058 50768 524400 50824
rect 519997 50766 524400 50768
rect 519997 50763 520063 50766
rect 523200 50736 524400 50766
rect 519261 50146 519327 50149
rect 518788 50144 519327 50146
rect 518788 50088 519266 50144
rect 519322 50088 519327 50144
rect 518788 50086 519327 50088
rect 519261 50083 519327 50086
rect 520181 49330 520247 49333
rect 523200 49330 524400 49360
rect 520181 49328 524400 49330
rect 520181 49272 520186 49328
rect 520242 49272 524400 49328
rect 520181 49270 524400 49272
rect 520181 49267 520247 49270
rect 523200 49240 524400 49270
rect 110321 48378 110387 48381
rect 119110 48378 119170 49164
rect 520089 48786 520155 48789
rect 518788 48784 520155 48786
rect 518788 48728 520094 48784
rect 520150 48728 520155 48784
rect 518788 48726 520155 48728
rect 520089 48723 520155 48726
rect 110321 48376 119170 48378
rect 110321 48320 110326 48376
rect 110382 48320 119170 48376
rect 110321 48318 119170 48320
rect 110321 48315 110387 48318
rect 519445 47834 519511 47837
rect 523200 47834 524400 47864
rect 519445 47832 524400 47834
rect 519445 47776 519450 47832
rect 519506 47776 524400 47832
rect 519445 47774 524400 47776
rect 519445 47771 519511 47774
rect 523200 47744 524400 47774
rect 519997 47426 520063 47429
rect 518788 47424 520063 47426
rect 518788 47368 520002 47424
rect 520058 47368 520063 47424
rect 518788 47366 520063 47368
rect 519997 47363 520063 47366
rect 110321 47154 110387 47157
rect 110321 47152 119140 47154
rect 110321 47096 110326 47152
rect 110382 47096 119140 47152
rect 110321 47094 119140 47096
rect 110321 47091 110387 47094
rect 519905 46338 519971 46341
rect 523200 46338 524400 46368
rect 519905 46336 524400 46338
rect 519905 46280 519910 46336
rect 519966 46280 524400 46336
rect 519905 46278 524400 46280
rect 519905 46275 519971 46278
rect 523200 46248 524400 46278
rect 520181 46066 520247 46069
rect 518788 46064 520247 46066
rect 518788 46008 520186 46064
rect 520242 46008 520247 46064
rect 518788 46006 520247 46008
rect 520181 46003 520247 46006
rect 111057 44298 111123 44301
rect 119110 44298 119170 45220
rect 519445 44706 519511 44709
rect 518788 44704 519511 44706
rect 518788 44648 519450 44704
rect 519506 44648 519511 44704
rect 518788 44646 519511 44648
rect 519445 44643 519511 44646
rect 519813 44706 519879 44709
rect 523200 44706 524400 44736
rect 519813 44704 524400 44706
rect 519813 44648 519818 44704
rect 519874 44648 524400 44704
rect 519813 44646 524400 44648
rect 519813 44643 519879 44646
rect 523200 44616 524400 44646
rect 111057 44296 119170 44298
rect 111057 44240 111062 44296
rect 111118 44240 119170 44296
rect 111057 44238 119170 44240
rect 111057 44235 111123 44238
rect 116117 43346 116183 43349
rect 519905 43346 519971 43349
rect 116117 43344 119140 43346
rect 116117 43288 116122 43344
rect 116178 43288 119140 43344
rect 116117 43286 119140 43288
rect 518788 43344 519971 43346
rect 518788 43288 519910 43344
rect 519966 43288 519971 43344
rect 518788 43286 519971 43288
rect 116117 43283 116183 43286
rect 519905 43283 519971 43286
rect 520181 43210 520247 43213
rect 523200 43210 524400 43240
rect 520181 43208 524400 43210
rect 520181 43152 520186 43208
rect 520242 43152 524400 43208
rect 520181 43150 524400 43152
rect 520181 43147 520247 43150
rect 523200 43120 524400 43150
rect 110321 42938 110387 42941
rect 110873 42938 110939 42941
rect 110321 42936 110939 42938
rect 110321 42880 110326 42936
rect 110382 42880 110878 42936
rect 110934 42880 110939 42936
rect 110321 42878 110939 42880
rect 110321 42875 110387 42878
rect 110873 42875 110939 42878
rect 110321 42394 110387 42397
rect 110689 42394 110755 42397
rect 110321 42392 110755 42394
rect 110321 42336 110326 42392
rect 110382 42336 110694 42392
rect 110750 42336 110755 42392
rect 110321 42334 110755 42336
rect 110321 42331 110387 42334
rect 110689 42331 110755 42334
rect 519813 41986 519879 41989
rect 518788 41984 519879 41986
rect 518788 41928 519818 41984
rect 519874 41928 519879 41984
rect 518788 41926 519879 41928
rect 519813 41923 519879 41926
rect 114093 41850 114159 41853
rect 110860 41848 114159 41850
rect 110860 41792 114098 41848
rect 114154 41792 114159 41848
rect 110860 41790 114159 41792
rect 114093 41787 114159 41790
rect 520089 41714 520155 41717
rect 523200 41714 524400 41744
rect 520089 41712 524400 41714
rect 520089 41656 520094 41712
rect 520150 41656 524400 41712
rect 520089 41654 524400 41656
rect 520089 41651 520155 41654
rect 523200 41624 524400 41654
rect 110597 41442 110663 41445
rect 110597 41440 119140 41442
rect 110597 41384 110602 41440
rect 110658 41384 119140 41440
rect 110597 41382 119140 41384
rect 110597 41379 110663 41382
rect 520181 40626 520247 40629
rect 518788 40624 520247 40626
rect 518788 40568 520186 40624
rect 520242 40568 520247 40624
rect 518788 40566 520247 40568
rect 520181 40563 520247 40566
rect 520181 40218 520247 40221
rect 523200 40218 524400 40248
rect 520181 40216 524400 40218
rect 520181 40160 520186 40216
rect 520242 40160 524400 40216
rect 520181 40158 524400 40160
rect 520181 40155 520247 40158
rect 523200 40128 524400 40158
rect 116761 39538 116827 39541
rect 116761 39536 119140 39538
rect 116761 39480 116766 39536
rect 116822 39480 119140 39536
rect 116761 39478 119140 39480
rect 116761 39475 116827 39478
rect 520089 39266 520155 39269
rect 518788 39264 520155 39266
rect 518788 39208 520094 39264
rect 520150 39208 520155 39264
rect 518788 39206 520155 39208
rect 520089 39203 520155 39206
rect 519813 38722 519879 38725
rect 523200 38722 524400 38752
rect 519813 38720 524400 38722
rect 519813 38664 519818 38720
rect 519874 38664 524400 38720
rect 519813 38662 524400 38664
rect 519813 38659 519879 38662
rect 523200 38632 524400 38662
rect 520181 37906 520247 37909
rect 518788 37904 520247 37906
rect 518788 37848 520186 37904
rect 520242 37848 520247 37904
rect 518788 37846 520247 37848
rect 520181 37843 520247 37846
rect 116669 37634 116735 37637
rect 116669 37632 119140 37634
rect 116669 37576 116674 37632
rect 116730 37576 119140 37632
rect 116669 37574 119140 37576
rect 116669 37571 116735 37574
rect 521561 37226 521627 37229
rect 523200 37226 524400 37256
rect 521561 37224 524400 37226
rect 521561 37168 521566 37224
rect 521622 37168 524400 37224
rect 521561 37166 524400 37168
rect 521561 37163 521627 37166
rect 523200 37136 524400 37166
rect 519813 36546 519879 36549
rect 518788 36544 519879 36546
rect 518788 36488 519818 36544
rect 519874 36488 519879 36544
rect 518788 36486 519879 36488
rect 519813 36483 519879 36486
rect 521561 36002 521627 36005
rect 521561 36000 521670 36002
rect 521561 35944 521566 36000
rect 521622 35944 521670 36000
rect 521561 35939 521670 35944
rect 521610 35866 521670 35939
rect 518758 35806 521670 35866
rect 110413 35050 110479 35053
rect 110965 35050 111031 35053
rect 110413 35048 111031 35050
rect 110413 34992 110418 35048
rect 110474 34992 110970 35048
rect 111026 34992 111031 35048
rect 110413 34990 111031 34992
rect 110413 34987 110479 34990
rect 110965 34987 111031 34990
rect 110321 34778 110387 34781
rect 111241 34778 111307 34781
rect 110321 34776 111307 34778
rect 110321 34720 110326 34776
rect 110382 34720 111246 34776
rect 111302 34720 111307 34776
rect 110321 34718 111307 34720
rect 110321 34715 110387 34718
rect 111241 34715 111307 34718
rect 110321 34642 110387 34645
rect 110597 34642 110663 34645
rect 110321 34640 110663 34642
rect 110321 34584 110326 34640
rect 110382 34584 110602 34640
rect 110658 34584 110663 34640
rect 110321 34582 110663 34584
rect 110321 34579 110387 34582
rect 110597 34579 110663 34582
rect 111149 34642 111215 34645
rect 119110 34642 119170 35700
rect 518758 35156 518818 35806
rect 521101 35594 521167 35597
rect 523200 35594 524400 35624
rect 521101 35592 524400 35594
rect 521101 35536 521106 35592
rect 521162 35536 524400 35592
rect 521101 35534 524400 35536
rect 521101 35531 521167 35534
rect 523200 35504 524400 35534
rect 111149 34640 119170 34642
rect 111149 34584 111154 34640
rect 111210 34584 119170 34640
rect 111149 34582 119170 34584
rect 111149 34579 111215 34582
rect 521101 34506 521167 34509
rect 518758 34504 521167 34506
rect 518758 34448 521106 34504
rect 521162 34448 521167 34504
rect 518758 34446 521167 34448
rect 116945 33826 117011 33829
rect 116945 33824 119140 33826
rect 116945 33768 116950 33824
rect 117006 33768 119140 33824
rect 518758 33796 518818 34446
rect 521101 34443 521167 34446
rect 520917 34098 520983 34101
rect 523200 34098 524400 34128
rect 520917 34096 524400 34098
rect 520917 34040 520922 34096
rect 520978 34040 524400 34096
rect 520917 34038 524400 34040
rect 520917 34035 520983 34038
rect 523200 34008 524400 34038
rect 116945 33766 119140 33768
rect 116945 33763 117011 33766
rect 520917 33146 520983 33149
rect 518758 33144 520983 33146
rect 518758 33088 520922 33144
rect 520978 33088 520983 33144
rect 518758 33086 520983 33088
rect 518758 32436 518818 33086
rect 520917 33083 520983 33086
rect 520917 32602 520983 32605
rect 523200 32602 524400 32632
rect 520917 32600 524400 32602
rect 520917 32544 520922 32600
rect 520978 32544 524400 32600
rect 520917 32542 524400 32544
rect 520917 32539 520983 32542
rect 523200 32512 524400 32542
rect 116853 31786 116919 31789
rect 116853 31784 119140 31786
rect 116853 31728 116858 31784
rect 116914 31728 119140 31784
rect 116853 31726 119140 31728
rect 116853 31723 116919 31726
rect 520917 31650 520983 31653
rect 518758 31648 520983 31650
rect 518758 31592 520922 31648
rect 520978 31592 520983 31648
rect 518758 31590 520983 31592
rect 518758 31076 518818 31590
rect 520917 31587 520983 31590
rect 520917 31106 520983 31109
rect 523200 31106 524400 31136
rect 520917 31104 524400 31106
rect 520917 31048 520922 31104
rect 520978 31048 524400 31104
rect 520917 31046 524400 31048
rect 520917 31043 520983 31046
rect 523200 31016 524400 31046
rect 114001 30426 114067 30429
rect 110860 30424 114067 30426
rect 110860 30368 114006 30424
rect 114062 30368 114067 30424
rect 110860 30366 114067 30368
rect 114001 30363 114067 30366
rect 520917 30290 520983 30293
rect 518758 30288 520983 30290
rect 518758 30232 520922 30288
rect 520978 30232 520983 30288
rect 518758 30230 520983 30232
rect 110689 29882 110755 29885
rect 111333 29882 111399 29885
rect 110689 29880 111399 29882
rect 110689 29824 110694 29880
rect 110750 29824 111338 29880
rect 111394 29824 111399 29880
rect 110689 29822 111399 29824
rect 110689 29819 110755 29822
rect 111333 29819 111399 29822
rect 117037 29882 117103 29885
rect 117037 29880 119140 29882
rect 117037 29824 117042 29880
rect 117098 29824 119140 29880
rect 117037 29822 119140 29824
rect 117037 29819 117103 29822
rect 518758 29716 518818 30230
rect 520917 30227 520983 30230
rect 110505 29610 110571 29613
rect 111057 29610 111123 29613
rect 110505 29608 111123 29610
rect 110505 29552 110510 29608
rect 110566 29552 111062 29608
rect 111118 29552 111123 29608
rect 110505 29550 111123 29552
rect 110505 29547 110571 29550
rect 111057 29547 111123 29550
rect 521101 29610 521167 29613
rect 523200 29610 524400 29640
rect 521101 29608 524400 29610
rect 521101 29552 521106 29608
rect 521162 29552 524400 29608
rect 521101 29550 524400 29552
rect 521101 29547 521167 29550
rect 523200 29520 524400 29550
rect 110321 29474 110387 29477
rect 110781 29474 110847 29477
rect 110321 29472 110847 29474
rect 110321 29416 110326 29472
rect 110382 29416 110786 29472
rect 110842 29416 110847 29472
rect 110321 29414 110847 29416
rect 110321 29411 110387 29414
rect 110781 29411 110847 29414
rect 110321 29338 110387 29341
rect 111149 29338 111215 29341
rect 110321 29336 111215 29338
rect 110321 29280 110326 29336
rect 110382 29280 111154 29336
rect 111210 29280 111215 29336
rect 110321 29278 111215 29280
rect 110321 29275 110387 29278
rect 111149 29275 111215 29278
rect 110321 29202 110387 29205
rect 111241 29202 111307 29205
rect 110321 29200 111307 29202
rect 110321 29144 110326 29200
rect 110382 29144 111246 29200
rect 111302 29144 111307 29200
rect 110321 29142 111307 29144
rect 110321 29139 110387 29142
rect 111241 29139 111307 29142
rect 521101 28386 521167 28389
rect 518788 28384 521167 28386
rect 518788 28328 521106 28384
rect 521162 28328 521167 28384
rect 518788 28326 521167 28328
rect 521101 28323 521167 28326
rect 523200 28114 524400 28144
rect 518850 28054 524400 28114
rect 117129 27978 117195 27981
rect 117129 27976 119140 27978
rect 117129 27920 117134 27976
rect 117190 27920 119140 27976
rect 117129 27918 119140 27920
rect 117129 27915 117195 27918
rect 518850 27570 518910 28054
rect 523200 28024 524400 28054
rect 518758 27510 518910 27570
rect 518758 26996 518818 27510
rect 523200 26482 524400 26512
rect 521610 26422 524400 26482
rect 521610 26210 521670 26422
rect 523200 26392 524400 26422
rect 518758 26150 521670 26210
rect 116393 26074 116459 26077
rect 116393 26072 119140 26074
rect 116393 26016 116398 26072
rect 116454 26016 119140 26072
rect 116393 26014 119140 26016
rect 116393 26011 116459 26014
rect 518758 25636 518818 26150
rect 523200 24986 524400 25016
rect 518850 24926 524400 24986
rect 518850 24850 518910 24926
rect 523200 24896 524400 24926
rect 518758 24790 518910 24850
rect 518758 24276 518818 24790
rect 117221 24170 117287 24173
rect 117221 24168 119140 24170
rect 117221 24112 117226 24168
rect 117282 24112 119140 24168
rect 117221 24110 119140 24112
rect 117221 24107 117287 24110
rect 523200 23490 524400 23520
rect 518758 23430 524400 23490
rect 518758 22916 518818 23430
rect 523200 23400 524400 23430
rect 116485 22266 116551 22269
rect 116485 22264 119140 22266
rect 116485 22208 116490 22264
rect 116546 22208 119140 22264
rect 116485 22206 119140 22208
rect 116485 22203 116551 22206
rect 521101 21994 521167 21997
rect 523200 21994 524400 22024
rect 521101 21992 524400 21994
rect 521101 21936 521106 21992
rect 521162 21936 524400 21992
rect 521101 21934 524400 21936
rect 521101 21931 521167 21934
rect 523200 21904 524400 21934
rect 518758 20906 518818 21556
rect 521101 20906 521167 20909
rect 518758 20904 521167 20906
rect 518758 20848 521106 20904
rect 521162 20848 521167 20904
rect 518758 20846 521167 20848
rect 521101 20843 521167 20846
rect 520733 20498 520799 20501
rect 523200 20498 524400 20528
rect 520733 20496 524400 20498
rect 520733 20440 520738 20496
rect 520794 20440 524400 20496
rect 520733 20438 524400 20440
rect 520733 20435 520799 20438
rect 523200 20408 524400 20438
rect 116301 20362 116367 20365
rect 116301 20360 119140 20362
rect 116301 20304 116306 20360
rect 116362 20304 119140 20360
rect 116301 20302 119140 20304
rect 116301 20299 116367 20302
rect 110321 20226 110387 20229
rect 110781 20226 110847 20229
rect 110321 20224 110847 20226
rect 110321 20168 110326 20224
rect 110382 20168 110786 20224
rect 110842 20168 110847 20224
rect 110321 20166 110847 20168
rect 110321 20163 110387 20166
rect 110781 20163 110847 20166
rect 110597 20090 110663 20093
rect 110781 20090 110847 20093
rect 110597 20088 110847 20090
rect 110597 20032 110602 20088
rect 110658 20032 110786 20088
rect 110842 20032 110847 20088
rect 110597 20030 110847 20032
rect 110597 20027 110663 20030
rect 110781 20027 110847 20030
rect 518758 19546 518818 20196
rect 520733 19546 520799 19549
rect 518758 19544 520799 19546
rect 518758 19488 520738 19544
rect 520794 19488 520799 19544
rect 518758 19486 520799 19488
rect 520733 19483 520799 19486
rect 113909 19002 113975 19005
rect 110860 19000 113975 19002
rect 110860 18944 113914 19000
rect 113970 18944 113975 19000
rect 110860 18942 113975 18944
rect 113909 18939 113975 18942
rect 520917 19002 520983 19005
rect 523200 19002 524400 19032
rect 520917 19000 524400 19002
rect 520917 18944 520922 19000
rect 520978 18944 524400 19000
rect 520917 18942 524400 18944
rect 520917 18939 520983 18942
rect 523200 18912 524400 18942
rect 116209 18458 116275 18461
rect 116209 18456 119140 18458
rect 116209 18400 116214 18456
rect 116270 18400 119140 18456
rect 116209 18398 119140 18400
rect 116209 18395 116275 18398
rect 518758 18186 518818 18836
rect 520917 18186 520983 18189
rect 518758 18184 520983 18186
rect 518758 18128 520922 18184
rect 520978 18128 520983 18184
rect 518758 18126 520983 18128
rect 520917 18123 520983 18126
rect 518758 16826 518818 17476
rect 523200 17370 524400 17400
rect 521150 17310 524400 17370
rect 521150 16826 521210 17310
rect 523200 17280 524400 17310
rect 518758 16766 521210 16826
rect 116025 16418 116091 16421
rect 116025 16416 119140 16418
rect 116025 16360 116030 16416
rect 116086 16360 119140 16416
rect 116025 16358 119140 16360
rect 116025 16355 116091 16358
rect 518758 15466 518818 16116
rect 523200 15874 524400 15904
rect 521104 15814 524400 15874
rect 521104 15466 521164 15814
rect 523200 15784 524400 15814
rect 518758 15406 521164 15466
rect 116117 14514 116183 14517
rect 116117 14512 119140 14514
rect 116117 14456 116122 14512
rect 116178 14456 119140 14512
rect 116117 14454 119140 14456
rect 116117 14451 116183 14454
rect 518758 14106 518818 14756
rect 523200 14378 524400 14408
rect 521104 14318 524400 14378
rect 521104 14106 521164 14318
rect 523200 14288 524400 14318
rect 518758 14046 521164 14106
rect 518758 12746 518818 13396
rect 523200 12882 524400 12912
rect 521104 12822 524400 12882
rect 521104 12746 521164 12822
rect 523200 12792 524400 12822
rect 518758 12686 521164 12746
rect 115933 12610 115999 12613
rect 115933 12608 119140 12610
rect 115933 12552 115938 12608
rect 115994 12552 119140 12608
rect 115933 12550 119140 12552
rect 115933 12547 115999 12550
rect 110321 12474 110387 12477
rect 110965 12474 111031 12477
rect 110321 12472 111031 12474
rect 110321 12416 110326 12472
rect 110382 12416 110970 12472
rect 111026 12416 111031 12472
rect 110321 12414 111031 12416
rect 110321 12411 110387 12414
rect 110965 12411 111031 12414
rect 110321 12202 110387 12205
rect 110597 12202 110663 12205
rect 110321 12200 110663 12202
rect 110321 12144 110326 12200
rect 110382 12144 110602 12200
rect 110658 12144 110663 12200
rect 110321 12142 110663 12144
rect 110321 12139 110387 12142
rect 110597 12139 110663 12142
rect 518758 11386 518818 12036
rect 523200 11386 524400 11416
rect 518758 11326 524400 11386
rect 523200 11296 524400 11326
rect 116526 10644 116532 10708
rect 116596 10706 116602 10708
rect 116596 10646 119140 10706
rect 116596 10644 116602 10646
rect 518758 10026 518818 10676
rect 518758 9966 518910 10026
rect 518850 9890 518910 9966
rect 523200 9890 524400 9920
rect 518850 9830 524400 9890
rect 523200 9800 524400 9830
rect 110505 9754 110571 9757
rect 110873 9754 110939 9757
rect 110505 9752 110939 9754
rect 110505 9696 110510 9752
rect 110566 9696 110878 9752
rect 110934 9696 110939 9752
rect 110505 9694 110939 9696
rect 110505 9691 110571 9694
rect 110873 9691 110939 9694
rect 521101 9346 521167 9349
rect 518788 9344 521167 9346
rect 518788 9288 521106 9344
rect 521162 9288 521167 9344
rect 518788 9286 521167 9288
rect 521101 9283 521167 9286
rect 110321 9074 110387 9077
rect 110597 9074 110663 9077
rect 110321 9072 110663 9074
rect 110321 9016 110326 9072
rect 110382 9016 110602 9072
rect 110658 9016 110663 9072
rect 110321 9014 110663 9016
rect 110321 9011 110387 9014
rect 110597 9011 110663 9014
rect 110321 8802 110387 8805
rect 110965 8802 111031 8805
rect 110321 8800 111031 8802
rect 110321 8744 110326 8800
rect 110382 8744 110970 8800
rect 111026 8744 111031 8800
rect 110321 8742 111031 8744
rect 110321 8739 110387 8742
rect 110965 8739 111031 8742
rect 117262 8740 117268 8804
rect 117332 8802 117338 8804
rect 117332 8742 119140 8802
rect 117332 8740 117338 8742
rect 110321 8530 110387 8533
rect 111057 8530 111123 8533
rect 110321 8528 111123 8530
rect 110321 8472 110326 8528
rect 110382 8472 111062 8528
rect 111118 8472 111123 8528
rect 110321 8470 111123 8472
rect 110321 8467 110387 8470
rect 111057 8467 111123 8470
rect 110321 8394 110387 8397
rect 111333 8394 111399 8397
rect 110321 8392 111399 8394
rect 110321 8336 110326 8392
rect 110382 8336 111338 8392
rect 111394 8336 111399 8392
rect 110321 8334 111399 8336
rect 110321 8331 110387 8334
rect 111333 8331 111399 8334
rect 521101 8258 521167 8261
rect 523200 8258 524400 8288
rect 521101 8256 524400 8258
rect 521101 8200 521106 8256
rect 521162 8200 524400 8256
rect 521101 8198 524400 8200
rect 521101 8195 521167 8198
rect 523200 8168 524400 8198
rect 520365 7986 520431 7989
rect 518788 7984 520431 7986
rect 518788 7928 520370 7984
rect 520426 7928 520431 7984
rect 518788 7926 520431 7928
rect 520365 7923 520431 7926
rect 110413 7850 110479 7853
rect 110965 7850 111031 7853
rect 110413 7848 111031 7850
rect 110413 7792 110418 7848
rect 110474 7792 110970 7848
rect 111026 7792 111031 7848
rect 110413 7790 111031 7792
rect 110413 7787 110479 7790
rect 110965 7787 111031 7790
rect 113817 7714 113883 7717
rect 110860 7712 113883 7714
rect 110860 7656 113822 7712
rect 113878 7656 113883 7712
rect 110860 7654 113883 7656
rect 113817 7651 113883 7654
rect 116158 6836 116164 6900
rect 116228 6898 116234 6900
rect 116228 6838 119140 6898
rect 116228 6836 116234 6838
rect 520365 6762 520431 6765
rect 523200 6762 524400 6792
rect 520365 6760 524400 6762
rect 520365 6704 520370 6760
rect 520426 6704 524400 6760
rect 520365 6702 524400 6704
rect 520365 6699 520431 6702
rect 523200 6672 524400 6702
rect 521101 6626 521167 6629
rect 518788 6624 521167 6626
rect 518788 6568 521106 6624
rect 521162 6568 521167 6624
rect 518788 6566 521167 6568
rect 521101 6563 521167 6566
rect 110873 5674 110939 5677
rect 110324 5672 110939 5674
rect 110324 5616 110878 5672
rect 110934 5616 110939 5672
rect 110324 5614 110939 5616
rect 110324 5553 110384 5614
rect 110873 5611 110939 5614
rect 110321 5548 110387 5553
rect 110321 5492 110326 5548
rect 110382 5492 110387 5548
rect 110321 5487 110387 5492
rect 520917 5266 520983 5269
rect 518788 5264 520983 5266
rect 518788 5208 520922 5264
rect 520978 5208 520983 5264
rect 518788 5206 520983 5208
rect 520917 5203 520983 5206
rect 521101 5266 521167 5269
rect 523200 5266 524400 5296
rect 521101 5264 524400 5266
rect 521101 5208 521106 5264
rect 521162 5208 524400 5264
rect 521101 5206 524400 5208
rect 521101 5203 521167 5206
rect 523200 5176 524400 5206
rect 110689 4178 110755 4181
rect 119110 4178 119170 4964
rect 110689 4176 119170 4178
rect 110689 4120 110694 4176
rect 110750 4120 119170 4176
rect 110689 4118 119170 4120
rect 110689 4115 110755 4118
rect 71730 3982 91754 4042
rect 71730 3906 71790 3982
rect 70350 3846 71790 3906
rect 73110 3846 84026 3906
rect 70350 3634 70410 3846
rect 67590 3574 70410 3634
rect 67590 3498 67650 3574
rect 73110 3498 73170 3846
rect 83966 3770 84026 3846
rect 55170 3438 59554 3498
rect 42750 3302 46950 3362
rect 35850 3030 37290 3090
rect 35850 2818 35910 3030
rect 33182 2758 35910 2818
rect 33041 2682 33107 2685
rect 33182 2682 33242 2758
rect 33041 2680 33242 2682
rect 33041 2624 33046 2680
rect 33102 2624 33242 2680
rect 33041 2622 33242 2624
rect 37230 2682 37290 3030
rect 42750 2685 42810 3302
rect 46890 3226 46950 3302
rect 55170 3226 55230 3438
rect 46890 3166 55230 3226
rect 46890 3030 56610 3090
rect 42057 2682 42123 2685
rect 37230 2680 42123 2682
rect 37230 2624 42062 2680
rect 42118 2624 42123 2680
rect 37230 2622 42123 2624
rect 33041 2619 33107 2622
rect 42057 2619 42123 2622
rect 42701 2680 42810 2685
rect 42701 2624 42706 2680
rect 42762 2624 42810 2680
rect 42701 2622 42810 2624
rect 44725 2682 44791 2685
rect 46890 2682 46950 3030
rect 44725 2680 46950 2682
rect 44725 2624 44730 2680
rect 44786 2624 46950 2680
rect 44725 2622 46950 2624
rect 56550 2682 56610 3030
rect 59494 2954 59554 3438
rect 66210 3438 67650 3498
rect 70350 3438 73170 3498
rect 78078 3710 81450 3770
rect 83966 3710 84394 3770
rect 66210 3362 66270 3438
rect 59126 2894 59554 2954
rect 62806 3302 66270 3362
rect 67590 3302 69030 3362
rect 59126 2685 59186 2894
rect 62806 2685 62866 3302
rect 67590 3226 67650 3302
rect 66210 3166 67650 3226
rect 68970 3226 69030 3302
rect 70350 3226 70410 3438
rect 78078 3362 78138 3710
rect 68970 3166 70410 3226
rect 72926 3302 78138 3362
rect 81390 3362 81450 3710
rect 84334 3498 84394 3710
rect 84334 3438 90420 3498
rect 81390 3302 89914 3362
rect 66210 2954 66270 3166
rect 64462 2894 66270 2954
rect 58985 2682 59051 2685
rect 56550 2680 59051 2682
rect 56550 2624 58990 2680
rect 59046 2624 59051 2680
rect 56550 2622 59051 2624
rect 59126 2680 59235 2685
rect 59126 2624 59174 2680
rect 59230 2624 59235 2680
rect 59126 2622 59235 2624
rect 42701 2619 42767 2622
rect 44725 2619 44791 2622
rect 58985 2619 59051 2622
rect 59169 2619 59235 2622
rect 62757 2680 62866 2685
rect 62757 2624 62762 2680
rect 62818 2624 62866 2680
rect 62757 2622 62866 2624
rect 63033 2682 63099 2685
rect 64462 2682 64522 2894
rect 72926 2818 72986 3302
rect 66210 2758 72986 2818
rect 73110 3166 89178 3226
rect 63033 2680 64522 2682
rect 63033 2624 63038 2680
rect 63094 2624 64522 2680
rect 63033 2622 64522 2624
rect 64597 2682 64663 2685
rect 66210 2682 66270 2758
rect 64597 2680 66270 2682
rect 64597 2624 64602 2680
rect 64658 2624 66270 2680
rect 64597 2622 66270 2624
rect 66989 2682 67055 2685
rect 73110 2682 73170 3166
rect 89118 3090 89178 3166
rect 89118 3030 89362 3090
rect 66989 2680 73170 2682
rect 66989 2624 66994 2680
rect 67050 2624 73170 2680
rect 66989 2622 73170 2624
rect 76557 2682 76623 2685
rect 89161 2682 89227 2685
rect 76557 2680 89227 2682
rect 76557 2624 76562 2680
rect 76618 2624 89166 2680
rect 89222 2624 89227 2680
rect 76557 2622 89227 2624
rect 89302 2682 89362 3030
rect 89854 2685 89914 3302
rect 90360 2685 90420 3438
rect 89713 2682 89779 2685
rect 89302 2680 89779 2682
rect 89302 2624 89718 2680
rect 89774 2624 89779 2680
rect 89302 2622 89779 2624
rect 89854 2680 89963 2685
rect 89854 2624 89902 2680
rect 89958 2624 89963 2680
rect 89854 2622 89963 2624
rect 62757 2619 62823 2622
rect 63033 2619 63099 2622
rect 64597 2619 64663 2622
rect 66989 2619 67055 2622
rect 76557 2619 76623 2622
rect 89161 2619 89227 2622
rect 89713 2619 89779 2622
rect 89897 2619 89963 2622
rect 90357 2680 90423 2685
rect 90357 2624 90362 2680
rect 90418 2624 90423 2680
rect 90357 2619 90423 2624
rect 91694 2682 91754 3982
rect 96570 3982 99390 4042
rect 96570 3634 96630 3982
rect 99330 3906 99390 3982
rect 110045 3906 110111 3909
rect 521009 3906 521075 3909
rect 99330 3904 110111 3906
rect 99330 3848 110050 3904
rect 110106 3848 110111 3904
rect 99330 3846 110111 3848
rect 518788 3904 521075 3906
rect 518788 3848 521014 3904
rect 521070 3848 521075 3904
rect 518788 3846 521075 3848
rect 110045 3843 110111 3846
rect 521009 3843 521075 3846
rect 116945 3770 117011 3773
rect 92752 3574 96630 3634
rect 96846 3768 117011 3770
rect 96846 3712 116950 3768
rect 117006 3712 117011 3768
rect 96846 3710 117011 3712
rect 92752 2685 92812 3574
rect 96846 3498 96906 3710
rect 116945 3707 117011 3710
rect 520917 3770 520983 3773
rect 523200 3770 524400 3800
rect 520917 3768 524400 3770
rect 520917 3712 520922 3768
rect 520978 3712 524400 3768
rect 520917 3710 524400 3712
rect 520917 3707 520983 3710
rect 523200 3680 524400 3710
rect 110965 3634 111031 3637
rect 99238 3632 111031 3634
rect 99238 3576 110970 3632
rect 111026 3576 111031 3632
rect 99238 3574 111031 3576
rect 99238 3498 99298 3574
rect 110965 3571 111031 3574
rect 117129 3498 117195 3501
rect 96570 3438 96906 3498
rect 97030 3438 99298 3498
rect 99606 3496 117195 3498
rect 99606 3440 117134 3496
rect 117190 3440 117195 3496
rect 99606 3438 117195 3440
rect 96570 3226 96630 3438
rect 95144 3166 96630 3226
rect 95144 2685 95204 3166
rect 97030 3090 97090 3438
rect 96570 3030 97090 3090
rect 96570 2818 96630 3030
rect 95374 2758 96630 2818
rect 95374 2685 95434 2758
rect 92473 2682 92539 2685
rect 91694 2680 92539 2682
rect 91694 2624 92478 2680
rect 92534 2624 92539 2680
rect 91694 2622 92539 2624
rect 92473 2619 92539 2622
rect 92749 2680 92815 2685
rect 92749 2624 92754 2680
rect 92810 2624 92815 2680
rect 92749 2619 92815 2624
rect 95141 2680 95207 2685
rect 95141 2624 95146 2680
rect 95202 2624 95207 2680
rect 95141 2619 95207 2624
rect 95325 2680 95434 2685
rect 95325 2624 95330 2680
rect 95386 2624 95434 2680
rect 95325 2622 95434 2624
rect 96429 2682 96495 2685
rect 99606 2682 99666 3438
rect 117129 3435 117195 3438
rect 116301 3362 116367 3365
rect 100526 3360 116367 3362
rect 100526 3304 116306 3360
rect 116362 3304 116367 3360
rect 100526 3302 116367 3304
rect 96429 2680 99666 2682
rect 96429 2624 96434 2680
rect 96490 2624 99666 2680
rect 96429 2622 99666 2624
rect 99925 2682 99991 2685
rect 100526 2682 100586 3302
rect 116301 3299 116367 3302
rect 109861 3226 109927 3229
rect 116761 3226 116827 3229
rect 100894 3224 109927 3226
rect 100894 3168 109866 3224
rect 109922 3168 109927 3224
rect 100894 3166 109927 3168
rect 100894 2685 100954 3166
rect 109861 3163 109927 3166
rect 112854 3224 116827 3226
rect 112854 3168 116766 3224
rect 116822 3168 116827 3224
rect 112854 3166 116827 3168
rect 112854 3090 112914 3166
rect 116761 3163 116827 3166
rect 101814 3030 112914 3090
rect 116301 3090 116367 3093
rect 116301 3088 119140 3090
rect 116301 3032 116306 3088
rect 116362 3032 119140 3088
rect 116301 3030 119140 3032
rect 101814 2685 101874 3030
rect 116301 3027 116367 3030
rect 109861 2954 109927 2957
rect 102550 2952 109927 2954
rect 102550 2896 109866 2952
rect 109922 2896 109927 2952
rect 102550 2894 109927 2896
rect 102550 2790 102610 2894
rect 109861 2891 109927 2894
rect 110321 2954 110387 2957
rect 110689 2954 110755 2957
rect 110321 2952 110755 2954
rect 110321 2896 110326 2952
rect 110382 2896 110694 2952
rect 110750 2896 110755 2952
rect 110321 2894 110755 2896
rect 110321 2891 110387 2894
rect 110689 2891 110755 2894
rect 111701 2818 111767 2821
rect 102182 2730 102610 2790
rect 106230 2816 111767 2818
rect 106230 2760 111706 2816
rect 111762 2760 111767 2816
rect 106230 2758 111767 2760
rect 99925 2680 100586 2682
rect 99925 2624 99930 2680
rect 99986 2624 100586 2680
rect 99925 2622 100586 2624
rect 100845 2680 100954 2685
rect 100845 2624 100850 2680
rect 100906 2624 100954 2680
rect 100845 2622 100954 2624
rect 101765 2680 101874 2685
rect 101765 2624 101770 2680
rect 101826 2624 101874 2680
rect 101765 2622 101874 2624
rect 101949 2682 102015 2685
rect 102182 2682 102242 2730
rect 101949 2680 102242 2682
rect 101949 2624 101954 2680
rect 102010 2624 102242 2680
rect 101949 2622 102242 2624
rect 102777 2682 102843 2685
rect 106230 2682 106290 2758
rect 111701 2755 111767 2758
rect 521101 2682 521167 2685
rect 102777 2680 106290 2682
rect 102777 2624 102782 2680
rect 102838 2624 106290 2680
rect 102777 2622 106290 2624
rect 518788 2680 521167 2682
rect 518788 2624 521106 2680
rect 521162 2624 521167 2680
rect 518788 2622 521167 2624
rect 95325 2619 95391 2622
rect 96429 2619 96495 2622
rect 99925 2619 99991 2622
rect 100845 2619 100911 2622
rect 101765 2619 101831 2622
rect 101949 2619 102015 2622
rect 102777 2619 102843 2622
rect 521101 2619 521167 2622
rect 29545 2546 29611 2549
rect 116209 2546 116275 2549
rect 29545 2544 116275 2546
rect 29545 2488 29550 2544
rect 29606 2488 116214 2544
rect 116270 2488 116275 2544
rect 29545 2486 116275 2488
rect 29545 2483 29611 2486
rect 116209 2483 116275 2486
rect 26049 2410 26115 2413
rect 116025 2410 116091 2413
rect 26049 2408 116091 2410
rect 26049 2352 26054 2408
rect 26110 2352 116030 2408
rect 116086 2352 116091 2408
rect 26049 2350 116091 2352
rect 26049 2347 26115 2350
rect 116025 2347 116091 2350
rect 22921 2274 22987 2277
rect 116117 2274 116183 2277
rect 22921 2272 116183 2274
rect 22921 2216 22926 2272
rect 22982 2216 116122 2272
rect 116178 2216 116183 2272
rect 22921 2214 116183 2216
rect 22921 2211 22987 2214
rect 116117 2211 116183 2214
rect 521009 2274 521075 2277
rect 523200 2274 524400 2304
rect 521009 2272 524400 2274
rect 521009 2216 521014 2272
rect 521070 2216 524400 2272
rect 521009 2214 524400 2216
rect 521009 2211 521075 2214
rect 523200 2184 524400 2214
rect 19609 2138 19675 2141
rect 115933 2138 115999 2141
rect 19609 2136 115999 2138
rect 19609 2080 19614 2136
rect 19670 2080 115938 2136
rect 115994 2080 115999 2136
rect 19609 2078 115999 2080
rect 19609 2075 19675 2078
rect 115933 2075 115999 2078
rect 16205 2002 16271 2005
rect 116526 2002 116532 2004
rect 16205 2000 116532 2002
rect 16205 1944 16210 2000
rect 16266 1944 116532 2000
rect 16205 1942 116532 1944
rect 16205 1939 16271 1942
rect 116526 1940 116532 1942
rect 116596 1940 116602 2004
rect 5993 1866 6059 1869
rect 110321 1866 110387 1869
rect 5993 1864 110387 1866
rect 5993 1808 5998 1864
rect 6054 1808 110326 1864
rect 110382 1808 110387 1864
rect 5993 1806 110387 1808
rect 5993 1803 6059 1806
rect 110321 1803 110387 1806
rect 12617 1730 12683 1733
rect 117262 1730 117268 1732
rect 12617 1728 117268 1730
rect 12617 1672 12622 1728
rect 12678 1672 117268 1728
rect 12617 1670 117268 1672
rect 12617 1667 12683 1670
rect 117262 1668 117268 1670
rect 117332 1668 117338 1732
rect 229277 1730 229343 1733
rect 293585 1730 293651 1733
rect 229277 1728 293651 1730
rect 229277 1672 229282 1728
rect 229338 1672 293590 1728
rect 293646 1672 293651 1728
rect 229277 1670 293651 1672
rect 229277 1667 229343 1670
rect 293585 1667 293651 1670
rect 9305 1594 9371 1597
rect 116158 1594 116164 1596
rect 9305 1592 116164 1594
rect 9305 1536 9310 1592
rect 9366 1536 116164 1592
rect 9305 1534 116164 1536
rect 9305 1531 9371 1534
rect 116158 1532 116164 1534
rect 116228 1532 116234 1596
rect 163773 1594 163839 1597
rect 243629 1594 243695 1597
rect 163773 1592 243695 1594
rect 163773 1536 163778 1592
rect 163834 1536 243634 1592
rect 243690 1536 243695 1592
rect 163773 1534 243695 1536
rect 163773 1531 163839 1534
rect 243629 1531 243695 1534
rect 55949 1458 56015 1461
rect 294781 1458 294847 1461
rect 55949 1456 294847 1458
rect 55949 1400 55954 1456
rect 56010 1400 294786 1456
rect 294842 1400 294847 1456
rect 55949 1398 294847 1400
rect 55949 1395 56015 1398
rect 294781 1395 294847 1398
rect 360285 1458 360351 1461
rect 393589 1458 393655 1461
rect 360285 1456 393655 1458
rect 360285 1400 360290 1456
rect 360346 1400 393594 1456
rect 393650 1400 393655 1456
rect 360285 1398 393655 1400
rect 360285 1395 360351 1398
rect 393589 1395 393655 1398
rect 89897 1322 89963 1325
rect 96429 1322 96495 1325
rect 89897 1320 96495 1322
rect 89897 1264 89902 1320
rect 89958 1264 96434 1320
rect 96490 1264 96495 1320
rect 89897 1262 96495 1264
rect 89897 1259 89963 1262
rect 96429 1259 96495 1262
rect 98269 1322 98335 1325
rect 101949 1322 102015 1325
rect 98269 1320 102015 1322
rect 98269 1264 98274 1320
rect 98330 1264 101954 1320
rect 102010 1264 102015 1320
rect 98269 1262 102015 1264
rect 98269 1259 98335 1262
rect 101949 1259 102015 1262
rect 89161 1186 89227 1189
rect 95141 1186 95207 1189
rect 89161 1184 95207 1186
rect 89161 1128 89166 1184
rect 89222 1128 95146 1184
rect 95202 1128 95207 1184
rect 89161 1126 95207 1128
rect 89161 1123 89227 1126
rect 95141 1123 95207 1126
rect 521101 778 521167 781
rect 523200 778 524400 808
rect 521101 776 524400 778
rect 521101 720 521106 776
rect 521162 720 524400 776
rect 521101 718 524400 720
rect 521101 715 521167 718
rect 523200 688 524400 718
<< via3 >>
rect 116532 10644 116596 10708
rect 117268 8740 117332 8804
rect 116164 6836 116228 6900
rect 116532 1940 116596 2004
rect 117268 1668 117332 1732
rect 116164 1532 116228 1596
<< metal4 >>
rect 1664 144454 1984 144496
rect 1664 144218 1706 144454
rect 1942 144218 1984 144454
rect 1664 144134 1984 144218
rect 1664 143898 1706 144134
rect 1942 143898 1984 144134
rect 1664 143856 1984 143898
rect 109956 144454 110276 144496
rect 109956 144218 109998 144454
rect 110234 144218 110276 144454
rect 109956 144134 110276 144218
rect 109956 143898 109998 144134
rect 110234 143898 110276 144134
rect 109956 143856 110276 143898
rect 119664 144454 119984 144496
rect 119664 144218 119706 144454
rect 119942 144218 119984 144454
rect 119664 144134 119984 144218
rect 119664 143898 119706 144134
rect 119942 143898 119984 144134
rect 119664 143856 119984 143898
rect 517940 144454 518260 144496
rect 517940 144218 517982 144454
rect 518218 144218 518260 144454
rect 517940 144134 518260 144218
rect 517940 143898 517982 144134
rect 518218 143898 518260 144134
rect 517940 143856 518260 143898
rect 1096 131454 1332 131496
rect 1096 131134 1332 131218
rect 1096 130856 1332 130898
rect 110616 131454 110936 131496
rect 110616 131218 110658 131454
rect 110894 131218 110936 131454
rect 110616 131134 110936 131218
rect 110616 130898 110658 131134
rect 110894 130898 110936 131134
rect 110616 130856 110936 130898
rect 119004 131454 119324 131496
rect 119004 131218 119046 131454
rect 119282 131218 119324 131454
rect 119004 131134 119324 131218
rect 119004 130898 119046 131134
rect 119282 130898 119324 131134
rect 119004 130856 119324 130898
rect 518600 131454 518920 131496
rect 518600 131218 518642 131454
rect 518878 131218 518920 131454
rect 518600 131134 518920 131218
rect 518600 130898 518642 131134
rect 518878 130898 518920 131134
rect 518600 130856 518920 130898
rect 1664 118454 1984 118496
rect 1664 118218 1706 118454
rect 1942 118218 1984 118454
rect 1664 118134 1984 118218
rect 1664 117898 1706 118134
rect 1942 117898 1984 118134
rect 1664 117856 1984 117898
rect 109956 118454 110276 118496
rect 109956 118218 109998 118454
rect 110234 118218 110276 118454
rect 109956 118134 110276 118218
rect 109956 117898 109998 118134
rect 110234 117898 110276 118134
rect 109956 117856 110276 117898
rect 119664 118454 119984 118496
rect 119664 118218 119706 118454
rect 119942 118218 119984 118454
rect 119664 118134 119984 118218
rect 119664 117898 119706 118134
rect 119942 117898 119984 118134
rect 119664 117856 119984 117898
rect 517940 118454 518260 118496
rect 517940 118218 517982 118454
rect 518218 118218 518260 118454
rect 517940 118134 518260 118218
rect 517940 117898 517982 118134
rect 518218 117898 518260 118134
rect 517940 117856 518260 117898
rect 1096 105454 1332 105496
rect 1096 105134 1332 105218
rect 1096 104856 1332 104898
rect 110616 105454 110936 105496
rect 110616 105218 110658 105454
rect 110894 105218 110936 105454
rect 110616 105134 110936 105218
rect 110616 104898 110658 105134
rect 110894 104898 110936 105134
rect 110616 104856 110936 104898
rect 119004 105454 119324 105496
rect 119004 105218 119046 105454
rect 119282 105218 119324 105454
rect 119004 105134 119324 105218
rect 119004 104898 119046 105134
rect 119282 104898 119324 105134
rect 119004 104856 119324 104898
rect 518600 105454 518920 105496
rect 518600 105218 518642 105454
rect 518878 105218 518920 105454
rect 518600 105134 518920 105218
rect 518600 104898 518642 105134
rect 518878 104898 518920 105134
rect 518600 104856 518920 104898
rect 1664 92454 1984 92496
rect 1664 92218 1706 92454
rect 1942 92218 1984 92454
rect 1664 92134 1984 92218
rect 1664 91898 1706 92134
rect 1942 91898 1984 92134
rect 1664 91856 1984 91898
rect 109956 92454 110276 92496
rect 109956 92218 109998 92454
rect 110234 92218 110276 92454
rect 109956 92134 110276 92218
rect 109956 91898 109998 92134
rect 110234 91898 110276 92134
rect 109956 91856 110276 91898
rect 119664 92454 119984 92496
rect 119664 92218 119706 92454
rect 119942 92218 119984 92454
rect 119664 92134 119984 92218
rect 119664 91898 119706 92134
rect 119942 91898 119984 92134
rect 119664 91856 119984 91898
rect 517940 92454 518260 92496
rect 517940 92218 517982 92454
rect 518218 92218 518260 92454
rect 517940 92134 518260 92218
rect 517940 91898 517982 92134
rect 518218 91898 518260 92134
rect 517940 91856 518260 91898
rect 1096 79454 1332 79496
rect 1096 79134 1332 79218
rect 1096 78856 1332 78898
rect 110616 79454 110936 79496
rect 110616 79218 110658 79454
rect 110894 79218 110936 79454
rect 110616 79134 110936 79218
rect 110616 78898 110658 79134
rect 110894 78898 110936 79134
rect 110616 78856 110936 78898
rect 119004 79454 119324 79496
rect 119004 79218 119046 79454
rect 119282 79218 119324 79454
rect 119004 79134 119324 79218
rect 119004 78898 119046 79134
rect 119282 78898 119324 79134
rect 119004 78856 119324 78898
rect 518600 79454 518920 79496
rect 518600 79218 518642 79454
rect 518878 79218 518920 79454
rect 518600 79134 518920 79218
rect 518600 78898 518642 79134
rect 518878 78898 518920 79134
rect 518600 78856 518920 78898
rect 1664 66454 1984 66496
rect 1664 66218 1706 66454
rect 1942 66218 1984 66454
rect 1664 66134 1984 66218
rect 1664 65898 1706 66134
rect 1942 65898 1984 66134
rect 1664 65856 1984 65898
rect 109956 66454 110276 66496
rect 109956 66218 109998 66454
rect 110234 66218 110276 66454
rect 109956 66134 110276 66218
rect 109956 65898 109998 66134
rect 110234 65898 110276 66134
rect 109956 65856 110276 65898
rect 119664 66454 119984 66496
rect 119664 66218 119706 66454
rect 119942 66218 119984 66454
rect 119664 66134 119984 66218
rect 119664 65898 119706 66134
rect 119942 65898 119984 66134
rect 119664 65856 119984 65898
rect 517940 66454 518260 66496
rect 517940 66218 517982 66454
rect 518218 66218 518260 66454
rect 517940 66134 518260 66218
rect 517940 65898 517982 66134
rect 518218 65898 518260 66134
rect 517940 65856 518260 65898
rect 1096 53454 1332 53496
rect 1096 53134 1332 53218
rect 1096 52856 1332 52898
rect 110616 53454 110936 53496
rect 110616 53218 110658 53454
rect 110894 53218 110936 53454
rect 110616 53134 110936 53218
rect 110616 52898 110658 53134
rect 110894 52898 110936 53134
rect 110616 52856 110936 52898
rect 119004 53454 119324 53496
rect 119004 53218 119046 53454
rect 119282 53218 119324 53454
rect 119004 53134 119324 53218
rect 119004 52898 119046 53134
rect 119282 52898 119324 53134
rect 119004 52856 119324 52898
rect 518600 53454 518920 53496
rect 518600 53218 518642 53454
rect 518878 53218 518920 53454
rect 518600 53134 518920 53218
rect 518600 52898 518642 53134
rect 518878 52898 518920 53134
rect 518600 52856 518920 52898
rect 1664 40454 1984 40496
rect 1664 40218 1706 40454
rect 1942 40218 1984 40454
rect 1664 40134 1984 40218
rect 1664 39898 1706 40134
rect 1942 39898 1984 40134
rect 1664 39856 1984 39898
rect 109956 40454 110276 40496
rect 109956 40218 109998 40454
rect 110234 40218 110276 40454
rect 109956 40134 110276 40218
rect 109956 39898 109998 40134
rect 110234 39898 110276 40134
rect 109956 39856 110276 39898
rect 119664 40454 119984 40496
rect 119664 40218 119706 40454
rect 119942 40218 119984 40454
rect 119664 40134 119984 40218
rect 119664 39898 119706 40134
rect 119942 39898 119984 40134
rect 119664 39856 119984 39898
rect 517940 40454 518260 40496
rect 517940 40218 517982 40454
rect 518218 40218 518260 40454
rect 517940 40134 518260 40218
rect 517940 39898 517982 40134
rect 518218 39898 518260 40134
rect 517940 39856 518260 39898
rect 1096 27454 1332 27496
rect 1096 27134 1332 27218
rect 1096 26856 1332 26898
rect 110616 27454 110936 27496
rect 110616 27218 110658 27454
rect 110894 27218 110936 27454
rect 110616 27134 110936 27218
rect 110616 26898 110658 27134
rect 110894 26898 110936 27134
rect 110616 26856 110936 26898
rect 119004 27454 119324 27496
rect 119004 27218 119046 27454
rect 119282 27218 119324 27454
rect 119004 27134 119324 27218
rect 119004 26898 119046 27134
rect 119282 26898 119324 27134
rect 119004 26856 119324 26898
rect 518600 27454 518920 27496
rect 518600 27218 518642 27454
rect 518878 27218 518920 27454
rect 518600 27134 518920 27218
rect 518600 26898 518642 27134
rect 518878 26898 518920 27134
rect 518600 26856 518920 26898
rect 1664 14454 1984 14496
rect 1664 14218 1706 14454
rect 1942 14218 1984 14454
rect 1664 14134 1984 14218
rect 1664 13898 1706 14134
rect 1942 13898 1984 14134
rect 1664 13856 1984 13898
rect 109956 14454 110276 14496
rect 109956 14218 109998 14454
rect 110234 14218 110276 14454
rect 109956 14134 110276 14218
rect 109956 13898 109998 14134
rect 110234 13898 110276 14134
rect 109956 13856 110276 13898
rect 119664 14454 119984 14496
rect 119664 14218 119706 14454
rect 119942 14218 119984 14454
rect 119664 14134 119984 14218
rect 119664 13898 119706 14134
rect 119942 13898 119984 14134
rect 119664 13856 119984 13898
rect 517940 14454 518260 14496
rect 517940 14218 517982 14454
rect 518218 14218 518260 14454
rect 517940 14134 518260 14218
rect 517940 13898 517982 14134
rect 518218 13898 518260 14134
rect 517940 13856 518260 13898
rect 116531 10708 116597 10709
rect 116531 10644 116532 10708
rect 116596 10644 116597 10708
rect 116531 10643 116597 10644
rect 116163 6900 116229 6901
rect 116163 6836 116164 6900
rect 116228 6836 116229 6900
rect 116163 6835 116229 6836
rect 116166 1597 116226 6835
rect 116534 2005 116594 10643
rect 117267 8804 117333 8805
rect 117267 8740 117268 8804
rect 117332 8740 117333 8804
rect 117267 8739 117333 8740
rect 116531 2004 116597 2005
rect 116531 1940 116532 2004
rect 116596 1940 116597 2004
rect 116531 1939 116597 1940
rect 117270 1733 117330 8739
rect 117267 1732 117333 1733
rect 117267 1668 117268 1732
rect 117332 1668 117333 1732
rect 117267 1667 117333 1668
rect 116163 1596 116229 1597
rect 116163 1532 116164 1596
rect 116228 1532 116229 1596
rect 116163 1531 116229 1532
<< via4 >>
rect 1706 144218 1942 144454
rect 1706 143898 1942 144134
rect 109998 144218 110234 144454
rect 109998 143898 110234 144134
rect 119706 144218 119942 144454
rect 119706 143898 119942 144134
rect 517982 144218 518218 144454
rect 517982 143898 518218 144134
rect 1096 131218 1332 131454
rect 1096 130898 1332 131134
rect 110658 131218 110894 131454
rect 110658 130898 110894 131134
rect 119046 131218 119282 131454
rect 119046 130898 119282 131134
rect 518642 131218 518878 131454
rect 518642 130898 518878 131134
rect 1706 118218 1942 118454
rect 1706 117898 1942 118134
rect 109998 118218 110234 118454
rect 109998 117898 110234 118134
rect 119706 118218 119942 118454
rect 119706 117898 119942 118134
rect 517982 118218 518218 118454
rect 517982 117898 518218 118134
rect 1096 105218 1332 105454
rect 1096 104898 1332 105134
rect 110658 105218 110894 105454
rect 110658 104898 110894 105134
rect 119046 105218 119282 105454
rect 119046 104898 119282 105134
rect 518642 105218 518878 105454
rect 518642 104898 518878 105134
rect 1706 92218 1942 92454
rect 1706 91898 1942 92134
rect 109998 92218 110234 92454
rect 109998 91898 110234 92134
rect 119706 92218 119942 92454
rect 119706 91898 119942 92134
rect 517982 92218 518218 92454
rect 517982 91898 518218 92134
rect 1096 79218 1332 79454
rect 1096 78898 1332 79134
rect 110658 79218 110894 79454
rect 110658 78898 110894 79134
rect 119046 79218 119282 79454
rect 119046 78898 119282 79134
rect 518642 79218 518878 79454
rect 518642 78898 518878 79134
rect 1706 66218 1942 66454
rect 1706 65898 1942 66134
rect 109998 66218 110234 66454
rect 109998 65898 110234 66134
rect 119706 66218 119942 66454
rect 119706 65898 119942 66134
rect 517982 66218 518218 66454
rect 517982 65898 518218 66134
rect 1096 53218 1332 53454
rect 1096 52898 1332 53134
rect 110658 53218 110894 53454
rect 110658 52898 110894 53134
rect 119046 53218 119282 53454
rect 119046 52898 119282 53134
rect 518642 53218 518878 53454
rect 518642 52898 518878 53134
rect 1706 40218 1942 40454
rect 1706 39898 1942 40134
rect 109998 40218 110234 40454
rect 109998 39898 110234 40134
rect 119706 40218 119942 40454
rect 119706 39898 119942 40134
rect 517982 40218 518218 40454
rect 517982 39898 518218 40134
rect 1096 27218 1332 27454
rect 1096 26898 1332 27134
rect 110658 27218 110894 27454
rect 110658 26898 110894 27134
rect 119046 27218 119282 27454
rect 119046 26898 119282 27134
rect 518642 27218 518878 27454
rect 518642 26898 518878 27134
rect 1706 14218 1942 14454
rect 1706 13898 1942 14134
rect 109998 14218 110234 14454
rect 109998 13898 110234 14134
rect 119706 14218 119942 14454
rect 119706 13898 119942 14134
rect 517982 14218 518218 14454
rect 517982 13898 518218 14134
<< metal5 >>
rect 1104 156856 522836 157496
rect 1104 144454 2200 144496
rect 1104 144218 1706 144454
rect 1942 144218 2200 144454
rect 1104 144134 2200 144218
rect 1104 143898 1706 144134
rect 1942 143898 2200 144134
rect 1104 143856 2200 143898
rect 109800 144454 120200 144496
rect 109800 144218 109998 144454
rect 110234 144218 119706 144454
rect 119942 144218 120200 144454
rect 109800 144134 120200 144218
rect 109800 143898 109998 144134
rect 110234 143898 119706 144134
rect 119942 143898 120200 144134
rect 109800 143856 120200 143898
rect 517800 144454 522836 144496
rect 517800 144218 517982 144454
rect 518218 144218 522836 144454
rect 517800 144134 522836 144218
rect 517800 143898 517982 144134
rect 518218 143898 522836 144134
rect 517800 143856 522836 143898
rect 1072 131454 2200 131496
rect 1072 131218 1096 131454
rect 1332 131218 2200 131454
rect 1072 131134 2200 131218
rect 1072 130898 1096 131134
rect 1332 130898 2200 131134
rect 1072 130856 2200 130898
rect 109800 131454 120200 131496
rect 109800 131218 110658 131454
rect 110894 131218 119046 131454
rect 119282 131218 120200 131454
rect 109800 131134 120200 131218
rect 109800 130898 110658 131134
rect 110894 130898 119046 131134
rect 119282 130898 120200 131134
rect 109800 130856 120200 130898
rect 517800 131454 522836 131496
rect 517800 131218 518642 131454
rect 518878 131218 522836 131454
rect 517800 131134 522836 131218
rect 517800 130898 518642 131134
rect 518878 130898 522836 131134
rect 517800 130856 522836 130898
rect 1104 118454 2200 118496
rect 1104 118218 1706 118454
rect 1942 118218 2200 118454
rect 1104 118134 2200 118218
rect 1104 117898 1706 118134
rect 1942 117898 2200 118134
rect 1104 117856 2200 117898
rect 109800 118454 120200 118496
rect 109800 118218 109998 118454
rect 110234 118218 119706 118454
rect 119942 118218 120200 118454
rect 109800 118134 120200 118218
rect 109800 117898 109998 118134
rect 110234 117898 119706 118134
rect 119942 117898 120200 118134
rect 109800 117856 120200 117898
rect 517800 118454 522836 118496
rect 517800 118218 517982 118454
rect 518218 118218 522836 118454
rect 517800 118134 522836 118218
rect 517800 117898 517982 118134
rect 518218 117898 522836 118134
rect 517800 117856 522836 117898
rect 1072 105454 2200 105496
rect 1072 105218 1096 105454
rect 1332 105218 2200 105454
rect 1072 105134 2200 105218
rect 1072 104898 1096 105134
rect 1332 104898 2200 105134
rect 1072 104856 2200 104898
rect 109800 105454 120200 105496
rect 109800 105218 110658 105454
rect 110894 105218 119046 105454
rect 119282 105218 120200 105454
rect 109800 105134 120200 105218
rect 109800 104898 110658 105134
rect 110894 104898 119046 105134
rect 119282 104898 120200 105134
rect 109800 104856 120200 104898
rect 517800 105454 522836 105496
rect 517800 105218 518642 105454
rect 518878 105218 522836 105454
rect 517800 105134 522836 105218
rect 517800 104898 518642 105134
rect 518878 104898 522836 105134
rect 517800 104856 522836 104898
rect 1104 92454 2200 92496
rect 1104 92218 1706 92454
rect 1942 92218 2200 92454
rect 1104 92134 2200 92218
rect 1104 91898 1706 92134
rect 1942 91898 2200 92134
rect 1104 91856 2200 91898
rect 109800 92454 120200 92496
rect 109800 92218 109998 92454
rect 110234 92218 119706 92454
rect 119942 92218 120200 92454
rect 109800 92134 120200 92218
rect 109800 91898 109998 92134
rect 110234 91898 119706 92134
rect 119942 91898 120200 92134
rect 109800 91856 120200 91898
rect 517800 92454 522836 92496
rect 517800 92218 517982 92454
rect 518218 92218 522836 92454
rect 517800 92134 522836 92218
rect 517800 91898 517982 92134
rect 518218 91898 522836 92134
rect 517800 91856 522836 91898
rect 1072 79454 2200 79496
rect 1072 79218 1096 79454
rect 1332 79218 2200 79454
rect 1072 79134 2200 79218
rect 1072 78898 1096 79134
rect 1332 78898 2200 79134
rect 1072 78856 2200 78898
rect 109800 79454 120200 79496
rect 109800 79218 110658 79454
rect 110894 79218 119046 79454
rect 119282 79218 120200 79454
rect 109800 79134 120200 79218
rect 109800 78898 110658 79134
rect 110894 78898 119046 79134
rect 119282 78898 120200 79134
rect 109800 78856 120200 78898
rect 517800 79454 522836 79496
rect 517800 79218 518642 79454
rect 518878 79218 522836 79454
rect 517800 79134 522836 79218
rect 517800 78898 518642 79134
rect 518878 78898 522836 79134
rect 517800 78856 522836 78898
rect 1104 66454 2200 66496
rect 1104 66218 1706 66454
rect 1942 66218 2200 66454
rect 1104 66134 2200 66218
rect 1104 65898 1706 66134
rect 1942 65898 2200 66134
rect 1104 65856 2200 65898
rect 109800 66454 120200 66496
rect 109800 66218 109998 66454
rect 110234 66218 119706 66454
rect 119942 66218 120200 66454
rect 109800 66134 120200 66218
rect 109800 65898 109998 66134
rect 110234 65898 119706 66134
rect 119942 65898 120200 66134
rect 109800 65856 120200 65898
rect 517800 66454 522836 66496
rect 517800 66218 517982 66454
rect 518218 66218 522836 66454
rect 517800 66134 522836 66218
rect 517800 65898 517982 66134
rect 518218 65898 522836 66134
rect 517800 65856 522836 65898
rect 1072 53454 2200 53496
rect 1072 53218 1096 53454
rect 1332 53218 2200 53454
rect 1072 53134 2200 53218
rect 1072 52898 1096 53134
rect 1332 52898 2200 53134
rect 1072 52856 2200 52898
rect 109800 53454 120200 53496
rect 109800 53218 110658 53454
rect 110894 53218 119046 53454
rect 119282 53218 120200 53454
rect 109800 53134 120200 53218
rect 109800 52898 110658 53134
rect 110894 52898 119046 53134
rect 119282 52898 120200 53134
rect 109800 52856 120200 52898
rect 517800 53454 522836 53496
rect 517800 53218 518642 53454
rect 518878 53218 522836 53454
rect 517800 53134 522836 53218
rect 517800 52898 518642 53134
rect 518878 52898 522836 53134
rect 517800 52856 522836 52898
rect 1104 40454 2200 40496
rect 1104 40218 1706 40454
rect 1942 40218 2200 40454
rect 1104 40134 2200 40218
rect 1104 39898 1706 40134
rect 1942 39898 2200 40134
rect 1104 39856 2200 39898
rect 109800 40454 120200 40496
rect 109800 40218 109998 40454
rect 110234 40218 119706 40454
rect 119942 40218 120200 40454
rect 109800 40134 120200 40218
rect 109800 39898 109998 40134
rect 110234 39898 119706 40134
rect 119942 39898 120200 40134
rect 109800 39856 120200 39898
rect 517800 40454 522836 40496
rect 517800 40218 517982 40454
rect 518218 40218 522836 40454
rect 517800 40134 522836 40218
rect 517800 39898 517982 40134
rect 518218 39898 522836 40134
rect 517800 39856 522836 39898
rect 1072 27454 2200 27496
rect 1072 27218 1096 27454
rect 1332 27218 2200 27454
rect 1072 27134 2200 27218
rect 1072 26898 1096 27134
rect 1332 26898 2200 27134
rect 1072 26856 2200 26898
rect 109800 27454 120200 27496
rect 109800 27218 110658 27454
rect 110894 27218 119046 27454
rect 119282 27218 120200 27454
rect 109800 27134 120200 27218
rect 109800 26898 110658 27134
rect 110894 26898 119046 27134
rect 119282 26898 120200 27134
rect 109800 26856 120200 26898
rect 517800 27454 522836 27496
rect 517800 27218 518642 27454
rect 518878 27218 522836 27454
rect 517800 27134 522836 27218
rect 517800 26898 518642 27134
rect 518878 26898 522836 27134
rect 517800 26856 522836 26898
rect 1104 14454 2200 14496
rect 1104 14218 1706 14454
rect 1942 14218 2200 14454
rect 1104 14134 2200 14218
rect 1104 13898 1706 14134
rect 1942 13898 2200 14134
rect 1104 13856 2200 13898
rect 109800 14454 120200 14496
rect 109800 14218 109998 14454
rect 110234 14218 119706 14454
rect 119942 14218 120200 14454
rect 109800 14134 120200 14218
rect 109800 13898 109998 14134
rect 110234 13898 119706 14134
rect 119942 13898 120200 14134
rect 109800 13856 120200 13898
rect 517800 14454 522836 14496
rect 517800 14218 517982 14454
rect 518218 14218 522836 14454
rect 517800 14134 522836 14218
rect 517800 13898 517982 14134
rect 518218 13898 522836 14134
rect 517800 13856 522836 13898
use mgmt_core  core
timestamp 1638229739
transform 1 0 119000 0 1 2000
box 0 0 400000 148000
use DFFRAM  DFFRAM
timestamp 1638229739
transform 1 0 1000 0 1 2000
box 4 0 110000 148000
<< labels >>
rlabel metal5 s 1104 26856 2200 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 26856 120200 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 26856 522836 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 52856 2200 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 52856 120200 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 52856 522836 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 78856 2200 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 78856 120200 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 78856 522836 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 104856 2200 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 104856 120200 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 104856 522836 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 130856 2200 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 130856 120200 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 130856 522836 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 156856 522836 157496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 13856 2200 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 13856 120200 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 13856 522836 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 39856 2200 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 39856 120200 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 39856 522836 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 65856 2200 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 65856 120200 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 65856 522836 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 91856 2200 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 91856 120200 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 91856 522836 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 117856 2200 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 117856 120200 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 117856 522836 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 143856 2200 144496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 143856 120200 144496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 143856 522836 144496 6 VPWR
port 1 nsew power input
rlabel metal2 s 294786 -400 294842 800 6 core_clk
port 2 nsew signal input
rlabel metal2 s 98274 -400 98330 800 6 core_rstn
port 3 nsew signal input
rlabel metal3 s 523200 64472 524400 64592 6 debug_in
port 4 nsew signal input
rlabel metal3 s 523200 65968 524400 66088 6 debug_mode
port 5 nsew signal tristate
rlabel metal3 s 523200 67464 524400 67584 6 debug_oeb
port 6 nsew signal tristate
rlabel metal3 s 523200 68960 524400 69080 6 debug_out
port 7 nsew signal tristate
rlabel metal3 s 523200 144848 524400 144968 6 flash_clk
port 8 nsew signal tristate
rlabel metal3 s 523200 143352 524400 143472 6 flash_csb
port 9 nsew signal tristate
rlabel metal3 s 523200 146480 524400 146600 6 flash_io0_di
port 10 nsew signal input
rlabel metal3 s 523200 147976 524400 148096 6 flash_io0_do
port 11 nsew signal tristate
rlabel metal3 s 523200 149472 524400 149592 6 flash_io0_oeb
port 12 nsew signal tristate
rlabel metal3 s 523200 150968 524400 151088 6 flash_io1_di
port 13 nsew signal input
rlabel metal3 s 523200 152464 524400 152584 6 flash_io1_do
port 14 nsew signal tristate
rlabel metal3 s 523200 153960 524400 154080 6 flash_io1_oeb
port 15 nsew signal tristate
rlabel metal3 s 523200 155592 524400 155712 6 flash_io2_di
port 16 nsew signal input
rlabel metal3 s 523200 157088 524400 157208 6 flash_io2_do
port 17 nsew signal tristate
rlabel metal3 s 523200 158584 524400 158704 6 flash_io2_oeb
port 18 nsew signal tristate
rlabel metal3 s 523200 160080 524400 160200 6 flash_io3_di
port 19 nsew signal input
rlabel metal3 s 523200 161576 524400 161696 6 flash_io3_do
port 20 nsew signal tristate
rlabel metal3 s 523200 163072 524400 163192 6 flash_io3_oeb
port 21 nsew signal tristate
rlabel metal2 s 32770 -400 32826 800 6 gpio_in_pad
port 22 nsew signal input
rlabel metal2 s 163778 -400 163834 800 6 gpio_inenb_pad
port 23 nsew signal tristate
rlabel metal2 s 229282 -400 229338 800 6 gpio_mode0_pad
port 24 nsew signal tristate
rlabel metal2 s 360290 -400 360346 800 6 gpio_mode1_pad
port 25 nsew signal tristate
rlabel metal2 s 425794 -400 425850 800 6 gpio_out_pad
port 26 nsew signal tristate
rlabel metal2 s 491298 -400 491354 800 6 gpio_outenb_pad
port 27 nsew signal tristate
rlabel metal3 s 523200 91808 524400 91928 6 hk_ack_i
port 28 nsew signal input
rlabel metal3 s 523200 94800 524400 94920 6 hk_dat_i[0]
port 29 nsew signal input
rlabel metal3 s 523200 110032 524400 110152 6 hk_dat_i[10]
port 30 nsew signal input
rlabel metal3 s 523200 111528 524400 111648 6 hk_dat_i[11]
port 31 nsew signal input
rlabel metal3 s 523200 113024 524400 113144 6 hk_dat_i[12]
port 32 nsew signal input
rlabel metal3 s 523200 114520 524400 114640 6 hk_dat_i[13]
port 33 nsew signal input
rlabel metal3 s 523200 116016 524400 116136 6 hk_dat_i[14]
port 34 nsew signal input
rlabel metal3 s 523200 117512 524400 117632 6 hk_dat_i[15]
port 35 nsew signal input
rlabel metal3 s 523200 119144 524400 119264 6 hk_dat_i[16]
port 36 nsew signal input
rlabel metal3 s 523200 120640 524400 120760 6 hk_dat_i[17]
port 37 nsew signal input
rlabel metal3 s 523200 122136 524400 122256 6 hk_dat_i[18]
port 38 nsew signal input
rlabel metal3 s 523200 123632 524400 123752 6 hk_dat_i[19]
port 39 nsew signal input
rlabel metal3 s 523200 96296 524400 96416 6 hk_dat_i[1]
port 40 nsew signal input
rlabel metal3 s 523200 125128 524400 125248 6 hk_dat_i[20]
port 41 nsew signal input
rlabel metal3 s 523200 126624 524400 126744 6 hk_dat_i[21]
port 42 nsew signal input
rlabel metal3 s 523200 128256 524400 128376 6 hk_dat_i[22]
port 43 nsew signal input
rlabel metal3 s 523200 129752 524400 129872 6 hk_dat_i[23]
port 44 nsew signal input
rlabel metal3 s 523200 131248 524400 131368 6 hk_dat_i[24]
port 45 nsew signal input
rlabel metal3 s 523200 132744 524400 132864 6 hk_dat_i[25]
port 46 nsew signal input
rlabel metal3 s 523200 134240 524400 134360 6 hk_dat_i[26]
port 47 nsew signal input
rlabel metal3 s 523200 135736 524400 135856 6 hk_dat_i[27]
port 48 nsew signal input
rlabel metal3 s 523200 137368 524400 137488 6 hk_dat_i[28]
port 49 nsew signal input
rlabel metal3 s 523200 138864 524400 138984 6 hk_dat_i[29]
port 50 nsew signal input
rlabel metal3 s 523200 97792 524400 97912 6 hk_dat_i[2]
port 51 nsew signal input
rlabel metal3 s 523200 140360 524400 140480 6 hk_dat_i[30]
port 52 nsew signal input
rlabel metal3 s 523200 141856 524400 141976 6 hk_dat_i[31]
port 53 nsew signal input
rlabel metal3 s 523200 99288 524400 99408 6 hk_dat_i[3]
port 54 nsew signal input
rlabel metal3 s 523200 100920 524400 101040 6 hk_dat_i[4]
port 55 nsew signal input
rlabel metal3 s 523200 102416 524400 102536 6 hk_dat_i[5]
port 56 nsew signal input
rlabel metal3 s 523200 103912 524400 104032 6 hk_dat_i[6]
port 57 nsew signal input
rlabel metal3 s 523200 105408 524400 105528 6 hk_dat_i[7]
port 58 nsew signal input
rlabel metal3 s 523200 106904 524400 107024 6 hk_dat_i[8]
port 59 nsew signal input
rlabel metal3 s 523200 108400 524400 108520 6 hk_dat_i[9]
port 60 nsew signal input
rlabel metal3 s 523200 93304 524400 93424 6 hk_stb_o
port 61 nsew signal tristate
rlabel metal2 s 521842 163200 521898 164400 6 irq[0]
port 62 nsew signal input
rlabel metal2 s 522670 163200 522726 164400 6 irq[1]
port 63 nsew signal input
rlabel metal2 s 523498 163200 523554 164400 6 irq[2]
port 64 nsew signal input
rlabel metal3 s 523200 75080 524400 75200 6 irq[3]
port 65 nsew signal input
rlabel metal3 s 523200 73584 524400 73704 6 irq[4]
port 66 nsew signal input
rlabel metal3 s 523200 71952 524400 72072 6 irq[5]
port 67 nsew signal input
rlabel metal2 s 386 163200 442 164400 6 la_iena[0]
port 68 nsew signal tristate
rlabel metal2 s 336830 163200 336886 164400 6 la_iena[100]
port 69 nsew signal tristate
rlabel metal2 s 340142 163200 340198 164400 6 la_iena[101]
port 70 nsew signal tristate
rlabel metal2 s 343546 163200 343602 164400 6 la_iena[102]
port 71 nsew signal tristate
rlabel metal2 s 346858 163200 346914 164400 6 la_iena[103]
port 72 nsew signal tristate
rlabel metal2 s 350262 163200 350318 164400 6 la_iena[104]
port 73 nsew signal tristate
rlabel metal2 s 353666 163200 353722 164400 6 la_iena[105]
port 74 nsew signal tristate
rlabel metal2 s 356978 163200 357034 164400 6 la_iena[106]
port 75 nsew signal tristate
rlabel metal2 s 360382 163200 360438 164400 6 la_iena[107]
port 76 nsew signal tristate
rlabel metal2 s 363694 163200 363750 164400 6 la_iena[108]
port 77 nsew signal tristate
rlabel metal2 s 367098 163200 367154 164400 6 la_iena[109]
port 78 nsew signal tristate
rlabel metal2 s 33966 163200 34022 164400 6 la_iena[10]
port 79 nsew signal tristate
rlabel metal2 s 370410 163200 370466 164400 6 la_iena[110]
port 80 nsew signal tristate
rlabel metal2 s 373814 163200 373870 164400 6 la_iena[111]
port 81 nsew signal tristate
rlabel metal2 s 377218 163200 377274 164400 6 la_iena[112]
port 82 nsew signal tristate
rlabel metal2 s 380530 163200 380586 164400 6 la_iena[113]
port 83 nsew signal tristate
rlabel metal2 s 383934 163200 383990 164400 6 la_iena[114]
port 84 nsew signal tristate
rlabel metal2 s 387246 163200 387302 164400 6 la_iena[115]
port 85 nsew signal tristate
rlabel metal2 s 390650 163200 390706 164400 6 la_iena[116]
port 86 nsew signal tristate
rlabel metal2 s 393962 163200 394018 164400 6 la_iena[117]
port 87 nsew signal tristate
rlabel metal2 s 397366 163200 397422 164400 6 la_iena[118]
port 88 nsew signal tristate
rlabel metal2 s 400770 163200 400826 164400 6 la_iena[119]
port 89 nsew signal tristate
rlabel metal2 s 37370 163200 37426 164400 6 la_iena[11]
port 90 nsew signal tristate
rlabel metal2 s 404082 163200 404138 164400 6 la_iena[120]
port 91 nsew signal tristate
rlabel metal2 s 407486 163200 407542 164400 6 la_iena[121]
port 92 nsew signal tristate
rlabel metal2 s 410798 163200 410854 164400 6 la_iena[122]
port 93 nsew signal tristate
rlabel metal2 s 414202 163200 414258 164400 6 la_iena[123]
port 94 nsew signal tristate
rlabel metal2 s 417514 163200 417570 164400 6 la_iena[124]
port 95 nsew signal tristate
rlabel metal2 s 420918 163200 420974 164400 6 la_iena[125]
port 96 nsew signal tristate
rlabel metal2 s 424322 163200 424378 164400 6 la_iena[126]
port 97 nsew signal tristate
rlabel metal2 s 427634 163200 427690 164400 6 la_iena[127]
port 98 nsew signal tristate
rlabel metal2 s 40682 163200 40738 164400 6 la_iena[12]
port 99 nsew signal tristate
rlabel metal2 s 44086 163200 44142 164400 6 la_iena[13]
port 100 nsew signal tristate
rlabel metal2 s 47490 163200 47546 164400 6 la_iena[14]
port 101 nsew signal tristate
rlabel metal2 s 50802 163200 50858 164400 6 la_iena[15]
port 102 nsew signal tristate
rlabel metal2 s 54206 163200 54262 164400 6 la_iena[16]
port 103 nsew signal tristate
rlabel metal2 s 57518 163200 57574 164400 6 la_iena[17]
port 104 nsew signal tristate
rlabel metal2 s 60922 163200 60978 164400 6 la_iena[18]
port 105 nsew signal tristate
rlabel metal2 s 64234 163200 64290 164400 6 la_iena[19]
port 106 nsew signal tristate
rlabel metal2 s 3698 163200 3754 164400 6 la_iena[1]
port 107 nsew signal tristate
rlabel metal2 s 67638 163200 67694 164400 6 la_iena[20]
port 108 nsew signal tristate
rlabel metal2 s 71042 163200 71098 164400 6 la_iena[21]
port 109 nsew signal tristate
rlabel metal2 s 74354 163200 74410 164400 6 la_iena[22]
port 110 nsew signal tristate
rlabel metal2 s 77758 163200 77814 164400 6 la_iena[23]
port 111 nsew signal tristate
rlabel metal2 s 81070 163200 81126 164400 6 la_iena[24]
port 112 nsew signal tristate
rlabel metal2 s 84474 163200 84530 164400 6 la_iena[25]
port 113 nsew signal tristate
rlabel metal2 s 87786 163200 87842 164400 6 la_iena[26]
port 114 nsew signal tristate
rlabel metal2 s 91190 163200 91246 164400 6 la_iena[27]
port 115 nsew signal tristate
rlabel metal2 s 94594 163200 94650 164400 6 la_iena[28]
port 116 nsew signal tristate
rlabel metal2 s 97906 163200 97962 164400 6 la_iena[29]
port 117 nsew signal tristate
rlabel metal2 s 7102 163200 7158 164400 6 la_iena[2]
port 118 nsew signal tristate
rlabel metal2 s 101310 163200 101366 164400 6 la_iena[30]
port 119 nsew signal tristate
rlabel metal2 s 104622 163200 104678 164400 6 la_iena[31]
port 120 nsew signal tristate
rlabel metal2 s 108026 163200 108082 164400 6 la_iena[32]
port 121 nsew signal tristate
rlabel metal2 s 111338 163200 111394 164400 6 la_iena[33]
port 122 nsew signal tristate
rlabel metal2 s 114742 163200 114798 164400 6 la_iena[34]
port 123 nsew signal tristate
rlabel metal2 s 118146 163200 118202 164400 6 la_iena[35]
port 124 nsew signal tristate
rlabel metal2 s 121458 163200 121514 164400 6 la_iena[36]
port 125 nsew signal tristate
rlabel metal2 s 124862 163200 124918 164400 6 la_iena[37]
port 126 nsew signal tristate
rlabel metal2 s 128174 163200 128230 164400 6 la_iena[38]
port 127 nsew signal tristate
rlabel metal2 s 131578 163200 131634 164400 6 la_iena[39]
port 128 nsew signal tristate
rlabel metal2 s 10414 163200 10470 164400 6 la_iena[3]
port 129 nsew signal tristate
rlabel metal2 s 134890 163200 134946 164400 6 la_iena[40]
port 130 nsew signal tristate
rlabel metal2 s 138294 163200 138350 164400 6 la_iena[41]
port 131 nsew signal tristate
rlabel metal2 s 141698 163200 141754 164400 6 la_iena[42]
port 132 nsew signal tristate
rlabel metal2 s 145010 163200 145066 164400 6 la_iena[43]
port 133 nsew signal tristate
rlabel metal2 s 148414 163200 148470 164400 6 la_iena[44]
port 134 nsew signal tristate
rlabel metal2 s 151726 163200 151782 164400 6 la_iena[45]
port 135 nsew signal tristate
rlabel metal2 s 155130 163200 155186 164400 6 la_iena[46]
port 136 nsew signal tristate
rlabel metal2 s 158442 163200 158498 164400 6 la_iena[47]
port 137 nsew signal tristate
rlabel metal2 s 161846 163200 161902 164400 6 la_iena[48]
port 138 nsew signal tristate
rlabel metal2 s 165250 163200 165306 164400 6 la_iena[49]
port 139 nsew signal tristate
rlabel metal2 s 13818 163200 13874 164400 6 la_iena[4]
port 140 nsew signal tristate
rlabel metal2 s 168562 163200 168618 164400 6 la_iena[50]
port 141 nsew signal tristate
rlabel metal2 s 171966 163200 172022 164400 6 la_iena[51]
port 142 nsew signal tristate
rlabel metal2 s 175278 163200 175334 164400 6 la_iena[52]
port 143 nsew signal tristate
rlabel metal2 s 178682 163200 178738 164400 6 la_iena[53]
port 144 nsew signal tristate
rlabel metal2 s 181994 163200 182050 164400 6 la_iena[54]
port 145 nsew signal tristate
rlabel metal2 s 185398 163200 185454 164400 6 la_iena[55]
port 146 nsew signal tristate
rlabel metal2 s 188802 163200 188858 164400 6 la_iena[56]
port 147 nsew signal tristate
rlabel metal2 s 192114 163200 192170 164400 6 la_iena[57]
port 148 nsew signal tristate
rlabel metal2 s 195518 163200 195574 164400 6 la_iena[58]
port 149 nsew signal tristate
rlabel metal2 s 198830 163200 198886 164400 6 la_iena[59]
port 150 nsew signal tristate
rlabel metal2 s 17130 163200 17186 164400 6 la_iena[5]
port 151 nsew signal tristate
rlabel metal2 s 202234 163200 202290 164400 6 la_iena[60]
port 152 nsew signal tristate
rlabel metal2 s 205546 163200 205602 164400 6 la_iena[61]
port 153 nsew signal tristate
rlabel metal2 s 208950 163200 209006 164400 6 la_iena[62]
port 154 nsew signal tristate
rlabel metal2 s 212354 163200 212410 164400 6 la_iena[63]
port 155 nsew signal tristate
rlabel metal2 s 215666 163200 215722 164400 6 la_iena[64]
port 156 nsew signal tristate
rlabel metal2 s 219070 163200 219126 164400 6 la_iena[65]
port 157 nsew signal tristate
rlabel metal2 s 222382 163200 222438 164400 6 la_iena[66]
port 158 nsew signal tristate
rlabel metal2 s 225786 163200 225842 164400 6 la_iena[67]
port 159 nsew signal tristate
rlabel metal2 s 229098 163200 229154 164400 6 la_iena[68]
port 160 nsew signal tristate
rlabel metal2 s 232502 163200 232558 164400 6 la_iena[69]
port 161 nsew signal tristate
rlabel metal2 s 20534 163200 20590 164400 6 la_iena[6]
port 162 nsew signal tristate
rlabel metal2 s 235906 163200 235962 164400 6 la_iena[70]
port 163 nsew signal tristate
rlabel metal2 s 239218 163200 239274 164400 6 la_iena[71]
port 164 nsew signal tristate
rlabel metal2 s 242622 163200 242678 164400 6 la_iena[72]
port 165 nsew signal tristate
rlabel metal2 s 245934 163200 245990 164400 6 la_iena[73]
port 166 nsew signal tristate
rlabel metal2 s 249338 163200 249394 164400 6 la_iena[74]
port 167 nsew signal tristate
rlabel metal2 s 252650 163200 252706 164400 6 la_iena[75]
port 168 nsew signal tristate
rlabel metal2 s 256054 163200 256110 164400 6 la_iena[76]
port 169 nsew signal tristate
rlabel metal2 s 259458 163200 259514 164400 6 la_iena[77]
port 170 nsew signal tristate
rlabel metal2 s 262770 163200 262826 164400 6 la_iena[78]
port 171 nsew signal tristate
rlabel metal2 s 266174 163200 266230 164400 6 la_iena[79]
port 172 nsew signal tristate
rlabel metal2 s 23938 163200 23994 164400 6 la_iena[7]
port 173 nsew signal tristate
rlabel metal2 s 269486 163200 269542 164400 6 la_iena[80]
port 174 nsew signal tristate
rlabel metal2 s 272890 163200 272946 164400 6 la_iena[81]
port 175 nsew signal tristate
rlabel metal2 s 276202 163200 276258 164400 6 la_iena[82]
port 176 nsew signal tristate
rlabel metal2 s 279606 163200 279662 164400 6 la_iena[83]
port 177 nsew signal tristate
rlabel metal2 s 283010 163200 283066 164400 6 la_iena[84]
port 178 nsew signal tristate
rlabel metal2 s 286322 163200 286378 164400 6 la_iena[85]
port 179 nsew signal tristate
rlabel metal2 s 289726 163200 289782 164400 6 la_iena[86]
port 180 nsew signal tristate
rlabel metal2 s 293038 163200 293094 164400 6 la_iena[87]
port 181 nsew signal tristate
rlabel metal2 s 296442 163200 296498 164400 6 la_iena[88]
port 182 nsew signal tristate
rlabel metal2 s 299754 163200 299810 164400 6 la_iena[89]
port 183 nsew signal tristate
rlabel metal2 s 27250 163200 27306 164400 6 la_iena[8]
port 184 nsew signal tristate
rlabel metal2 s 303158 163200 303214 164400 6 la_iena[90]
port 185 nsew signal tristate
rlabel metal2 s 306562 163200 306618 164400 6 la_iena[91]
port 186 nsew signal tristate
rlabel metal2 s 309874 163200 309930 164400 6 la_iena[92]
port 187 nsew signal tristate
rlabel metal2 s 313278 163200 313334 164400 6 la_iena[93]
port 188 nsew signal tristate
rlabel metal2 s 316590 163200 316646 164400 6 la_iena[94]
port 189 nsew signal tristate
rlabel metal2 s 319994 163200 320050 164400 6 la_iena[95]
port 190 nsew signal tristate
rlabel metal2 s 323306 163200 323362 164400 6 la_iena[96]
port 191 nsew signal tristate
rlabel metal2 s 326710 163200 326766 164400 6 la_iena[97]
port 192 nsew signal tristate
rlabel metal2 s 330114 163200 330170 164400 6 la_iena[98]
port 193 nsew signal tristate
rlabel metal2 s 333426 163200 333482 164400 6 la_iena[99]
port 194 nsew signal tristate
rlabel metal2 s 30654 163200 30710 164400 6 la_iena[9]
port 195 nsew signal tristate
rlabel metal2 s 1214 163200 1270 164400 6 la_input[0]
port 196 nsew signal input
rlabel metal2 s 337658 163200 337714 164400 6 la_input[100]
port 197 nsew signal input
rlabel metal2 s 340970 163200 341026 164400 6 la_input[101]
port 198 nsew signal input
rlabel metal2 s 344374 163200 344430 164400 6 la_input[102]
port 199 nsew signal input
rlabel metal2 s 347778 163200 347834 164400 6 la_input[103]
port 200 nsew signal input
rlabel metal2 s 351090 163200 351146 164400 6 la_input[104]
port 201 nsew signal input
rlabel metal2 s 354494 163200 354550 164400 6 la_input[105]
port 202 nsew signal input
rlabel metal2 s 357806 163200 357862 164400 6 la_input[106]
port 203 nsew signal input
rlabel metal2 s 361210 163200 361266 164400 6 la_input[107]
port 204 nsew signal input
rlabel metal2 s 364522 163200 364578 164400 6 la_input[108]
port 205 nsew signal input
rlabel metal2 s 367926 163200 367982 164400 6 la_input[109]
port 206 nsew signal input
rlabel metal2 s 34794 163200 34850 164400 6 la_input[10]
port 207 nsew signal input
rlabel metal2 s 371330 163200 371386 164400 6 la_input[110]
port 208 nsew signal input
rlabel metal2 s 374642 163200 374698 164400 6 la_input[111]
port 209 nsew signal input
rlabel metal2 s 378046 163200 378102 164400 6 la_input[112]
port 210 nsew signal input
rlabel metal2 s 381358 163200 381414 164400 6 la_input[113]
port 211 nsew signal input
rlabel metal2 s 384762 163200 384818 164400 6 la_input[114]
port 212 nsew signal input
rlabel metal2 s 388074 163200 388130 164400 6 la_input[115]
port 213 nsew signal input
rlabel metal2 s 391478 163200 391534 164400 6 la_input[116]
port 214 nsew signal input
rlabel metal2 s 394882 163200 394938 164400 6 la_input[117]
port 215 nsew signal input
rlabel metal2 s 398194 163200 398250 164400 6 la_input[118]
port 216 nsew signal input
rlabel metal2 s 401598 163200 401654 164400 6 la_input[119]
port 217 nsew signal input
rlabel metal2 s 38198 163200 38254 164400 6 la_input[11]
port 218 nsew signal input
rlabel metal2 s 404910 163200 404966 164400 6 la_input[120]
port 219 nsew signal input
rlabel metal2 s 408314 163200 408370 164400 6 la_input[121]
port 220 nsew signal input
rlabel metal2 s 411626 163200 411682 164400 6 la_input[122]
port 221 nsew signal input
rlabel metal2 s 415030 163200 415086 164400 6 la_input[123]
port 222 nsew signal input
rlabel metal2 s 418434 163200 418490 164400 6 la_input[124]
port 223 nsew signal input
rlabel metal2 s 421746 163200 421802 164400 6 la_input[125]
port 224 nsew signal input
rlabel metal2 s 425150 163200 425206 164400 6 la_input[126]
port 225 nsew signal input
rlabel metal2 s 428462 163200 428518 164400 6 la_input[127]
port 226 nsew signal input
rlabel metal2 s 41602 163200 41658 164400 6 la_input[12]
port 227 nsew signal input
rlabel metal2 s 44914 163200 44970 164400 6 la_input[13]
port 228 nsew signal input
rlabel metal2 s 48318 163200 48374 164400 6 la_input[14]
port 229 nsew signal input
rlabel metal2 s 51630 163200 51686 164400 6 la_input[15]
port 230 nsew signal input
rlabel metal2 s 55034 163200 55090 164400 6 la_input[16]
port 231 nsew signal input
rlabel metal2 s 58346 163200 58402 164400 6 la_input[17]
port 232 nsew signal input
rlabel metal2 s 61750 163200 61806 164400 6 la_input[18]
port 233 nsew signal input
rlabel metal2 s 65154 163200 65210 164400 6 la_input[19]
port 234 nsew signal input
rlabel metal2 s 4526 163200 4582 164400 6 la_input[1]
port 235 nsew signal input
rlabel metal2 s 68466 163200 68522 164400 6 la_input[20]
port 236 nsew signal input
rlabel metal2 s 71870 163200 71926 164400 6 la_input[21]
port 237 nsew signal input
rlabel metal2 s 75182 163200 75238 164400 6 la_input[22]
port 238 nsew signal input
rlabel metal2 s 78586 163200 78642 164400 6 la_input[23]
port 239 nsew signal input
rlabel metal2 s 81898 163200 81954 164400 6 la_input[24]
port 240 nsew signal input
rlabel metal2 s 85302 163200 85358 164400 6 la_input[25]
port 241 nsew signal input
rlabel metal2 s 88706 163200 88762 164400 6 la_input[26]
port 242 nsew signal input
rlabel metal2 s 92018 163200 92074 164400 6 la_input[27]
port 243 nsew signal input
rlabel metal2 s 95422 163200 95478 164400 6 la_input[28]
port 244 nsew signal input
rlabel metal2 s 98734 163200 98790 164400 6 la_input[29]
port 245 nsew signal input
rlabel metal2 s 7930 163200 7986 164400 6 la_input[2]
port 246 nsew signal input
rlabel metal2 s 102138 163200 102194 164400 6 la_input[30]
port 247 nsew signal input
rlabel metal2 s 105450 163200 105506 164400 6 la_input[31]
port 248 nsew signal input
rlabel metal2 s 108854 163200 108910 164400 6 la_input[32]
port 249 nsew signal input
rlabel metal2 s 112258 163200 112314 164400 6 la_input[33]
port 250 nsew signal input
rlabel metal2 s 115570 163200 115626 164400 6 la_input[34]
port 251 nsew signal input
rlabel metal2 s 118974 163200 119030 164400 6 la_input[35]
port 252 nsew signal input
rlabel metal2 s 122286 163200 122342 164400 6 la_input[36]
port 253 nsew signal input
rlabel metal2 s 125690 163200 125746 164400 6 la_input[37]
port 254 nsew signal input
rlabel metal2 s 129002 163200 129058 164400 6 la_input[38]
port 255 nsew signal input
rlabel metal2 s 132406 163200 132462 164400 6 la_input[39]
port 256 nsew signal input
rlabel metal2 s 11242 163200 11298 164400 6 la_input[3]
port 257 nsew signal input
rlabel metal2 s 135810 163200 135866 164400 6 la_input[40]
port 258 nsew signal input
rlabel metal2 s 139122 163200 139178 164400 6 la_input[41]
port 259 nsew signal input
rlabel metal2 s 142526 163200 142582 164400 6 la_input[42]
port 260 nsew signal input
rlabel metal2 s 145838 163200 145894 164400 6 la_input[43]
port 261 nsew signal input
rlabel metal2 s 149242 163200 149298 164400 6 la_input[44]
port 262 nsew signal input
rlabel metal2 s 152554 163200 152610 164400 6 la_input[45]
port 263 nsew signal input
rlabel metal2 s 155958 163200 156014 164400 6 la_input[46]
port 264 nsew signal input
rlabel metal2 s 159362 163200 159418 164400 6 la_input[47]
port 265 nsew signal input
rlabel metal2 s 162674 163200 162730 164400 6 la_input[48]
port 266 nsew signal input
rlabel metal2 s 166078 163200 166134 164400 6 la_input[49]
port 267 nsew signal input
rlabel metal2 s 14646 163200 14702 164400 6 la_input[4]
port 268 nsew signal input
rlabel metal2 s 169390 163200 169446 164400 6 la_input[50]
port 269 nsew signal input
rlabel metal2 s 172794 163200 172850 164400 6 la_input[51]
port 270 nsew signal input
rlabel metal2 s 176106 163200 176162 164400 6 la_input[52]
port 271 nsew signal input
rlabel metal2 s 179510 163200 179566 164400 6 la_input[53]
port 272 nsew signal input
rlabel metal2 s 182914 163200 182970 164400 6 la_input[54]
port 273 nsew signal input
rlabel metal2 s 186226 163200 186282 164400 6 la_input[55]
port 274 nsew signal input
rlabel metal2 s 189630 163200 189686 164400 6 la_input[56]
port 275 nsew signal input
rlabel metal2 s 192942 163200 192998 164400 6 la_input[57]
port 276 nsew signal input
rlabel metal2 s 196346 163200 196402 164400 6 la_input[58]
port 277 nsew signal input
rlabel metal2 s 199658 163200 199714 164400 6 la_input[59]
port 278 nsew signal input
rlabel metal2 s 18050 163200 18106 164400 6 la_input[5]
port 279 nsew signal input
rlabel metal2 s 203062 163200 203118 164400 6 la_input[60]
port 280 nsew signal input
rlabel metal2 s 206466 163200 206522 164400 6 la_input[61]
port 281 nsew signal input
rlabel metal2 s 209778 163200 209834 164400 6 la_input[62]
port 282 nsew signal input
rlabel metal2 s 213182 163200 213238 164400 6 la_input[63]
port 283 nsew signal input
rlabel metal2 s 216494 163200 216550 164400 6 la_input[64]
port 284 nsew signal input
rlabel metal2 s 219898 163200 219954 164400 6 la_input[65]
port 285 nsew signal input
rlabel metal2 s 223210 163200 223266 164400 6 la_input[66]
port 286 nsew signal input
rlabel metal2 s 226614 163200 226670 164400 6 la_input[67]
port 287 nsew signal input
rlabel metal2 s 230018 163200 230074 164400 6 la_input[68]
port 288 nsew signal input
rlabel metal2 s 233330 163200 233386 164400 6 la_input[69]
port 289 nsew signal input
rlabel metal2 s 21362 163200 21418 164400 6 la_input[6]
port 290 nsew signal input
rlabel metal2 s 236734 163200 236790 164400 6 la_input[70]
port 291 nsew signal input
rlabel metal2 s 240046 163200 240102 164400 6 la_input[71]
port 292 nsew signal input
rlabel metal2 s 243450 163200 243506 164400 6 la_input[72]
port 293 nsew signal input
rlabel metal2 s 246762 163200 246818 164400 6 la_input[73]
port 294 nsew signal input
rlabel metal2 s 250166 163200 250222 164400 6 la_input[74]
port 295 nsew signal input
rlabel metal2 s 253570 163200 253626 164400 6 la_input[75]
port 296 nsew signal input
rlabel metal2 s 256882 163200 256938 164400 6 la_input[76]
port 297 nsew signal input
rlabel metal2 s 260286 163200 260342 164400 6 la_input[77]
port 298 nsew signal input
rlabel metal2 s 263598 163200 263654 164400 6 la_input[78]
port 299 nsew signal input
rlabel metal2 s 267002 163200 267058 164400 6 la_input[79]
port 300 nsew signal input
rlabel metal2 s 24766 163200 24822 164400 6 la_input[7]
port 301 nsew signal input
rlabel metal2 s 270314 163200 270370 164400 6 la_input[80]
port 302 nsew signal input
rlabel metal2 s 273718 163200 273774 164400 6 la_input[81]
port 303 nsew signal input
rlabel metal2 s 277122 163200 277178 164400 6 la_input[82]
port 304 nsew signal input
rlabel metal2 s 280434 163200 280490 164400 6 la_input[83]
port 305 nsew signal input
rlabel metal2 s 283838 163200 283894 164400 6 la_input[84]
port 306 nsew signal input
rlabel metal2 s 287150 163200 287206 164400 6 la_input[85]
port 307 nsew signal input
rlabel metal2 s 290554 163200 290610 164400 6 la_input[86]
port 308 nsew signal input
rlabel metal2 s 293866 163200 293922 164400 6 la_input[87]
port 309 nsew signal input
rlabel metal2 s 297270 163200 297326 164400 6 la_input[88]
port 310 nsew signal input
rlabel metal2 s 300674 163200 300730 164400 6 la_input[89]
port 311 nsew signal input
rlabel metal2 s 28078 163200 28134 164400 6 la_input[8]
port 312 nsew signal input
rlabel metal2 s 303986 163200 304042 164400 6 la_input[90]
port 313 nsew signal input
rlabel metal2 s 307390 163200 307446 164400 6 la_input[91]
port 314 nsew signal input
rlabel metal2 s 310702 163200 310758 164400 6 la_input[92]
port 315 nsew signal input
rlabel metal2 s 314106 163200 314162 164400 6 la_input[93]
port 316 nsew signal input
rlabel metal2 s 317418 163200 317474 164400 6 la_input[94]
port 317 nsew signal input
rlabel metal2 s 320822 163200 320878 164400 6 la_input[95]
port 318 nsew signal input
rlabel metal2 s 324226 163200 324282 164400 6 la_input[96]
port 319 nsew signal input
rlabel metal2 s 327538 163200 327594 164400 6 la_input[97]
port 320 nsew signal input
rlabel metal2 s 330942 163200 330998 164400 6 la_input[98]
port 321 nsew signal input
rlabel metal2 s 334254 163200 334310 164400 6 la_input[99]
port 322 nsew signal input
rlabel metal2 s 31482 163200 31538 164400 6 la_input[9]
port 323 nsew signal input
rlabel metal2 s 2042 163200 2098 164400 6 la_oenb[0]
port 324 nsew signal tristate
rlabel metal2 s 338486 163200 338542 164400 6 la_oenb[100]
port 325 nsew signal tristate
rlabel metal2 s 341890 163200 341946 164400 6 la_oenb[101]
port 326 nsew signal tristate
rlabel metal2 s 345202 163200 345258 164400 6 la_oenb[102]
port 327 nsew signal tristate
rlabel metal2 s 348606 163200 348662 164400 6 la_oenb[103]
port 328 nsew signal tristate
rlabel metal2 s 351918 163200 351974 164400 6 la_oenb[104]
port 329 nsew signal tristate
rlabel metal2 s 355322 163200 355378 164400 6 la_oenb[105]
port 330 nsew signal tristate
rlabel metal2 s 358634 163200 358690 164400 6 la_oenb[106]
port 331 nsew signal tristate
rlabel metal2 s 362038 163200 362094 164400 6 la_oenb[107]
port 332 nsew signal tristate
rlabel metal2 s 365442 163200 365498 164400 6 la_oenb[108]
port 333 nsew signal tristate
rlabel metal2 s 368754 163200 368810 164400 6 la_oenb[109]
port 334 nsew signal tristate
rlabel metal2 s 35714 163200 35770 164400 6 la_oenb[10]
port 335 nsew signal tristate
rlabel metal2 s 372158 163200 372214 164400 6 la_oenb[110]
port 336 nsew signal tristate
rlabel metal2 s 375470 163200 375526 164400 6 la_oenb[111]
port 337 nsew signal tristate
rlabel metal2 s 378874 163200 378930 164400 6 la_oenb[112]
port 338 nsew signal tristate
rlabel metal2 s 382186 163200 382242 164400 6 la_oenb[113]
port 339 nsew signal tristate
rlabel metal2 s 385590 163200 385646 164400 6 la_oenb[114]
port 340 nsew signal tristate
rlabel metal2 s 388994 163200 389050 164400 6 la_oenb[115]
port 341 nsew signal tristate
rlabel metal2 s 392306 163200 392362 164400 6 la_oenb[116]
port 342 nsew signal tristate
rlabel metal2 s 395710 163200 395766 164400 6 la_oenb[117]
port 343 nsew signal tristate
rlabel metal2 s 399022 163200 399078 164400 6 la_oenb[118]
port 344 nsew signal tristate
rlabel metal2 s 402426 163200 402482 164400 6 la_oenb[119]
port 345 nsew signal tristate
rlabel metal2 s 39026 163200 39082 164400 6 la_oenb[11]
port 346 nsew signal tristate
rlabel metal2 s 405738 163200 405794 164400 6 la_oenb[120]
port 347 nsew signal tristate
rlabel metal2 s 409142 163200 409198 164400 6 la_oenb[121]
port 348 nsew signal tristate
rlabel metal2 s 412546 163200 412602 164400 6 la_oenb[122]
port 349 nsew signal tristate
rlabel metal2 s 415858 163200 415914 164400 6 la_oenb[123]
port 350 nsew signal tristate
rlabel metal2 s 419262 163200 419318 164400 6 la_oenb[124]
port 351 nsew signal tristate
rlabel metal2 s 422574 163200 422630 164400 6 la_oenb[125]
port 352 nsew signal tristate
rlabel metal2 s 425978 163200 426034 164400 6 la_oenb[126]
port 353 nsew signal tristate
rlabel metal2 s 429290 163200 429346 164400 6 la_oenb[127]
port 354 nsew signal tristate
rlabel metal2 s 42430 163200 42486 164400 6 la_oenb[12]
port 355 nsew signal tristate
rlabel metal2 s 45742 163200 45798 164400 6 la_oenb[13]
port 356 nsew signal tristate
rlabel metal2 s 49146 163200 49202 164400 6 la_oenb[14]
port 357 nsew signal tristate
rlabel metal2 s 52458 163200 52514 164400 6 la_oenb[15]
port 358 nsew signal tristate
rlabel metal2 s 55862 163200 55918 164400 6 la_oenb[16]
port 359 nsew signal tristate
rlabel metal2 s 59266 163200 59322 164400 6 la_oenb[17]
port 360 nsew signal tristate
rlabel metal2 s 62578 163200 62634 164400 6 la_oenb[18]
port 361 nsew signal tristate
rlabel metal2 s 65982 163200 66038 164400 6 la_oenb[19]
port 362 nsew signal tristate
rlabel metal2 s 5354 163200 5410 164400 6 la_oenb[1]
port 363 nsew signal tristate
rlabel metal2 s 69294 163200 69350 164400 6 la_oenb[20]
port 364 nsew signal tristate
rlabel metal2 s 72698 163200 72754 164400 6 la_oenb[21]
port 365 nsew signal tristate
rlabel metal2 s 76010 163200 76066 164400 6 la_oenb[22]
port 366 nsew signal tristate
rlabel metal2 s 79414 163200 79470 164400 6 la_oenb[23]
port 367 nsew signal tristate
rlabel metal2 s 82818 163200 82874 164400 6 la_oenb[24]
port 368 nsew signal tristate
rlabel metal2 s 86130 163200 86186 164400 6 la_oenb[25]
port 369 nsew signal tristate
rlabel metal2 s 89534 163200 89590 164400 6 la_oenb[26]
port 370 nsew signal tristate
rlabel metal2 s 92846 163200 92902 164400 6 la_oenb[27]
port 371 nsew signal tristate
rlabel metal2 s 96250 163200 96306 164400 6 la_oenb[28]
port 372 nsew signal tristate
rlabel metal2 s 99562 163200 99618 164400 6 la_oenb[29]
port 373 nsew signal tristate
rlabel metal2 s 8758 163200 8814 164400 6 la_oenb[2]
port 374 nsew signal tristate
rlabel metal2 s 102966 163200 103022 164400 6 la_oenb[30]
port 375 nsew signal tristate
rlabel metal2 s 106370 163200 106426 164400 6 la_oenb[31]
port 376 nsew signal tristate
rlabel metal2 s 109682 163200 109738 164400 6 la_oenb[32]
port 377 nsew signal tristate
rlabel metal2 s 113086 163200 113142 164400 6 la_oenb[33]
port 378 nsew signal tristate
rlabel metal2 s 116398 163200 116454 164400 6 la_oenb[34]
port 379 nsew signal tristate
rlabel metal2 s 119802 163200 119858 164400 6 la_oenb[35]
port 380 nsew signal tristate
rlabel metal2 s 123114 163200 123170 164400 6 la_oenb[36]
port 381 nsew signal tristate
rlabel metal2 s 126518 163200 126574 164400 6 la_oenb[37]
port 382 nsew signal tristate
rlabel metal2 s 129922 163200 129978 164400 6 la_oenb[38]
port 383 nsew signal tristate
rlabel metal2 s 133234 163200 133290 164400 6 la_oenb[39]
port 384 nsew signal tristate
rlabel metal2 s 12162 163200 12218 164400 6 la_oenb[3]
port 385 nsew signal tristate
rlabel metal2 s 136638 163200 136694 164400 6 la_oenb[40]
port 386 nsew signal tristate
rlabel metal2 s 139950 163200 140006 164400 6 la_oenb[41]
port 387 nsew signal tristate
rlabel metal2 s 143354 163200 143410 164400 6 la_oenb[42]
port 388 nsew signal tristate
rlabel metal2 s 146666 163200 146722 164400 6 la_oenb[43]
port 389 nsew signal tristate
rlabel metal2 s 150070 163200 150126 164400 6 la_oenb[44]
port 390 nsew signal tristate
rlabel metal2 s 153474 163200 153530 164400 6 la_oenb[45]
port 391 nsew signal tristate
rlabel metal2 s 156786 163200 156842 164400 6 la_oenb[46]
port 392 nsew signal tristate
rlabel metal2 s 160190 163200 160246 164400 6 la_oenb[47]
port 393 nsew signal tristate
rlabel metal2 s 163502 163200 163558 164400 6 la_oenb[48]
port 394 nsew signal tristate
rlabel metal2 s 166906 163200 166962 164400 6 la_oenb[49]
port 395 nsew signal tristate
rlabel metal2 s 15474 163200 15530 164400 6 la_oenb[4]
port 396 nsew signal tristate
rlabel metal2 s 170218 163200 170274 164400 6 la_oenb[50]
port 397 nsew signal tristate
rlabel metal2 s 173622 163200 173678 164400 6 la_oenb[51]
port 398 nsew signal tristate
rlabel metal2 s 177026 163200 177082 164400 6 la_oenb[52]
port 399 nsew signal tristate
rlabel metal2 s 180338 163200 180394 164400 6 la_oenb[53]
port 400 nsew signal tristate
rlabel metal2 s 183742 163200 183798 164400 6 la_oenb[54]
port 401 nsew signal tristate
rlabel metal2 s 187054 163200 187110 164400 6 la_oenb[55]
port 402 nsew signal tristate
rlabel metal2 s 190458 163200 190514 164400 6 la_oenb[56]
port 403 nsew signal tristate
rlabel metal2 s 193770 163200 193826 164400 6 la_oenb[57]
port 404 nsew signal tristate
rlabel metal2 s 197174 163200 197230 164400 6 la_oenb[58]
port 405 nsew signal tristate
rlabel metal2 s 200578 163200 200634 164400 6 la_oenb[59]
port 406 nsew signal tristate
rlabel metal2 s 18878 163200 18934 164400 6 la_oenb[5]
port 407 nsew signal tristate
rlabel metal2 s 203890 163200 203946 164400 6 la_oenb[60]
port 408 nsew signal tristate
rlabel metal2 s 207294 163200 207350 164400 6 la_oenb[61]
port 409 nsew signal tristate
rlabel metal2 s 210606 163200 210662 164400 6 la_oenb[62]
port 410 nsew signal tristate
rlabel metal2 s 214010 163200 214066 164400 6 la_oenb[63]
port 411 nsew signal tristate
rlabel metal2 s 217322 163200 217378 164400 6 la_oenb[64]
port 412 nsew signal tristate
rlabel metal2 s 220726 163200 220782 164400 6 la_oenb[65]
port 413 nsew signal tristate
rlabel metal2 s 224130 163200 224186 164400 6 la_oenb[66]
port 414 nsew signal tristate
rlabel metal2 s 227442 163200 227498 164400 6 la_oenb[67]
port 415 nsew signal tristate
rlabel metal2 s 230846 163200 230902 164400 6 la_oenb[68]
port 416 nsew signal tristate
rlabel metal2 s 234158 163200 234214 164400 6 la_oenb[69]
port 417 nsew signal tristate
rlabel metal2 s 22190 163200 22246 164400 6 la_oenb[6]
port 418 nsew signal tristate
rlabel metal2 s 237562 163200 237618 164400 6 la_oenb[70]
port 419 nsew signal tristate
rlabel metal2 s 240874 163200 240930 164400 6 la_oenb[71]
port 420 nsew signal tristate
rlabel metal2 s 244278 163200 244334 164400 6 la_oenb[72]
port 421 nsew signal tristate
rlabel metal2 s 247682 163200 247738 164400 6 la_oenb[73]
port 422 nsew signal tristate
rlabel metal2 s 250994 163200 251050 164400 6 la_oenb[74]
port 423 nsew signal tristate
rlabel metal2 s 254398 163200 254454 164400 6 la_oenb[75]
port 424 nsew signal tristate
rlabel metal2 s 257710 163200 257766 164400 6 la_oenb[76]
port 425 nsew signal tristate
rlabel metal2 s 261114 163200 261170 164400 6 la_oenb[77]
port 426 nsew signal tristate
rlabel metal2 s 264426 163200 264482 164400 6 la_oenb[78]
port 427 nsew signal tristate
rlabel metal2 s 267830 163200 267886 164400 6 la_oenb[79]
port 428 nsew signal tristate
rlabel metal2 s 25594 163200 25650 164400 6 la_oenb[7]
port 429 nsew signal tristate
rlabel metal2 s 271234 163200 271290 164400 6 la_oenb[80]
port 430 nsew signal tristate
rlabel metal2 s 274546 163200 274602 164400 6 la_oenb[81]
port 431 nsew signal tristate
rlabel metal2 s 277950 163200 278006 164400 6 la_oenb[82]
port 432 nsew signal tristate
rlabel metal2 s 281262 163200 281318 164400 6 la_oenb[83]
port 433 nsew signal tristate
rlabel metal2 s 284666 163200 284722 164400 6 la_oenb[84]
port 434 nsew signal tristate
rlabel metal2 s 287978 163200 288034 164400 6 la_oenb[85]
port 435 nsew signal tristate
rlabel metal2 s 291382 163200 291438 164400 6 la_oenb[86]
port 436 nsew signal tristate
rlabel metal2 s 294786 163200 294842 164400 6 la_oenb[87]
port 437 nsew signal tristate
rlabel metal2 s 298098 163200 298154 164400 6 la_oenb[88]
port 438 nsew signal tristate
rlabel metal2 s 301502 163200 301558 164400 6 la_oenb[89]
port 439 nsew signal tristate
rlabel metal2 s 28906 163200 28962 164400 6 la_oenb[8]
port 440 nsew signal tristate
rlabel metal2 s 304814 163200 304870 164400 6 la_oenb[90]
port 441 nsew signal tristate
rlabel metal2 s 308218 163200 308274 164400 6 la_oenb[91]
port 442 nsew signal tristate
rlabel metal2 s 311530 163200 311586 164400 6 la_oenb[92]
port 443 nsew signal tristate
rlabel metal2 s 314934 163200 314990 164400 6 la_oenb[93]
port 444 nsew signal tristate
rlabel metal2 s 318338 163200 318394 164400 6 la_oenb[94]
port 445 nsew signal tristate
rlabel metal2 s 321650 163200 321706 164400 6 la_oenb[95]
port 446 nsew signal tristate
rlabel metal2 s 325054 163200 325110 164400 6 la_oenb[96]
port 447 nsew signal tristate
rlabel metal2 s 328366 163200 328422 164400 6 la_oenb[97]
port 448 nsew signal tristate
rlabel metal2 s 331770 163200 331826 164400 6 la_oenb[98]
port 449 nsew signal tristate
rlabel metal2 s 335082 163200 335138 164400 6 la_oenb[99]
port 450 nsew signal tristate
rlabel metal2 s 32310 163200 32366 164400 6 la_oenb[9]
port 451 nsew signal tristate
rlabel metal2 s 2870 163200 2926 164400 6 la_output[0]
port 452 nsew signal tristate
rlabel metal2 s 339314 163200 339370 164400 6 la_output[100]
port 453 nsew signal tristate
rlabel metal2 s 342718 163200 342774 164400 6 la_output[101]
port 454 nsew signal tristate
rlabel metal2 s 346030 163200 346086 164400 6 la_output[102]
port 455 nsew signal tristate
rlabel metal2 s 349434 163200 349490 164400 6 la_output[103]
port 456 nsew signal tristate
rlabel metal2 s 352746 163200 352802 164400 6 la_output[104]
port 457 nsew signal tristate
rlabel metal2 s 356150 163200 356206 164400 6 la_output[105]
port 458 nsew signal tristate
rlabel metal2 s 359554 163200 359610 164400 6 la_output[106]
port 459 nsew signal tristate
rlabel metal2 s 362866 163200 362922 164400 6 la_output[107]
port 460 nsew signal tristate
rlabel metal2 s 366270 163200 366326 164400 6 la_output[108]
port 461 nsew signal tristate
rlabel metal2 s 369582 163200 369638 164400 6 la_output[109]
port 462 nsew signal tristate
rlabel metal2 s 36542 163200 36598 164400 6 la_output[10]
port 463 nsew signal tristate
rlabel metal2 s 372986 163200 373042 164400 6 la_output[110]
port 464 nsew signal tristate
rlabel metal2 s 376298 163200 376354 164400 6 la_output[111]
port 465 nsew signal tristate
rlabel metal2 s 379702 163200 379758 164400 6 la_output[112]
port 466 nsew signal tristate
rlabel metal2 s 383106 163200 383162 164400 6 la_output[113]
port 467 nsew signal tristate
rlabel metal2 s 386418 163200 386474 164400 6 la_output[114]
port 468 nsew signal tristate
rlabel metal2 s 389822 163200 389878 164400 6 la_output[115]
port 469 nsew signal tristate
rlabel metal2 s 393134 163200 393190 164400 6 la_output[116]
port 470 nsew signal tristate
rlabel metal2 s 396538 163200 396594 164400 6 la_output[117]
port 471 nsew signal tristate
rlabel metal2 s 399850 163200 399906 164400 6 la_output[118]
port 472 nsew signal tristate
rlabel metal2 s 403254 163200 403310 164400 6 la_output[119]
port 473 nsew signal tristate
rlabel metal2 s 39854 163200 39910 164400 6 la_output[11]
port 474 nsew signal tristate
rlabel metal2 s 406658 163200 406714 164400 6 la_output[120]
port 475 nsew signal tristate
rlabel metal2 s 409970 163200 410026 164400 6 la_output[121]
port 476 nsew signal tristate
rlabel metal2 s 413374 163200 413430 164400 6 la_output[122]
port 477 nsew signal tristate
rlabel metal2 s 416686 163200 416742 164400 6 la_output[123]
port 478 nsew signal tristate
rlabel metal2 s 420090 163200 420146 164400 6 la_output[124]
port 479 nsew signal tristate
rlabel metal2 s 423402 163200 423458 164400 6 la_output[125]
port 480 nsew signal tristate
rlabel metal2 s 426806 163200 426862 164400 6 la_output[126]
port 481 nsew signal tristate
rlabel metal2 s 430210 163200 430266 164400 6 la_output[127]
port 482 nsew signal tristate
rlabel metal2 s 43258 163200 43314 164400 6 la_output[12]
port 483 nsew signal tristate
rlabel metal2 s 46570 163200 46626 164400 6 la_output[13]
port 484 nsew signal tristate
rlabel metal2 s 49974 163200 50030 164400 6 la_output[14]
port 485 nsew signal tristate
rlabel metal2 s 53378 163200 53434 164400 6 la_output[15]
port 486 nsew signal tristate
rlabel metal2 s 56690 163200 56746 164400 6 la_output[16]
port 487 nsew signal tristate
rlabel metal2 s 60094 163200 60150 164400 6 la_output[17]
port 488 nsew signal tristate
rlabel metal2 s 63406 163200 63462 164400 6 la_output[18]
port 489 nsew signal tristate
rlabel metal2 s 66810 163200 66866 164400 6 la_output[19]
port 490 nsew signal tristate
rlabel metal2 s 6274 163200 6330 164400 6 la_output[1]
port 491 nsew signal tristate
rlabel metal2 s 70122 163200 70178 164400 6 la_output[20]
port 492 nsew signal tristate
rlabel metal2 s 73526 163200 73582 164400 6 la_output[21]
port 493 nsew signal tristate
rlabel metal2 s 76930 163200 76986 164400 6 la_output[22]
port 494 nsew signal tristate
rlabel metal2 s 80242 163200 80298 164400 6 la_output[23]
port 495 nsew signal tristate
rlabel metal2 s 83646 163200 83702 164400 6 la_output[24]
port 496 nsew signal tristate
rlabel metal2 s 86958 163200 87014 164400 6 la_output[25]
port 497 nsew signal tristate
rlabel metal2 s 90362 163200 90418 164400 6 la_output[26]
port 498 nsew signal tristate
rlabel metal2 s 93674 163200 93730 164400 6 la_output[27]
port 499 nsew signal tristate
rlabel metal2 s 97078 163200 97134 164400 6 la_output[28]
port 500 nsew signal tristate
rlabel metal2 s 100482 163200 100538 164400 6 la_output[29]
port 501 nsew signal tristate
rlabel metal2 s 9586 163200 9642 164400 6 la_output[2]
port 502 nsew signal tristate
rlabel metal2 s 103794 163200 103850 164400 6 la_output[30]
port 503 nsew signal tristate
rlabel metal2 s 107198 163200 107254 164400 6 la_output[31]
port 504 nsew signal tristate
rlabel metal2 s 110510 163200 110566 164400 6 la_output[32]
port 505 nsew signal tristate
rlabel metal2 s 113914 163200 113970 164400 6 la_output[33]
port 506 nsew signal tristate
rlabel metal2 s 117226 163200 117282 164400 6 la_output[34]
port 507 nsew signal tristate
rlabel metal2 s 120630 163200 120686 164400 6 la_output[35]
port 508 nsew signal tristate
rlabel metal2 s 124034 163200 124090 164400 6 la_output[36]
port 509 nsew signal tristate
rlabel metal2 s 127346 163200 127402 164400 6 la_output[37]
port 510 nsew signal tristate
rlabel metal2 s 130750 163200 130806 164400 6 la_output[38]
port 511 nsew signal tristate
rlabel metal2 s 134062 163200 134118 164400 6 la_output[39]
port 512 nsew signal tristate
rlabel metal2 s 12990 163200 13046 164400 6 la_output[3]
port 513 nsew signal tristate
rlabel metal2 s 137466 163200 137522 164400 6 la_output[40]
port 514 nsew signal tristate
rlabel metal2 s 140778 163200 140834 164400 6 la_output[41]
port 515 nsew signal tristate
rlabel metal2 s 144182 163200 144238 164400 6 la_output[42]
port 516 nsew signal tristate
rlabel metal2 s 147586 163200 147642 164400 6 la_output[43]
port 517 nsew signal tristate
rlabel metal2 s 150898 163200 150954 164400 6 la_output[44]
port 518 nsew signal tristate
rlabel metal2 s 154302 163200 154358 164400 6 la_output[45]
port 519 nsew signal tristate
rlabel metal2 s 157614 163200 157670 164400 6 la_output[46]
port 520 nsew signal tristate
rlabel metal2 s 161018 163200 161074 164400 6 la_output[47]
port 521 nsew signal tristate
rlabel metal2 s 164330 163200 164386 164400 6 la_output[48]
port 522 nsew signal tristate
rlabel metal2 s 167734 163200 167790 164400 6 la_output[49]
port 523 nsew signal tristate
rlabel metal2 s 16302 163200 16358 164400 6 la_output[4]
port 524 nsew signal tristate
rlabel metal2 s 171138 163200 171194 164400 6 la_output[50]
port 525 nsew signal tristate
rlabel metal2 s 174450 163200 174506 164400 6 la_output[51]
port 526 nsew signal tristate
rlabel metal2 s 177854 163200 177910 164400 6 la_output[52]
port 527 nsew signal tristate
rlabel metal2 s 181166 163200 181222 164400 6 la_output[53]
port 528 nsew signal tristate
rlabel metal2 s 184570 163200 184626 164400 6 la_output[54]
port 529 nsew signal tristate
rlabel metal2 s 187882 163200 187938 164400 6 la_output[55]
port 530 nsew signal tristate
rlabel metal2 s 191286 163200 191342 164400 6 la_output[56]
port 531 nsew signal tristate
rlabel metal2 s 194690 163200 194746 164400 6 la_output[57]
port 532 nsew signal tristate
rlabel metal2 s 198002 163200 198058 164400 6 la_output[58]
port 533 nsew signal tristate
rlabel metal2 s 201406 163200 201462 164400 6 la_output[59]
port 534 nsew signal tristate
rlabel metal2 s 19706 163200 19762 164400 6 la_output[5]
port 535 nsew signal tristate
rlabel metal2 s 204718 163200 204774 164400 6 la_output[60]
port 536 nsew signal tristate
rlabel metal2 s 208122 163200 208178 164400 6 la_output[61]
port 537 nsew signal tristate
rlabel metal2 s 211434 163200 211490 164400 6 la_output[62]
port 538 nsew signal tristate
rlabel metal2 s 214838 163200 214894 164400 6 la_output[63]
port 539 nsew signal tristate
rlabel metal2 s 218242 163200 218298 164400 6 la_output[64]
port 540 nsew signal tristate
rlabel metal2 s 221554 163200 221610 164400 6 la_output[65]
port 541 nsew signal tristate
rlabel metal2 s 224958 163200 225014 164400 6 la_output[66]
port 542 nsew signal tristate
rlabel metal2 s 228270 163200 228326 164400 6 la_output[67]
port 543 nsew signal tristate
rlabel metal2 s 231674 163200 231730 164400 6 la_output[68]
port 544 nsew signal tristate
rlabel metal2 s 234986 163200 235042 164400 6 la_output[69]
port 545 nsew signal tristate
rlabel metal2 s 23018 163200 23074 164400 6 la_output[6]
port 546 nsew signal tristate
rlabel metal2 s 238390 163200 238446 164400 6 la_output[70]
port 547 nsew signal tristate
rlabel metal2 s 241794 163200 241850 164400 6 la_output[71]
port 548 nsew signal tristate
rlabel metal2 s 245106 163200 245162 164400 6 la_output[72]
port 549 nsew signal tristate
rlabel metal2 s 248510 163200 248566 164400 6 la_output[73]
port 550 nsew signal tristate
rlabel metal2 s 251822 163200 251878 164400 6 la_output[74]
port 551 nsew signal tristate
rlabel metal2 s 255226 163200 255282 164400 6 la_output[75]
port 552 nsew signal tristate
rlabel metal2 s 258538 163200 258594 164400 6 la_output[76]
port 553 nsew signal tristate
rlabel metal2 s 261942 163200 261998 164400 6 la_output[77]
port 554 nsew signal tristate
rlabel metal2 s 265346 163200 265402 164400 6 la_output[78]
port 555 nsew signal tristate
rlabel metal2 s 268658 163200 268714 164400 6 la_output[79]
port 556 nsew signal tristate
rlabel metal2 s 26422 163200 26478 164400 6 la_output[7]
port 557 nsew signal tristate
rlabel metal2 s 272062 163200 272118 164400 6 la_output[80]
port 558 nsew signal tristate
rlabel metal2 s 275374 163200 275430 164400 6 la_output[81]
port 559 nsew signal tristate
rlabel metal2 s 278778 163200 278834 164400 6 la_output[82]
port 560 nsew signal tristate
rlabel metal2 s 282090 163200 282146 164400 6 la_output[83]
port 561 nsew signal tristate
rlabel metal2 s 285494 163200 285550 164400 6 la_output[84]
port 562 nsew signal tristate
rlabel metal2 s 288898 163200 288954 164400 6 la_output[85]
port 563 nsew signal tristate
rlabel metal2 s 292210 163200 292266 164400 6 la_output[86]
port 564 nsew signal tristate
rlabel metal2 s 295614 163200 295670 164400 6 la_output[87]
port 565 nsew signal tristate
rlabel metal2 s 298926 163200 298982 164400 6 la_output[88]
port 566 nsew signal tristate
rlabel metal2 s 302330 163200 302386 164400 6 la_output[89]
port 567 nsew signal tristate
rlabel metal2 s 29826 163200 29882 164400 6 la_output[8]
port 568 nsew signal tristate
rlabel metal2 s 305642 163200 305698 164400 6 la_output[90]
port 569 nsew signal tristate
rlabel metal2 s 309046 163200 309102 164400 6 la_output[91]
port 570 nsew signal tristate
rlabel metal2 s 312450 163200 312506 164400 6 la_output[92]
port 571 nsew signal tristate
rlabel metal2 s 315762 163200 315818 164400 6 la_output[93]
port 572 nsew signal tristate
rlabel metal2 s 319166 163200 319222 164400 6 la_output[94]
port 573 nsew signal tristate
rlabel metal2 s 322478 163200 322534 164400 6 la_output[95]
port 574 nsew signal tristate
rlabel metal2 s 325882 163200 325938 164400 6 la_output[96]
port 575 nsew signal tristate
rlabel metal2 s 329194 163200 329250 164400 6 la_output[97]
port 576 nsew signal tristate
rlabel metal2 s 332598 163200 332654 164400 6 la_output[98]
port 577 nsew signal tristate
rlabel metal2 s 336002 163200 336058 164400 6 la_output[99]
port 578 nsew signal tristate
rlabel metal2 s 33138 163200 33194 164400 6 la_output[9]
port 579 nsew signal tristate
rlabel metal2 s 431038 163200 431094 164400 6 mprj_ack_i
port 580 nsew signal input
rlabel metal2 s 435178 163200 435234 164400 6 mprj_adr_o[0]
port 581 nsew signal tristate
rlabel metal2 s 463790 163200 463846 164400 6 mprj_adr_o[10]
port 582 nsew signal tristate
rlabel metal2 s 466366 163200 466422 164400 6 mprj_adr_o[11]
port 583 nsew signal tristate
rlabel metal2 s 468850 163200 468906 164400 6 mprj_adr_o[12]
port 584 nsew signal tristate
rlabel metal2 s 471426 163200 471482 164400 6 mprj_adr_o[13]
port 585 nsew signal tristate
rlabel metal2 s 473910 163200 473966 164400 6 mprj_adr_o[14]
port 586 nsew signal tristate
rlabel metal2 s 476394 163200 476450 164400 6 mprj_adr_o[15]
port 587 nsew signal tristate
rlabel metal2 s 478970 163200 479026 164400 6 mprj_adr_o[16]
port 588 nsew signal tristate
rlabel metal2 s 481454 163200 481510 164400 6 mprj_adr_o[17]
port 589 nsew signal tristate
rlabel metal2 s 484030 163200 484086 164400 6 mprj_adr_o[18]
port 590 nsew signal tristate
rlabel metal2 s 486514 163200 486570 164400 6 mprj_adr_o[19]
port 591 nsew signal tristate
rlabel metal2 s 438582 163200 438638 164400 6 mprj_adr_o[1]
port 592 nsew signal tristate
rlabel metal2 s 489090 163200 489146 164400 6 mprj_adr_o[20]
port 593 nsew signal tristate
rlabel metal2 s 491574 163200 491630 164400 6 mprj_adr_o[21]
port 594 nsew signal tristate
rlabel metal2 s 494058 163200 494114 164400 6 mprj_adr_o[22]
port 595 nsew signal tristate
rlabel metal2 s 496634 163200 496690 164400 6 mprj_adr_o[23]
port 596 nsew signal tristate
rlabel metal2 s 499118 163200 499174 164400 6 mprj_adr_o[24]
port 597 nsew signal tristate
rlabel metal2 s 501694 163200 501750 164400 6 mprj_adr_o[25]
port 598 nsew signal tristate
rlabel metal2 s 504178 163200 504234 164400 6 mprj_adr_o[26]
port 599 nsew signal tristate
rlabel metal2 s 506754 163200 506810 164400 6 mprj_adr_o[27]
port 600 nsew signal tristate
rlabel metal2 s 509238 163200 509294 164400 6 mprj_adr_o[28]
port 601 nsew signal tristate
rlabel metal2 s 511722 163200 511778 164400 6 mprj_adr_o[29]
port 602 nsew signal tristate
rlabel metal2 s 441986 163200 442042 164400 6 mprj_adr_o[2]
port 603 nsew signal tristate
rlabel metal2 s 514298 163200 514354 164400 6 mprj_adr_o[30]
port 604 nsew signal tristate
rlabel metal2 s 516782 163200 516838 164400 6 mprj_adr_o[31]
port 605 nsew signal tristate
rlabel metal2 s 445298 163200 445354 164400 6 mprj_adr_o[3]
port 606 nsew signal tristate
rlabel metal2 s 448702 163200 448758 164400 6 mprj_adr_o[4]
port 607 nsew signal tristate
rlabel metal2 s 451186 163200 451242 164400 6 mprj_adr_o[5]
port 608 nsew signal tristate
rlabel metal2 s 453762 163200 453818 164400 6 mprj_adr_o[6]
port 609 nsew signal tristate
rlabel metal2 s 456246 163200 456302 164400 6 mprj_adr_o[7]
port 610 nsew signal tristate
rlabel metal2 s 458730 163200 458786 164400 6 mprj_adr_o[8]
port 611 nsew signal tristate
rlabel metal2 s 461306 163200 461362 164400 6 mprj_adr_o[9]
port 612 nsew signal tristate
rlabel metal2 s 431866 163200 431922 164400 6 mprj_cyc_o
port 613 nsew signal tristate
rlabel metal2 s 436098 163200 436154 164400 6 mprj_dat_i[0]
port 614 nsew signal input
rlabel metal2 s 464618 163200 464674 164400 6 mprj_dat_i[10]
port 615 nsew signal input
rlabel metal2 s 467194 163200 467250 164400 6 mprj_dat_i[11]
port 616 nsew signal input
rlabel metal2 s 469678 163200 469734 164400 6 mprj_dat_i[12]
port 617 nsew signal input
rlabel metal2 s 472254 163200 472310 164400 6 mprj_dat_i[13]
port 618 nsew signal input
rlabel metal2 s 474738 163200 474794 164400 6 mprj_dat_i[14]
port 619 nsew signal input
rlabel metal2 s 477314 163200 477370 164400 6 mprj_dat_i[15]
port 620 nsew signal input
rlabel metal2 s 479798 163200 479854 164400 6 mprj_dat_i[16]
port 621 nsew signal input
rlabel metal2 s 482282 163200 482338 164400 6 mprj_dat_i[17]
port 622 nsew signal input
rlabel metal2 s 484858 163200 484914 164400 6 mprj_dat_i[18]
port 623 nsew signal input
rlabel metal2 s 487342 163200 487398 164400 6 mprj_dat_i[19]
port 624 nsew signal input
rlabel metal2 s 439410 163200 439466 164400 6 mprj_dat_i[1]
port 625 nsew signal input
rlabel metal2 s 489918 163200 489974 164400 6 mprj_dat_i[20]
port 626 nsew signal input
rlabel metal2 s 492402 163200 492458 164400 6 mprj_dat_i[21]
port 627 nsew signal input
rlabel metal2 s 494978 163200 495034 164400 6 mprj_dat_i[22]
port 628 nsew signal input
rlabel metal2 s 497462 163200 497518 164400 6 mprj_dat_i[23]
port 629 nsew signal input
rlabel metal2 s 499946 163200 500002 164400 6 mprj_dat_i[24]
port 630 nsew signal input
rlabel metal2 s 502522 163200 502578 164400 6 mprj_dat_i[25]
port 631 nsew signal input
rlabel metal2 s 505006 163200 505062 164400 6 mprj_dat_i[26]
port 632 nsew signal input
rlabel metal2 s 507582 163200 507638 164400 6 mprj_dat_i[27]
port 633 nsew signal input
rlabel metal2 s 510066 163200 510122 164400 6 mprj_dat_i[28]
port 634 nsew signal input
rlabel metal2 s 512642 163200 512698 164400 6 mprj_dat_i[29]
port 635 nsew signal input
rlabel metal2 s 442814 163200 442870 164400 6 mprj_dat_i[2]
port 636 nsew signal input
rlabel metal2 s 515126 163200 515182 164400 6 mprj_dat_i[30]
port 637 nsew signal input
rlabel metal2 s 517610 163200 517666 164400 6 mprj_dat_i[31]
port 638 nsew signal input
rlabel metal2 s 446126 163200 446182 164400 6 mprj_dat_i[3]
port 639 nsew signal input
rlabel metal2 s 449530 163200 449586 164400 6 mprj_dat_i[4]
port 640 nsew signal input
rlabel metal2 s 452014 163200 452070 164400 6 mprj_dat_i[5]
port 641 nsew signal input
rlabel metal2 s 454590 163200 454646 164400 6 mprj_dat_i[6]
port 642 nsew signal input
rlabel metal2 s 457074 163200 457130 164400 6 mprj_dat_i[7]
port 643 nsew signal input
rlabel metal2 s 459650 163200 459706 164400 6 mprj_dat_i[8]
port 644 nsew signal input
rlabel metal2 s 462134 163200 462190 164400 6 mprj_dat_i[9]
port 645 nsew signal input
rlabel metal2 s 436926 163200 436982 164400 6 mprj_dat_o[0]
port 646 nsew signal tristate
rlabel metal2 s 465538 163200 465594 164400 6 mprj_dat_o[10]
port 647 nsew signal tristate
rlabel metal2 s 468022 163200 468078 164400 6 mprj_dat_o[11]
port 648 nsew signal tristate
rlabel metal2 s 470506 163200 470562 164400 6 mprj_dat_o[12]
port 649 nsew signal tristate
rlabel metal2 s 473082 163200 473138 164400 6 mprj_dat_o[13]
port 650 nsew signal tristate
rlabel metal2 s 475566 163200 475622 164400 6 mprj_dat_o[14]
port 651 nsew signal tristate
rlabel metal2 s 478142 163200 478198 164400 6 mprj_dat_o[15]
port 652 nsew signal tristate
rlabel metal2 s 480626 163200 480682 164400 6 mprj_dat_o[16]
port 653 nsew signal tristate
rlabel metal2 s 483202 163200 483258 164400 6 mprj_dat_o[17]
port 654 nsew signal tristate
rlabel metal2 s 485686 163200 485742 164400 6 mprj_dat_o[18]
port 655 nsew signal tristate
rlabel metal2 s 488170 163200 488226 164400 6 mprj_dat_o[19]
port 656 nsew signal tristate
rlabel metal2 s 440238 163200 440294 164400 6 mprj_dat_o[1]
port 657 nsew signal tristate
rlabel metal2 s 490746 163200 490802 164400 6 mprj_dat_o[20]
port 658 nsew signal tristate
rlabel metal2 s 493230 163200 493286 164400 6 mprj_dat_o[21]
port 659 nsew signal tristate
rlabel metal2 s 495806 163200 495862 164400 6 mprj_dat_o[22]
port 660 nsew signal tristate
rlabel metal2 s 498290 163200 498346 164400 6 mprj_dat_o[23]
port 661 nsew signal tristate
rlabel metal2 s 500866 163200 500922 164400 6 mprj_dat_o[24]
port 662 nsew signal tristate
rlabel metal2 s 503350 163200 503406 164400 6 mprj_dat_o[25]
port 663 nsew signal tristate
rlabel metal2 s 505834 163200 505890 164400 6 mprj_dat_o[26]
port 664 nsew signal tristate
rlabel metal2 s 508410 163200 508466 164400 6 mprj_dat_o[27]
port 665 nsew signal tristate
rlabel metal2 s 510894 163200 510950 164400 6 mprj_dat_o[28]
port 666 nsew signal tristate
rlabel metal2 s 513470 163200 513526 164400 6 mprj_dat_o[29]
port 667 nsew signal tristate
rlabel metal2 s 443642 163200 443698 164400 6 mprj_dat_o[2]
port 668 nsew signal tristate
rlabel metal2 s 515954 163200 516010 164400 6 mprj_dat_o[30]
port 669 nsew signal tristate
rlabel metal2 s 518530 163200 518586 164400 6 mprj_dat_o[31]
port 670 nsew signal tristate
rlabel metal2 s 446954 163200 447010 164400 6 mprj_dat_o[3]
port 671 nsew signal tristate
rlabel metal2 s 450358 163200 450414 164400 6 mprj_dat_o[4]
port 672 nsew signal tristate
rlabel metal2 s 452842 163200 452898 164400 6 mprj_dat_o[5]
port 673 nsew signal tristate
rlabel metal2 s 455418 163200 455474 164400 6 mprj_dat_o[6]
port 674 nsew signal tristate
rlabel metal2 s 457902 163200 457958 164400 6 mprj_dat_o[7]
port 675 nsew signal tristate
rlabel metal2 s 460478 163200 460534 164400 6 mprj_dat_o[8]
port 676 nsew signal tristate
rlabel metal2 s 462962 163200 463018 164400 6 mprj_dat_o[9]
port 677 nsew signal tristate
rlabel metal2 s 437754 163200 437810 164400 6 mprj_sel_o[0]
port 678 nsew signal tristate
rlabel metal2 s 441066 163200 441122 164400 6 mprj_sel_o[1]
port 679 nsew signal tristate
rlabel metal2 s 444470 163200 444526 164400 6 mprj_sel_o[2]
port 680 nsew signal tristate
rlabel metal2 s 447874 163200 447930 164400 6 mprj_sel_o[3]
port 681 nsew signal tristate
rlabel metal2 s 432694 163200 432750 164400 6 mprj_stb_o
port 682 nsew signal tristate
rlabel metal2 s 433522 163200 433578 164400 6 mprj_wb_iena
port 683 nsew signal tristate
rlabel metal2 s 434350 163200 434406 164400 6 mprj_we_o
port 684 nsew signal tristate
rlabel metal3 s 523200 90176 524400 90296 6 qspi_enabled
port 685 nsew signal tristate
rlabel metal3 s 523200 84192 524400 84312 6 ser_rx
port 686 nsew signal input
rlabel metal3 s 523200 85688 524400 85808 6 ser_tx
port 687 nsew signal tristate
rlabel metal3 s 523200 81064 524400 81184 6 spi_csb
port 688 nsew signal tristate
rlabel metal3 s 523200 87184 524400 87304 6 spi_enabled
port 689 nsew signal tristate
rlabel metal3 s 523200 79568 524400 79688 6 spi_sck
port 690 nsew signal tristate
rlabel metal3 s 523200 82696 524400 82816 6 spi_sdi
port 691 nsew signal input
rlabel metal3 s 523200 78072 524400 78192 6 spi_sdo
port 692 nsew signal tristate
rlabel metal3 s 523200 76576 524400 76696 6 spi_sdoenb
port 693 nsew signal tristate
rlabel metal3 s 523200 2184 524400 2304 6 sram_ro_addr[0]
port 694 nsew signal input
rlabel metal3 s 523200 3680 524400 3800 6 sram_ro_addr[1]
port 695 nsew signal input
rlabel metal3 s 523200 5176 524400 5296 6 sram_ro_addr[2]
port 696 nsew signal input
rlabel metal3 s 523200 6672 524400 6792 6 sram_ro_addr[3]
port 697 nsew signal input
rlabel metal3 s 523200 8168 524400 8288 6 sram_ro_addr[4]
port 698 nsew signal input
rlabel metal3 s 523200 9800 524400 9920 6 sram_ro_addr[5]
port 699 nsew signal input
rlabel metal3 s 523200 11296 524400 11416 6 sram_ro_addr[6]
port 700 nsew signal input
rlabel metal3 s 523200 12792 524400 12912 6 sram_ro_addr[7]
port 701 nsew signal input
rlabel metal3 s 523200 14288 524400 14408 6 sram_ro_clk
port 702 nsew signal input
rlabel metal3 s 523200 688 524400 808 6 sram_ro_csb
port 703 nsew signal input
rlabel metal3 s 523200 15784 524400 15904 6 sram_ro_data[0]
port 704 nsew signal tristate
rlabel metal3 s 523200 31016 524400 31136 6 sram_ro_data[10]
port 705 nsew signal tristate
rlabel metal3 s 523200 32512 524400 32632 6 sram_ro_data[11]
port 706 nsew signal tristate
rlabel metal3 s 523200 34008 524400 34128 6 sram_ro_data[12]
port 707 nsew signal tristate
rlabel metal3 s 523200 35504 524400 35624 6 sram_ro_data[13]
port 708 nsew signal tristate
rlabel metal3 s 523200 37136 524400 37256 6 sram_ro_data[14]
port 709 nsew signal tristate
rlabel metal3 s 523200 38632 524400 38752 6 sram_ro_data[15]
port 710 nsew signal tristate
rlabel metal3 s 523200 40128 524400 40248 6 sram_ro_data[16]
port 711 nsew signal tristate
rlabel metal3 s 523200 41624 524400 41744 6 sram_ro_data[17]
port 712 nsew signal tristate
rlabel metal3 s 523200 43120 524400 43240 6 sram_ro_data[18]
port 713 nsew signal tristate
rlabel metal3 s 523200 44616 524400 44736 6 sram_ro_data[19]
port 714 nsew signal tristate
rlabel metal3 s 523200 17280 524400 17400 6 sram_ro_data[1]
port 715 nsew signal tristate
rlabel metal3 s 523200 46248 524400 46368 6 sram_ro_data[20]
port 716 nsew signal tristate
rlabel metal3 s 523200 47744 524400 47864 6 sram_ro_data[21]
port 717 nsew signal tristate
rlabel metal3 s 523200 49240 524400 49360 6 sram_ro_data[22]
port 718 nsew signal tristate
rlabel metal3 s 523200 50736 524400 50856 6 sram_ro_data[23]
port 719 nsew signal tristate
rlabel metal3 s 523200 52232 524400 52352 6 sram_ro_data[24]
port 720 nsew signal tristate
rlabel metal3 s 523200 53728 524400 53848 6 sram_ro_data[25]
port 721 nsew signal tristate
rlabel metal3 s 523200 55360 524400 55480 6 sram_ro_data[26]
port 722 nsew signal tristate
rlabel metal3 s 523200 56856 524400 56976 6 sram_ro_data[27]
port 723 nsew signal tristate
rlabel metal3 s 523200 58352 524400 58472 6 sram_ro_data[28]
port 724 nsew signal tristate
rlabel metal3 s 523200 59848 524400 59968 6 sram_ro_data[29]
port 725 nsew signal tristate
rlabel metal3 s 523200 18912 524400 19032 6 sram_ro_data[2]
port 726 nsew signal tristate
rlabel metal3 s 523200 61344 524400 61464 6 sram_ro_data[30]
port 727 nsew signal tristate
rlabel metal3 s 523200 62840 524400 62960 6 sram_ro_data[31]
port 728 nsew signal tristate
rlabel metal3 s 523200 20408 524400 20528 6 sram_ro_data[3]
port 729 nsew signal tristate
rlabel metal3 s 523200 21904 524400 22024 6 sram_ro_data[4]
port 730 nsew signal tristate
rlabel metal3 s 523200 23400 524400 23520 6 sram_ro_data[5]
port 731 nsew signal tristate
rlabel metal3 s 523200 24896 524400 25016 6 sram_ro_data[6]
port 732 nsew signal tristate
rlabel metal3 s 523200 26392 524400 26512 6 sram_ro_data[7]
port 733 nsew signal tristate
rlabel metal3 s 523200 28024 524400 28144 6 sram_ro_data[8]
port 734 nsew signal tristate
rlabel metal3 s 523200 29520 524400 29640 6 sram_ro_data[9]
port 735 nsew signal tristate
rlabel metal3 s 523200 70456 524400 70576 6 trap
port 736 nsew signal tristate
rlabel metal3 s 523200 88680 524400 88800 6 uart_enabled
port 737 nsew signal tristate
rlabel metal2 s 519358 163200 519414 164400 6 user_irq_ena[0]
port 738 nsew signal tristate
rlabel metal2 s 520186 163200 520242 164400 6 user_irq_ena[1]
port 739 nsew signal tristate
rlabel metal2 s 521014 163200 521070 164400 6 user_irq_ena[2]
port 740 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 524000 164000
<< end >>
