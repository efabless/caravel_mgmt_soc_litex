magic
tech sky130A
magscale 1 2
timestamp 1675791412
<< obsli1 >>
rect 552 527 79948 93585
<< obsm1 >>
rect 198 76 80486 94104
<< metal2 >>
rect 1674 93712 1730 94112
rect 4158 93712 4214 94112
rect 6642 93712 6698 94112
rect 9126 93712 9182 94112
rect 11610 93712 11666 94112
rect 14094 93712 14150 94112
rect 16578 93712 16634 94112
rect 19062 93712 19118 94112
rect 21546 93712 21602 94112
rect 24030 93712 24086 94112
rect 26514 93712 26570 94112
rect 28998 93712 29054 94112
rect 31482 93712 31538 94112
rect 33966 93712 34022 94112
rect 36450 93712 36506 94112
rect 38934 93712 38990 94112
rect 41418 93712 41474 94112
rect 43902 93712 43958 94112
rect 46386 93712 46442 94112
rect 48870 93712 48926 94112
rect 51354 93712 51410 94112
rect 53838 93712 53894 94112
rect 56322 93712 56378 94112
rect 58806 93712 58862 94112
rect 61290 93712 61346 94112
rect 63774 93712 63830 94112
rect 66258 93712 66314 94112
rect 68742 93712 68798 94112
rect 71226 93712 71282 94112
rect 73710 93712 73766 94112
rect 76194 93712 76250 94112
rect 78678 93712 78734 94112
rect 1674 0 1730 400
rect 4158 0 4214 400
rect 6642 0 6698 400
rect 9126 0 9182 400
rect 11610 0 11666 400
rect 14094 0 14150 400
rect 16578 0 16634 400
rect 19062 0 19118 400
rect 21546 0 21602 400
rect 24030 0 24086 400
rect 26514 0 26570 400
rect 28998 0 29054 400
rect 31482 0 31538 400
rect 33966 0 34022 400
rect 36450 0 36506 400
rect 38934 0 38990 400
rect 41418 0 41474 400
rect 43902 0 43958 400
rect 46386 0 46442 400
rect 48870 0 48926 400
rect 51354 0 51410 400
rect 53838 0 53894 400
rect 56322 0 56378 400
rect 58806 0 58862 400
rect 61290 0 61346 400
rect 63774 0 63830 400
rect 66258 0 66314 400
rect 68742 0 68798 400
rect 71226 0 71282 400
rect 73710 0 73766 400
rect 76194 0 76250 400
rect 78678 0 78734 400
<< obsm2 >>
rect 204 93656 1618 94110
rect 1786 93656 4102 94110
rect 4270 93656 6586 94110
rect 6754 93656 9070 94110
rect 9238 93656 11554 94110
rect 11722 93656 14038 94110
rect 14206 93656 16522 94110
rect 16690 93656 19006 94110
rect 19174 93656 21490 94110
rect 21658 93656 23974 94110
rect 24142 93656 26458 94110
rect 26626 93656 28942 94110
rect 29110 93656 31426 94110
rect 31594 93656 33910 94110
rect 34078 93656 36394 94110
rect 36562 93656 38878 94110
rect 39046 93656 41362 94110
rect 41530 93656 43846 94110
rect 44014 93656 46330 94110
rect 46498 93656 48814 94110
rect 48982 93656 51298 94110
rect 51466 93656 53782 94110
rect 53950 93656 56266 94110
rect 56434 93656 58750 94110
rect 58918 93656 61234 94110
rect 61402 93656 63718 94110
rect 63886 93656 66202 94110
rect 66370 93656 68686 94110
rect 68854 93656 71170 94110
rect 71338 93656 73654 94110
rect 73822 93656 76138 94110
rect 76306 93656 78622 94110
rect 78790 93656 80480 94110
rect 204 456 80480 93656
rect 204 70 1618 456
rect 1786 70 4102 456
rect 4270 70 6586 456
rect 6754 70 9070 456
rect 9238 70 11554 456
rect 11722 70 14038 456
rect 14206 70 16522 456
rect 16690 70 19006 456
rect 19174 70 21490 456
rect 21658 70 23974 456
rect 24142 70 26458 456
rect 26626 70 28942 456
rect 29110 70 31426 456
rect 31594 70 33910 456
rect 34078 70 36394 456
rect 36562 70 38878 456
rect 39046 70 41362 456
rect 41530 70 43846 456
rect 44014 70 46330 456
rect 46498 70 48814 456
rect 48982 70 51298 456
rect 51466 70 53782 456
rect 53950 70 56266 456
rect 56434 70 58750 456
rect 58918 70 61234 456
rect 61402 70 63718 456
rect 63886 70 66202 456
rect 66370 70 68686 456
rect 68854 70 71170 456
rect 71338 70 73654 456
rect 73822 70 76138 456
rect 76306 70 78622 456
rect 78790 70 80480 456
<< metal3 >>
rect 80100 89632 80500 89752
rect 80100 81880 80500 82000
rect 80100 74128 80500 74248
rect 80100 66376 80500 66496
rect 80100 58624 80500 58744
rect 80100 50872 80500 50992
rect 0 46928 400 47048
rect 80100 43120 80500 43240
rect 80100 35368 80500 35488
rect 80100 27616 80500 27736
rect 80100 19864 80500 19984
rect 80100 12112 80500 12232
rect 80100 4360 80500 4480
<< obsm3 >>
rect 400 89832 80395 94108
rect 400 89552 80020 89832
rect 400 82080 80395 89552
rect 400 81800 80020 82080
rect 400 74328 80395 81800
rect 400 74048 80020 74328
rect 400 66576 80395 74048
rect 400 66296 80020 66576
rect 400 58824 80395 66296
rect 400 58544 80020 58824
rect 400 51072 80395 58544
rect 400 50792 80020 51072
rect 400 47128 80395 50792
rect 480 46848 80395 47128
rect 400 43320 80395 46848
rect 400 43040 80020 43320
rect 400 35568 80395 43040
rect 400 35288 80020 35568
rect 400 27816 80395 35288
rect 400 27536 80020 27816
rect 400 20064 80395 27536
rect 400 19784 80020 20064
rect 400 12312 80395 19784
rect 400 12032 80020 12312
rect 400 4560 80395 12032
rect 400 4280 80020 4560
rect 400 171 80395 4280
<< metal4 >>
rect 3656 496 3976 93616
rect 19016 496 19336 93616
rect 34376 496 34696 93616
rect 49736 496 50056 93616
rect 65096 496 65416 93616
<< obsm4 >>
rect 2267 93696 78877 94077
rect 2267 3435 3576 93696
rect 4056 3435 18936 93696
rect 19416 3435 34296 93696
rect 34776 3435 49656 93696
rect 50136 3435 65016 93696
rect 65496 3435 78877 93696
<< labels >>
rlabel metal3 s 80100 43120 80500 43240 6 A0[0]
port 1 nsew signal input
rlabel metal3 s 80100 50872 80500 50992 6 A0[1]
port 2 nsew signal input
rlabel metal3 s 80100 58624 80500 58744 6 A0[2]
port 3 nsew signal input
rlabel metal3 s 80100 66376 80500 66496 6 A0[3]
port 4 nsew signal input
rlabel metal3 s 80100 74128 80500 74248 6 A0[4]
port 5 nsew signal input
rlabel metal3 s 80100 81880 80500 82000 6 A0[5]
port 6 nsew signal input
rlabel metal3 s 80100 89632 80500 89752 6 A0[6]
port 7 nsew signal input
rlabel metal3 s 0 46928 400 47048 6 CLK
port 8 nsew signal input
rlabel metal2 s 1674 0 1730 400 6 Di0[0]
port 9 nsew signal input
rlabel metal2 s 26514 0 26570 400 6 Di0[10]
port 10 nsew signal input
rlabel metal2 s 28998 0 29054 400 6 Di0[11]
port 11 nsew signal input
rlabel metal2 s 31482 0 31538 400 6 Di0[12]
port 12 nsew signal input
rlabel metal2 s 33966 0 34022 400 6 Di0[13]
port 13 nsew signal input
rlabel metal2 s 36450 0 36506 400 6 Di0[14]
port 14 nsew signal input
rlabel metal2 s 38934 0 38990 400 6 Di0[15]
port 15 nsew signal input
rlabel metal2 s 41418 0 41474 400 6 Di0[16]
port 16 nsew signal input
rlabel metal2 s 43902 0 43958 400 6 Di0[17]
port 17 nsew signal input
rlabel metal2 s 46386 0 46442 400 6 Di0[18]
port 18 nsew signal input
rlabel metal2 s 48870 0 48926 400 6 Di0[19]
port 19 nsew signal input
rlabel metal2 s 4158 0 4214 400 6 Di0[1]
port 20 nsew signal input
rlabel metal2 s 51354 0 51410 400 6 Di0[20]
port 21 nsew signal input
rlabel metal2 s 53838 0 53894 400 6 Di0[21]
port 22 nsew signal input
rlabel metal2 s 56322 0 56378 400 6 Di0[22]
port 23 nsew signal input
rlabel metal2 s 58806 0 58862 400 6 Di0[23]
port 24 nsew signal input
rlabel metal2 s 61290 0 61346 400 6 Di0[24]
port 25 nsew signal input
rlabel metal2 s 63774 0 63830 400 6 Di0[25]
port 26 nsew signal input
rlabel metal2 s 66258 0 66314 400 6 Di0[26]
port 27 nsew signal input
rlabel metal2 s 68742 0 68798 400 6 Di0[27]
port 28 nsew signal input
rlabel metal2 s 71226 0 71282 400 6 Di0[28]
port 29 nsew signal input
rlabel metal2 s 73710 0 73766 400 6 Di0[29]
port 30 nsew signal input
rlabel metal2 s 6642 0 6698 400 6 Di0[2]
port 31 nsew signal input
rlabel metal2 s 76194 0 76250 400 6 Di0[30]
port 32 nsew signal input
rlabel metal2 s 78678 0 78734 400 6 Di0[31]
port 33 nsew signal input
rlabel metal2 s 9126 0 9182 400 6 Di0[3]
port 34 nsew signal input
rlabel metal2 s 11610 0 11666 400 6 Di0[4]
port 35 nsew signal input
rlabel metal2 s 14094 0 14150 400 6 Di0[5]
port 36 nsew signal input
rlabel metal2 s 16578 0 16634 400 6 Di0[6]
port 37 nsew signal input
rlabel metal2 s 19062 0 19118 400 6 Di0[7]
port 38 nsew signal input
rlabel metal2 s 21546 0 21602 400 6 Di0[8]
port 39 nsew signal input
rlabel metal2 s 24030 0 24086 400 6 Di0[9]
port 40 nsew signal input
rlabel metal2 s 1674 93712 1730 94112 6 Do0[0]
port 41 nsew signal output
rlabel metal2 s 26514 93712 26570 94112 6 Do0[10]
port 42 nsew signal output
rlabel metal2 s 28998 93712 29054 94112 6 Do0[11]
port 43 nsew signal output
rlabel metal2 s 31482 93712 31538 94112 6 Do0[12]
port 44 nsew signal output
rlabel metal2 s 33966 93712 34022 94112 6 Do0[13]
port 45 nsew signal output
rlabel metal2 s 36450 93712 36506 94112 6 Do0[14]
port 46 nsew signal output
rlabel metal2 s 38934 93712 38990 94112 6 Do0[15]
port 47 nsew signal output
rlabel metal2 s 41418 93712 41474 94112 6 Do0[16]
port 48 nsew signal output
rlabel metal2 s 43902 93712 43958 94112 6 Do0[17]
port 49 nsew signal output
rlabel metal2 s 46386 93712 46442 94112 6 Do0[18]
port 50 nsew signal output
rlabel metal2 s 48870 93712 48926 94112 6 Do0[19]
port 51 nsew signal output
rlabel metal2 s 4158 93712 4214 94112 6 Do0[1]
port 52 nsew signal output
rlabel metal2 s 51354 93712 51410 94112 6 Do0[20]
port 53 nsew signal output
rlabel metal2 s 53838 93712 53894 94112 6 Do0[21]
port 54 nsew signal output
rlabel metal2 s 56322 93712 56378 94112 6 Do0[22]
port 55 nsew signal output
rlabel metal2 s 58806 93712 58862 94112 6 Do0[23]
port 56 nsew signal output
rlabel metal2 s 61290 93712 61346 94112 6 Do0[24]
port 57 nsew signal output
rlabel metal2 s 63774 93712 63830 94112 6 Do0[25]
port 58 nsew signal output
rlabel metal2 s 66258 93712 66314 94112 6 Do0[26]
port 59 nsew signal output
rlabel metal2 s 68742 93712 68798 94112 6 Do0[27]
port 60 nsew signal output
rlabel metal2 s 71226 93712 71282 94112 6 Do0[28]
port 61 nsew signal output
rlabel metal2 s 73710 93712 73766 94112 6 Do0[29]
port 62 nsew signal output
rlabel metal2 s 6642 93712 6698 94112 6 Do0[2]
port 63 nsew signal output
rlabel metal2 s 76194 93712 76250 94112 6 Do0[30]
port 64 nsew signal output
rlabel metal2 s 78678 93712 78734 94112 6 Do0[31]
port 65 nsew signal output
rlabel metal2 s 9126 93712 9182 94112 6 Do0[3]
port 66 nsew signal output
rlabel metal2 s 11610 93712 11666 94112 6 Do0[4]
port 67 nsew signal output
rlabel metal2 s 14094 93712 14150 94112 6 Do0[5]
port 68 nsew signal output
rlabel metal2 s 16578 93712 16634 94112 6 Do0[6]
port 69 nsew signal output
rlabel metal2 s 19062 93712 19118 94112 6 Do0[7]
port 70 nsew signal output
rlabel metal2 s 21546 93712 21602 94112 6 Do0[8]
port 71 nsew signal output
rlabel metal2 s 24030 93712 24086 94112 6 Do0[9]
port 72 nsew signal output
rlabel metal3 s 80100 4360 80500 4480 6 EN0
port 73 nsew signal input
rlabel metal4 s 19016 496 19336 93616 6 VGND
port 74 nsew ground bidirectional
rlabel metal4 s 49736 496 50056 93616 6 VGND
port 74 nsew ground bidirectional
rlabel metal4 s 3656 496 3976 93616 6 VPWR
port 75 nsew power bidirectional
rlabel metal4 s 34376 496 34696 93616 6 VPWR
port 75 nsew power bidirectional
rlabel metal4 s 65096 496 65416 93616 6 VPWR
port 75 nsew power bidirectional
rlabel metal3 s 80100 12112 80500 12232 6 WE0[0]
port 76 nsew signal input
rlabel metal3 s 80100 19864 80500 19984 6 WE0[1]
port 77 nsew signal input
rlabel metal3 s 80100 27616 80500 27736 6 WE0[2]
port 78 nsew signal input
rlabel metal3 s 80100 35368 80500 35488 6 WE0[3]
port 79 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 80500 94112
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 24017876
string GDS_FILE /mnt/dffram/build/128x32_DEFAULT/openlane/runs/RUN_2023.02.07_17.13.21/results/signoff/RAM128.magic.gds
string GDS_START 183640
<< end >>

