magic
tech sky130A
magscale 1 2
timestamp 1639080793
<< obsli1 >>
rect 2869 4159 516900 147809
<< obsm1 >>
rect 382 756 523558 160064
<< metal2 >>
rect 386 163200 442 164400
rect 1214 163200 1270 164400
rect 2042 163200 2098 164400
rect 2870 163200 2926 164400
rect 3698 163200 3754 164400
rect 4526 163200 4582 164400
rect 5354 163200 5410 164400
rect 6274 163200 6330 164400
rect 7102 163200 7158 164400
rect 7930 163200 7986 164400
rect 8758 163200 8814 164400
rect 9586 163200 9642 164400
rect 10414 163200 10470 164400
rect 11242 163200 11298 164400
rect 12162 163200 12218 164400
rect 12990 163200 13046 164400
rect 13818 163200 13874 164400
rect 14646 163200 14702 164400
rect 15474 163200 15530 164400
rect 16302 163200 16358 164400
rect 17130 163200 17186 164400
rect 18050 163200 18106 164400
rect 18878 163200 18934 164400
rect 19706 163200 19762 164400
rect 20534 163200 20590 164400
rect 21362 163200 21418 164400
rect 22190 163200 22246 164400
rect 23018 163200 23074 164400
rect 23938 163200 23994 164400
rect 24766 163200 24822 164400
rect 25594 163200 25650 164400
rect 26422 163200 26478 164400
rect 27250 163200 27306 164400
rect 28078 163200 28134 164400
rect 28906 163200 28962 164400
rect 29826 163200 29882 164400
rect 30654 163200 30710 164400
rect 31482 163200 31538 164400
rect 32310 163200 32366 164400
rect 33138 163200 33194 164400
rect 33966 163200 34022 164400
rect 34794 163200 34850 164400
rect 35714 163200 35770 164400
rect 36542 163200 36598 164400
rect 37370 163200 37426 164400
rect 38198 163200 38254 164400
rect 39026 163200 39082 164400
rect 39854 163200 39910 164400
rect 40682 163200 40738 164400
rect 41602 163200 41658 164400
rect 42430 163200 42486 164400
rect 43258 163200 43314 164400
rect 44086 163200 44142 164400
rect 44914 163200 44970 164400
rect 45742 163200 45798 164400
rect 46570 163200 46626 164400
rect 47490 163200 47546 164400
rect 48318 163200 48374 164400
rect 49146 163200 49202 164400
rect 49974 163200 50030 164400
rect 50802 163200 50858 164400
rect 51630 163200 51686 164400
rect 52458 163200 52514 164400
rect 53378 163200 53434 164400
rect 54206 163200 54262 164400
rect 55034 163200 55090 164400
rect 55862 163200 55918 164400
rect 56690 163200 56746 164400
rect 57518 163200 57574 164400
rect 58346 163200 58402 164400
rect 59266 163200 59322 164400
rect 60094 163200 60150 164400
rect 60922 163200 60978 164400
rect 61750 163200 61806 164400
rect 62578 163200 62634 164400
rect 63406 163200 63462 164400
rect 64234 163200 64290 164400
rect 65154 163200 65210 164400
rect 65982 163200 66038 164400
rect 66810 163200 66866 164400
rect 67638 163200 67694 164400
rect 68466 163200 68522 164400
rect 69294 163200 69350 164400
rect 70122 163200 70178 164400
rect 71042 163200 71098 164400
rect 71870 163200 71926 164400
rect 72698 163200 72754 164400
rect 73526 163200 73582 164400
rect 74354 163200 74410 164400
rect 75182 163200 75238 164400
rect 76010 163200 76066 164400
rect 76930 163200 76986 164400
rect 77758 163200 77814 164400
rect 78586 163200 78642 164400
rect 79414 163200 79470 164400
rect 80242 163200 80298 164400
rect 81070 163200 81126 164400
rect 81898 163200 81954 164400
rect 82818 163200 82874 164400
rect 83646 163200 83702 164400
rect 84474 163200 84530 164400
rect 85302 163200 85358 164400
rect 86130 163200 86186 164400
rect 86958 163200 87014 164400
rect 87786 163200 87842 164400
rect 88706 163200 88762 164400
rect 89534 163200 89590 164400
rect 90362 163200 90418 164400
rect 91190 163200 91246 164400
rect 92018 163200 92074 164400
rect 92846 163200 92902 164400
rect 93674 163200 93730 164400
rect 94594 163200 94650 164400
rect 95422 163200 95478 164400
rect 96250 163200 96306 164400
rect 97078 163200 97134 164400
rect 97906 163200 97962 164400
rect 98734 163200 98790 164400
rect 99562 163200 99618 164400
rect 100482 163200 100538 164400
rect 101310 163200 101366 164400
rect 102138 163200 102194 164400
rect 102966 163200 103022 164400
rect 103794 163200 103850 164400
rect 104622 163200 104678 164400
rect 105450 163200 105506 164400
rect 106370 163200 106426 164400
rect 107198 163200 107254 164400
rect 108026 163200 108082 164400
rect 108854 163200 108910 164400
rect 109682 163200 109738 164400
rect 110510 163200 110566 164400
rect 111338 163200 111394 164400
rect 112258 163200 112314 164400
rect 113086 163200 113142 164400
rect 113914 163200 113970 164400
rect 114742 163200 114798 164400
rect 115570 163200 115626 164400
rect 116398 163200 116454 164400
rect 117226 163200 117282 164400
rect 118146 163200 118202 164400
rect 118974 163200 119030 164400
rect 119802 163200 119858 164400
rect 120630 163200 120686 164400
rect 121458 163200 121514 164400
rect 122286 163200 122342 164400
rect 123114 163200 123170 164400
rect 124034 163200 124090 164400
rect 124862 163200 124918 164400
rect 125690 163200 125746 164400
rect 126518 163200 126574 164400
rect 127346 163200 127402 164400
rect 128174 163200 128230 164400
rect 129002 163200 129058 164400
rect 129922 163200 129978 164400
rect 130750 163200 130806 164400
rect 131578 163200 131634 164400
rect 132406 163200 132462 164400
rect 133234 163200 133290 164400
rect 134062 163200 134118 164400
rect 134890 163200 134946 164400
rect 135810 163200 135866 164400
rect 136638 163200 136694 164400
rect 137466 163200 137522 164400
rect 138294 163200 138350 164400
rect 139122 163200 139178 164400
rect 139950 163200 140006 164400
rect 140778 163200 140834 164400
rect 141698 163200 141754 164400
rect 142526 163200 142582 164400
rect 143354 163200 143410 164400
rect 144182 163200 144238 164400
rect 145010 163200 145066 164400
rect 145838 163200 145894 164400
rect 146666 163200 146722 164400
rect 147586 163200 147642 164400
rect 148414 163200 148470 164400
rect 149242 163200 149298 164400
rect 150070 163200 150126 164400
rect 150898 163200 150954 164400
rect 151726 163200 151782 164400
rect 152554 163200 152610 164400
rect 153474 163200 153530 164400
rect 154302 163200 154358 164400
rect 155130 163200 155186 164400
rect 155958 163200 156014 164400
rect 156786 163200 156842 164400
rect 157614 163200 157670 164400
rect 158442 163200 158498 164400
rect 159362 163200 159418 164400
rect 160190 163200 160246 164400
rect 161018 163200 161074 164400
rect 161846 163200 161902 164400
rect 162674 163200 162730 164400
rect 163502 163200 163558 164400
rect 164330 163200 164386 164400
rect 165250 163200 165306 164400
rect 166078 163200 166134 164400
rect 166906 163200 166962 164400
rect 167734 163200 167790 164400
rect 168562 163200 168618 164400
rect 169390 163200 169446 164400
rect 170218 163200 170274 164400
rect 171138 163200 171194 164400
rect 171966 163200 172022 164400
rect 172794 163200 172850 164400
rect 173622 163200 173678 164400
rect 174450 163200 174506 164400
rect 175278 163200 175334 164400
rect 176106 163200 176162 164400
rect 177026 163200 177082 164400
rect 177854 163200 177910 164400
rect 178682 163200 178738 164400
rect 179510 163200 179566 164400
rect 180338 163200 180394 164400
rect 181166 163200 181222 164400
rect 181994 163200 182050 164400
rect 182914 163200 182970 164400
rect 183742 163200 183798 164400
rect 184570 163200 184626 164400
rect 185398 163200 185454 164400
rect 186226 163200 186282 164400
rect 187054 163200 187110 164400
rect 187882 163200 187938 164400
rect 188802 163200 188858 164400
rect 189630 163200 189686 164400
rect 190458 163200 190514 164400
rect 191286 163200 191342 164400
rect 192114 163200 192170 164400
rect 192942 163200 192998 164400
rect 193770 163200 193826 164400
rect 194690 163200 194746 164400
rect 195518 163200 195574 164400
rect 196346 163200 196402 164400
rect 197174 163200 197230 164400
rect 198002 163200 198058 164400
rect 198830 163200 198886 164400
rect 199658 163200 199714 164400
rect 200578 163200 200634 164400
rect 201406 163200 201462 164400
rect 202234 163200 202290 164400
rect 203062 163200 203118 164400
rect 203890 163200 203946 164400
rect 204718 163200 204774 164400
rect 205546 163200 205602 164400
rect 206466 163200 206522 164400
rect 207294 163200 207350 164400
rect 208122 163200 208178 164400
rect 208950 163200 209006 164400
rect 209778 163200 209834 164400
rect 210606 163200 210662 164400
rect 211434 163200 211490 164400
rect 212354 163200 212410 164400
rect 213182 163200 213238 164400
rect 214010 163200 214066 164400
rect 214838 163200 214894 164400
rect 215666 163200 215722 164400
rect 216494 163200 216550 164400
rect 217322 163200 217378 164400
rect 218242 163200 218298 164400
rect 219070 163200 219126 164400
rect 219898 163200 219954 164400
rect 220726 163200 220782 164400
rect 221554 163200 221610 164400
rect 222382 163200 222438 164400
rect 223210 163200 223266 164400
rect 224130 163200 224186 164400
rect 224958 163200 225014 164400
rect 225786 163200 225842 164400
rect 226614 163200 226670 164400
rect 227442 163200 227498 164400
rect 228270 163200 228326 164400
rect 229098 163200 229154 164400
rect 230018 163200 230074 164400
rect 230846 163200 230902 164400
rect 231674 163200 231730 164400
rect 232502 163200 232558 164400
rect 233330 163200 233386 164400
rect 234158 163200 234214 164400
rect 234986 163200 235042 164400
rect 235906 163200 235962 164400
rect 236734 163200 236790 164400
rect 237562 163200 237618 164400
rect 238390 163200 238446 164400
rect 239218 163200 239274 164400
rect 240046 163200 240102 164400
rect 240874 163200 240930 164400
rect 241794 163200 241850 164400
rect 242622 163200 242678 164400
rect 243450 163200 243506 164400
rect 244278 163200 244334 164400
rect 245106 163200 245162 164400
rect 245934 163200 245990 164400
rect 246762 163200 246818 164400
rect 247682 163200 247738 164400
rect 248510 163200 248566 164400
rect 249338 163200 249394 164400
rect 250166 163200 250222 164400
rect 250994 163200 251050 164400
rect 251822 163200 251878 164400
rect 252650 163200 252706 164400
rect 253570 163200 253626 164400
rect 254398 163200 254454 164400
rect 255226 163200 255282 164400
rect 256054 163200 256110 164400
rect 256882 163200 256938 164400
rect 257710 163200 257766 164400
rect 258538 163200 258594 164400
rect 259458 163200 259514 164400
rect 260286 163200 260342 164400
rect 261114 163200 261170 164400
rect 261942 163200 261998 164400
rect 262770 163200 262826 164400
rect 263598 163200 263654 164400
rect 264426 163200 264482 164400
rect 265346 163200 265402 164400
rect 266174 163200 266230 164400
rect 267002 163200 267058 164400
rect 267830 163200 267886 164400
rect 268658 163200 268714 164400
rect 269486 163200 269542 164400
rect 270314 163200 270370 164400
rect 271234 163200 271290 164400
rect 272062 163200 272118 164400
rect 272890 163200 272946 164400
rect 273718 163200 273774 164400
rect 274546 163200 274602 164400
rect 275374 163200 275430 164400
rect 276202 163200 276258 164400
rect 277122 163200 277178 164400
rect 277950 163200 278006 164400
rect 278778 163200 278834 164400
rect 279606 163200 279662 164400
rect 280434 163200 280490 164400
rect 281262 163200 281318 164400
rect 282090 163200 282146 164400
rect 283010 163200 283066 164400
rect 283838 163200 283894 164400
rect 284666 163200 284722 164400
rect 285494 163200 285550 164400
rect 286322 163200 286378 164400
rect 287150 163200 287206 164400
rect 287978 163200 288034 164400
rect 288898 163200 288954 164400
rect 289726 163200 289782 164400
rect 290554 163200 290610 164400
rect 291382 163200 291438 164400
rect 292210 163200 292266 164400
rect 293038 163200 293094 164400
rect 293866 163200 293922 164400
rect 294786 163200 294842 164400
rect 295614 163200 295670 164400
rect 296442 163200 296498 164400
rect 297270 163200 297326 164400
rect 298098 163200 298154 164400
rect 298926 163200 298982 164400
rect 299754 163200 299810 164400
rect 300674 163200 300730 164400
rect 301502 163200 301558 164400
rect 302330 163200 302386 164400
rect 303158 163200 303214 164400
rect 303986 163200 304042 164400
rect 304814 163200 304870 164400
rect 305642 163200 305698 164400
rect 306562 163200 306618 164400
rect 307390 163200 307446 164400
rect 308218 163200 308274 164400
rect 309046 163200 309102 164400
rect 309874 163200 309930 164400
rect 310702 163200 310758 164400
rect 311530 163200 311586 164400
rect 312450 163200 312506 164400
rect 313278 163200 313334 164400
rect 314106 163200 314162 164400
rect 314934 163200 314990 164400
rect 315762 163200 315818 164400
rect 316590 163200 316646 164400
rect 317418 163200 317474 164400
rect 318338 163200 318394 164400
rect 319166 163200 319222 164400
rect 319994 163200 320050 164400
rect 320822 163200 320878 164400
rect 321650 163200 321706 164400
rect 322478 163200 322534 164400
rect 323306 163200 323362 164400
rect 324226 163200 324282 164400
rect 325054 163200 325110 164400
rect 325882 163200 325938 164400
rect 326710 163200 326766 164400
rect 327538 163200 327594 164400
rect 328366 163200 328422 164400
rect 329194 163200 329250 164400
rect 330114 163200 330170 164400
rect 330942 163200 330998 164400
rect 331770 163200 331826 164400
rect 332598 163200 332654 164400
rect 333426 163200 333482 164400
rect 334254 163200 334310 164400
rect 335082 163200 335138 164400
rect 336002 163200 336058 164400
rect 336830 163200 336886 164400
rect 337658 163200 337714 164400
rect 338486 163200 338542 164400
rect 339314 163200 339370 164400
rect 340142 163200 340198 164400
rect 340970 163200 341026 164400
rect 341890 163200 341946 164400
rect 342718 163200 342774 164400
rect 343546 163200 343602 164400
rect 344374 163200 344430 164400
rect 345202 163200 345258 164400
rect 346030 163200 346086 164400
rect 346858 163200 346914 164400
rect 347778 163200 347834 164400
rect 348606 163200 348662 164400
rect 349434 163200 349490 164400
rect 350262 163200 350318 164400
rect 351090 163200 351146 164400
rect 351918 163200 351974 164400
rect 352746 163200 352802 164400
rect 353666 163200 353722 164400
rect 354494 163200 354550 164400
rect 355322 163200 355378 164400
rect 356150 163200 356206 164400
rect 356978 163200 357034 164400
rect 357806 163200 357862 164400
rect 358634 163200 358690 164400
rect 359554 163200 359610 164400
rect 360382 163200 360438 164400
rect 361210 163200 361266 164400
rect 362038 163200 362094 164400
rect 362866 163200 362922 164400
rect 363694 163200 363750 164400
rect 364522 163200 364578 164400
rect 365442 163200 365498 164400
rect 366270 163200 366326 164400
rect 367098 163200 367154 164400
rect 367926 163200 367982 164400
rect 368754 163200 368810 164400
rect 369582 163200 369638 164400
rect 370410 163200 370466 164400
rect 371330 163200 371386 164400
rect 372158 163200 372214 164400
rect 372986 163200 373042 164400
rect 373814 163200 373870 164400
rect 374642 163200 374698 164400
rect 375470 163200 375526 164400
rect 376298 163200 376354 164400
rect 377218 163200 377274 164400
rect 378046 163200 378102 164400
rect 378874 163200 378930 164400
rect 379702 163200 379758 164400
rect 380530 163200 380586 164400
rect 381358 163200 381414 164400
rect 382186 163200 382242 164400
rect 383106 163200 383162 164400
rect 383934 163200 383990 164400
rect 384762 163200 384818 164400
rect 385590 163200 385646 164400
rect 386418 163200 386474 164400
rect 387246 163200 387302 164400
rect 388074 163200 388130 164400
rect 388994 163200 389050 164400
rect 389822 163200 389878 164400
rect 390650 163200 390706 164400
rect 391478 163200 391534 164400
rect 392306 163200 392362 164400
rect 393134 163200 393190 164400
rect 393962 163200 394018 164400
rect 394882 163200 394938 164400
rect 395710 163200 395766 164400
rect 396538 163200 396594 164400
rect 397366 163200 397422 164400
rect 398194 163200 398250 164400
rect 399022 163200 399078 164400
rect 399850 163200 399906 164400
rect 400770 163200 400826 164400
rect 401598 163200 401654 164400
rect 402426 163200 402482 164400
rect 403254 163200 403310 164400
rect 404082 163200 404138 164400
rect 404910 163200 404966 164400
rect 405738 163200 405794 164400
rect 406658 163200 406714 164400
rect 407486 163200 407542 164400
rect 408314 163200 408370 164400
rect 409142 163200 409198 164400
rect 409970 163200 410026 164400
rect 410798 163200 410854 164400
rect 411626 163200 411682 164400
rect 412546 163200 412602 164400
rect 413374 163200 413430 164400
rect 414202 163200 414258 164400
rect 415030 163200 415086 164400
rect 415858 163200 415914 164400
rect 416686 163200 416742 164400
rect 417514 163200 417570 164400
rect 418434 163200 418490 164400
rect 419262 163200 419318 164400
rect 420090 163200 420146 164400
rect 420918 163200 420974 164400
rect 421746 163200 421802 164400
rect 422574 163200 422630 164400
rect 423402 163200 423458 164400
rect 424322 163200 424378 164400
rect 425150 163200 425206 164400
rect 425978 163200 426034 164400
rect 426806 163200 426862 164400
rect 427634 163200 427690 164400
rect 428462 163200 428518 164400
rect 429290 163200 429346 164400
rect 430210 163200 430266 164400
rect 431038 163200 431094 164400
rect 431866 163200 431922 164400
rect 432694 163200 432750 164400
rect 433522 163200 433578 164400
rect 434350 163200 434406 164400
rect 435178 163200 435234 164400
rect 436098 163200 436154 164400
rect 436926 163200 436982 164400
rect 437754 163200 437810 164400
rect 438582 163200 438638 164400
rect 439410 163200 439466 164400
rect 440238 163200 440294 164400
rect 441066 163200 441122 164400
rect 441986 163200 442042 164400
rect 442814 163200 442870 164400
rect 443642 163200 443698 164400
rect 444470 163200 444526 164400
rect 445298 163200 445354 164400
rect 446126 163200 446182 164400
rect 446954 163200 447010 164400
rect 447874 163200 447930 164400
rect 448702 163200 448758 164400
rect 449530 163200 449586 164400
rect 450358 163200 450414 164400
rect 451186 163200 451242 164400
rect 452014 163200 452070 164400
rect 452842 163200 452898 164400
rect 453762 163200 453818 164400
rect 454590 163200 454646 164400
rect 455418 163200 455474 164400
rect 456246 163200 456302 164400
rect 457074 163200 457130 164400
rect 457902 163200 457958 164400
rect 458730 163200 458786 164400
rect 459650 163200 459706 164400
rect 460478 163200 460534 164400
rect 461306 163200 461362 164400
rect 462134 163200 462190 164400
rect 462962 163200 463018 164400
rect 463790 163200 463846 164400
rect 464618 163200 464674 164400
rect 465538 163200 465594 164400
rect 466366 163200 466422 164400
rect 467194 163200 467250 164400
rect 468022 163200 468078 164400
rect 468850 163200 468906 164400
rect 469678 163200 469734 164400
rect 470506 163200 470562 164400
rect 471426 163200 471482 164400
rect 472254 163200 472310 164400
rect 473082 163200 473138 164400
rect 473910 163200 473966 164400
rect 474738 163200 474794 164400
rect 475566 163200 475622 164400
rect 476394 163200 476450 164400
rect 477314 163200 477370 164400
rect 478142 163200 478198 164400
rect 478970 163200 479026 164400
rect 479798 163200 479854 164400
rect 480626 163200 480682 164400
rect 481454 163200 481510 164400
rect 482282 163200 482338 164400
rect 483202 163200 483258 164400
rect 484030 163200 484086 164400
rect 484858 163200 484914 164400
rect 485686 163200 485742 164400
rect 486514 163200 486570 164400
rect 487342 163200 487398 164400
rect 488170 163200 488226 164400
rect 489090 163200 489146 164400
rect 489918 163200 489974 164400
rect 490746 163200 490802 164400
rect 491574 163200 491630 164400
rect 492402 163200 492458 164400
rect 493230 163200 493286 164400
rect 494058 163200 494114 164400
rect 494978 163200 495034 164400
rect 495806 163200 495862 164400
rect 496634 163200 496690 164400
rect 497462 163200 497518 164400
rect 498290 163200 498346 164400
rect 499118 163200 499174 164400
rect 499946 163200 500002 164400
rect 500866 163200 500922 164400
rect 501694 163200 501750 164400
rect 502522 163200 502578 164400
rect 503350 163200 503406 164400
rect 504178 163200 504234 164400
rect 505006 163200 505062 164400
rect 505834 163200 505890 164400
rect 506754 163200 506810 164400
rect 507582 163200 507638 164400
rect 508410 163200 508466 164400
rect 509238 163200 509294 164400
rect 510066 163200 510122 164400
rect 510894 163200 510950 164400
rect 511722 163200 511778 164400
rect 512642 163200 512698 164400
rect 513470 163200 513526 164400
rect 514298 163200 514354 164400
rect 515126 163200 515182 164400
rect 515954 163200 516010 164400
rect 516782 163200 516838 164400
rect 517610 163200 517666 164400
rect 518530 163200 518586 164400
rect 519358 163200 519414 164400
rect 520186 163200 520242 164400
rect 521014 163200 521070 164400
rect 521842 163200 521898 164400
rect 522670 163200 522726 164400
rect 523498 163200 523554 164400
rect 32770 -400 32826 800
rect 98274 -400 98330 800
rect 163778 -400 163834 800
rect 229282 -400 229338 800
rect 294786 -400 294842 800
rect 360290 -400 360346 800
rect 425794 -400 425850 800
rect 491298 -400 491354 800
<< obsm2 >>
rect 498 163144 1158 163282
rect 1326 163144 1986 163282
rect 2154 163144 2814 163282
rect 2982 163144 3642 163282
rect 3810 163144 4470 163282
rect 4638 163144 5298 163282
rect 5466 163144 6218 163282
rect 6386 163144 7046 163282
rect 7214 163144 7874 163282
rect 8042 163144 8702 163282
rect 8870 163144 9530 163282
rect 9698 163144 10358 163282
rect 10526 163144 11186 163282
rect 11354 163144 12106 163282
rect 12274 163144 12934 163282
rect 13102 163144 13762 163282
rect 13930 163144 14590 163282
rect 14758 163144 15418 163282
rect 15586 163144 16246 163282
rect 16414 163144 17074 163282
rect 17242 163144 17994 163282
rect 18162 163144 18822 163282
rect 18990 163144 19650 163282
rect 19818 163144 20478 163282
rect 20646 163144 21306 163282
rect 21474 163144 22134 163282
rect 22302 163144 22962 163282
rect 23130 163144 23882 163282
rect 24050 163144 24710 163282
rect 24878 163144 25538 163282
rect 25706 163144 26366 163282
rect 26534 163144 27194 163282
rect 27362 163144 28022 163282
rect 28190 163144 28850 163282
rect 29018 163144 29770 163282
rect 29938 163144 30598 163282
rect 30766 163144 31426 163282
rect 31594 163144 32254 163282
rect 32422 163144 33082 163282
rect 33250 163144 33910 163282
rect 34078 163144 34738 163282
rect 34906 163144 35658 163282
rect 35826 163144 36486 163282
rect 36654 163144 37314 163282
rect 37482 163144 38142 163282
rect 38310 163144 38970 163282
rect 39138 163144 39798 163282
rect 39966 163144 40626 163282
rect 40794 163144 41546 163282
rect 41714 163144 42374 163282
rect 42542 163144 43202 163282
rect 43370 163144 44030 163282
rect 44198 163144 44858 163282
rect 45026 163144 45686 163282
rect 45854 163144 46514 163282
rect 46682 163144 47434 163282
rect 47602 163144 48262 163282
rect 48430 163144 49090 163282
rect 49258 163144 49918 163282
rect 50086 163144 50746 163282
rect 50914 163144 51574 163282
rect 51742 163144 52402 163282
rect 52570 163144 53322 163282
rect 53490 163144 54150 163282
rect 54318 163144 54978 163282
rect 55146 163144 55806 163282
rect 55974 163144 56634 163282
rect 56802 163144 57462 163282
rect 57630 163144 58290 163282
rect 58458 163144 59210 163282
rect 59378 163144 60038 163282
rect 60206 163144 60866 163282
rect 61034 163144 61694 163282
rect 61862 163144 62522 163282
rect 62690 163144 63350 163282
rect 63518 163144 64178 163282
rect 64346 163144 65098 163282
rect 65266 163144 65926 163282
rect 66094 163144 66754 163282
rect 66922 163144 67582 163282
rect 67750 163144 68410 163282
rect 68578 163144 69238 163282
rect 69406 163144 70066 163282
rect 70234 163144 70986 163282
rect 71154 163144 71814 163282
rect 71982 163144 72642 163282
rect 72810 163144 73470 163282
rect 73638 163144 74298 163282
rect 74466 163144 75126 163282
rect 75294 163144 75954 163282
rect 76122 163144 76874 163282
rect 77042 163144 77702 163282
rect 77870 163144 78530 163282
rect 78698 163144 79358 163282
rect 79526 163144 80186 163282
rect 80354 163144 81014 163282
rect 81182 163144 81842 163282
rect 82010 163144 82762 163282
rect 82930 163144 83590 163282
rect 83758 163144 84418 163282
rect 84586 163144 85246 163282
rect 85414 163144 86074 163282
rect 86242 163144 86902 163282
rect 87070 163144 87730 163282
rect 87898 163144 88650 163282
rect 88818 163144 89478 163282
rect 89646 163144 90306 163282
rect 90474 163144 91134 163282
rect 91302 163144 91962 163282
rect 92130 163144 92790 163282
rect 92958 163144 93618 163282
rect 93786 163144 94538 163282
rect 94706 163144 95366 163282
rect 95534 163144 96194 163282
rect 96362 163144 97022 163282
rect 97190 163144 97850 163282
rect 98018 163144 98678 163282
rect 98846 163144 99506 163282
rect 99674 163144 100426 163282
rect 100594 163144 101254 163282
rect 101422 163144 102082 163282
rect 102250 163144 102910 163282
rect 103078 163144 103738 163282
rect 103906 163144 104566 163282
rect 104734 163144 105394 163282
rect 105562 163144 106314 163282
rect 106482 163144 107142 163282
rect 107310 163144 107970 163282
rect 108138 163144 108798 163282
rect 108966 163144 109626 163282
rect 109794 163144 110454 163282
rect 110622 163144 111282 163282
rect 111450 163144 112202 163282
rect 112370 163144 113030 163282
rect 113198 163144 113858 163282
rect 114026 163144 114686 163282
rect 114854 163144 115514 163282
rect 115682 163144 116342 163282
rect 116510 163144 117170 163282
rect 117338 163144 118090 163282
rect 118258 163144 118918 163282
rect 119086 163144 119746 163282
rect 119914 163144 120574 163282
rect 120742 163144 121402 163282
rect 121570 163144 122230 163282
rect 122398 163144 123058 163282
rect 123226 163144 123978 163282
rect 124146 163144 124806 163282
rect 124974 163144 125634 163282
rect 125802 163144 126462 163282
rect 126630 163144 127290 163282
rect 127458 163144 128118 163282
rect 128286 163144 128946 163282
rect 129114 163144 129866 163282
rect 130034 163144 130694 163282
rect 130862 163144 131522 163282
rect 131690 163144 132350 163282
rect 132518 163144 133178 163282
rect 133346 163144 134006 163282
rect 134174 163144 134834 163282
rect 135002 163144 135754 163282
rect 135922 163144 136582 163282
rect 136750 163144 137410 163282
rect 137578 163144 138238 163282
rect 138406 163144 139066 163282
rect 139234 163144 139894 163282
rect 140062 163144 140722 163282
rect 140890 163144 141642 163282
rect 141810 163144 142470 163282
rect 142638 163144 143298 163282
rect 143466 163144 144126 163282
rect 144294 163144 144954 163282
rect 145122 163144 145782 163282
rect 145950 163144 146610 163282
rect 146778 163144 147530 163282
rect 147698 163144 148358 163282
rect 148526 163144 149186 163282
rect 149354 163144 150014 163282
rect 150182 163144 150842 163282
rect 151010 163144 151670 163282
rect 151838 163144 152498 163282
rect 152666 163144 153418 163282
rect 153586 163144 154246 163282
rect 154414 163144 155074 163282
rect 155242 163144 155902 163282
rect 156070 163144 156730 163282
rect 156898 163144 157558 163282
rect 157726 163144 158386 163282
rect 158554 163144 159306 163282
rect 159474 163144 160134 163282
rect 160302 163144 160962 163282
rect 161130 163144 161790 163282
rect 161958 163144 162618 163282
rect 162786 163144 163446 163282
rect 163614 163144 164274 163282
rect 164442 163144 165194 163282
rect 165362 163144 166022 163282
rect 166190 163144 166850 163282
rect 167018 163144 167678 163282
rect 167846 163144 168506 163282
rect 168674 163144 169334 163282
rect 169502 163144 170162 163282
rect 170330 163144 171082 163282
rect 171250 163144 171910 163282
rect 172078 163144 172738 163282
rect 172906 163144 173566 163282
rect 173734 163144 174394 163282
rect 174562 163144 175222 163282
rect 175390 163144 176050 163282
rect 176218 163144 176970 163282
rect 177138 163144 177798 163282
rect 177966 163144 178626 163282
rect 178794 163144 179454 163282
rect 179622 163144 180282 163282
rect 180450 163144 181110 163282
rect 181278 163144 181938 163282
rect 182106 163144 182858 163282
rect 183026 163144 183686 163282
rect 183854 163144 184514 163282
rect 184682 163144 185342 163282
rect 185510 163144 186170 163282
rect 186338 163144 186998 163282
rect 187166 163144 187826 163282
rect 187994 163144 188746 163282
rect 188914 163144 189574 163282
rect 189742 163144 190402 163282
rect 190570 163144 191230 163282
rect 191398 163144 192058 163282
rect 192226 163144 192886 163282
rect 193054 163144 193714 163282
rect 193882 163144 194634 163282
rect 194802 163144 195462 163282
rect 195630 163144 196290 163282
rect 196458 163144 197118 163282
rect 197286 163144 197946 163282
rect 198114 163144 198774 163282
rect 198942 163144 199602 163282
rect 199770 163144 200522 163282
rect 200690 163144 201350 163282
rect 201518 163144 202178 163282
rect 202346 163144 203006 163282
rect 203174 163144 203834 163282
rect 204002 163144 204662 163282
rect 204830 163144 205490 163282
rect 205658 163144 206410 163282
rect 206578 163144 207238 163282
rect 207406 163144 208066 163282
rect 208234 163144 208894 163282
rect 209062 163144 209722 163282
rect 209890 163144 210550 163282
rect 210718 163144 211378 163282
rect 211546 163144 212298 163282
rect 212466 163144 213126 163282
rect 213294 163144 213954 163282
rect 214122 163144 214782 163282
rect 214950 163144 215610 163282
rect 215778 163144 216438 163282
rect 216606 163144 217266 163282
rect 217434 163144 218186 163282
rect 218354 163144 219014 163282
rect 219182 163144 219842 163282
rect 220010 163144 220670 163282
rect 220838 163144 221498 163282
rect 221666 163144 222326 163282
rect 222494 163144 223154 163282
rect 223322 163144 224074 163282
rect 224242 163144 224902 163282
rect 225070 163144 225730 163282
rect 225898 163144 226558 163282
rect 226726 163144 227386 163282
rect 227554 163144 228214 163282
rect 228382 163144 229042 163282
rect 229210 163144 229962 163282
rect 230130 163144 230790 163282
rect 230958 163144 231618 163282
rect 231786 163144 232446 163282
rect 232614 163144 233274 163282
rect 233442 163144 234102 163282
rect 234270 163144 234930 163282
rect 235098 163144 235850 163282
rect 236018 163144 236678 163282
rect 236846 163144 237506 163282
rect 237674 163144 238334 163282
rect 238502 163144 239162 163282
rect 239330 163144 239990 163282
rect 240158 163144 240818 163282
rect 240986 163144 241738 163282
rect 241906 163144 242566 163282
rect 242734 163144 243394 163282
rect 243562 163144 244222 163282
rect 244390 163144 245050 163282
rect 245218 163144 245878 163282
rect 246046 163144 246706 163282
rect 246874 163144 247626 163282
rect 247794 163144 248454 163282
rect 248622 163144 249282 163282
rect 249450 163144 250110 163282
rect 250278 163144 250938 163282
rect 251106 163144 251766 163282
rect 251934 163144 252594 163282
rect 252762 163144 253514 163282
rect 253682 163144 254342 163282
rect 254510 163144 255170 163282
rect 255338 163144 255998 163282
rect 256166 163144 256826 163282
rect 256994 163144 257654 163282
rect 257822 163144 258482 163282
rect 258650 163144 259402 163282
rect 259570 163144 260230 163282
rect 260398 163144 261058 163282
rect 261226 163144 261886 163282
rect 262054 163144 262714 163282
rect 262882 163144 263542 163282
rect 263710 163144 264370 163282
rect 264538 163144 265290 163282
rect 265458 163144 266118 163282
rect 266286 163144 266946 163282
rect 267114 163144 267774 163282
rect 267942 163144 268602 163282
rect 268770 163144 269430 163282
rect 269598 163144 270258 163282
rect 270426 163144 271178 163282
rect 271346 163144 272006 163282
rect 272174 163144 272834 163282
rect 273002 163144 273662 163282
rect 273830 163144 274490 163282
rect 274658 163144 275318 163282
rect 275486 163144 276146 163282
rect 276314 163144 277066 163282
rect 277234 163144 277894 163282
rect 278062 163144 278722 163282
rect 278890 163144 279550 163282
rect 279718 163144 280378 163282
rect 280546 163144 281206 163282
rect 281374 163144 282034 163282
rect 282202 163144 282954 163282
rect 283122 163144 283782 163282
rect 283950 163144 284610 163282
rect 284778 163144 285438 163282
rect 285606 163144 286266 163282
rect 286434 163144 287094 163282
rect 287262 163144 287922 163282
rect 288090 163144 288842 163282
rect 289010 163144 289670 163282
rect 289838 163144 290498 163282
rect 290666 163144 291326 163282
rect 291494 163144 292154 163282
rect 292322 163144 292982 163282
rect 293150 163144 293810 163282
rect 293978 163144 294730 163282
rect 294898 163144 295558 163282
rect 295726 163144 296386 163282
rect 296554 163144 297214 163282
rect 297382 163144 298042 163282
rect 298210 163144 298870 163282
rect 299038 163144 299698 163282
rect 299866 163144 300618 163282
rect 300786 163144 301446 163282
rect 301614 163144 302274 163282
rect 302442 163144 303102 163282
rect 303270 163144 303930 163282
rect 304098 163144 304758 163282
rect 304926 163144 305586 163282
rect 305754 163144 306506 163282
rect 306674 163144 307334 163282
rect 307502 163144 308162 163282
rect 308330 163144 308990 163282
rect 309158 163144 309818 163282
rect 309986 163144 310646 163282
rect 310814 163144 311474 163282
rect 311642 163144 312394 163282
rect 312562 163144 313222 163282
rect 313390 163144 314050 163282
rect 314218 163144 314878 163282
rect 315046 163144 315706 163282
rect 315874 163144 316534 163282
rect 316702 163144 317362 163282
rect 317530 163144 318282 163282
rect 318450 163144 319110 163282
rect 319278 163144 319938 163282
rect 320106 163144 320766 163282
rect 320934 163144 321594 163282
rect 321762 163144 322422 163282
rect 322590 163144 323250 163282
rect 323418 163144 324170 163282
rect 324338 163144 324998 163282
rect 325166 163144 325826 163282
rect 325994 163144 326654 163282
rect 326822 163144 327482 163282
rect 327650 163144 328310 163282
rect 328478 163144 329138 163282
rect 329306 163144 330058 163282
rect 330226 163144 330886 163282
rect 331054 163144 331714 163282
rect 331882 163144 332542 163282
rect 332710 163144 333370 163282
rect 333538 163144 334198 163282
rect 334366 163144 335026 163282
rect 335194 163144 335946 163282
rect 336114 163144 336774 163282
rect 336942 163144 337602 163282
rect 337770 163144 338430 163282
rect 338598 163144 339258 163282
rect 339426 163144 340086 163282
rect 340254 163144 340914 163282
rect 341082 163144 341834 163282
rect 342002 163144 342662 163282
rect 342830 163144 343490 163282
rect 343658 163144 344318 163282
rect 344486 163144 345146 163282
rect 345314 163144 345974 163282
rect 346142 163144 346802 163282
rect 346970 163144 347722 163282
rect 347890 163144 348550 163282
rect 348718 163144 349378 163282
rect 349546 163144 350206 163282
rect 350374 163144 351034 163282
rect 351202 163144 351862 163282
rect 352030 163144 352690 163282
rect 352858 163144 353610 163282
rect 353778 163144 354438 163282
rect 354606 163144 355266 163282
rect 355434 163144 356094 163282
rect 356262 163144 356922 163282
rect 357090 163144 357750 163282
rect 357918 163144 358578 163282
rect 358746 163144 359498 163282
rect 359666 163144 360326 163282
rect 360494 163144 361154 163282
rect 361322 163144 361982 163282
rect 362150 163144 362810 163282
rect 362978 163144 363638 163282
rect 363806 163144 364466 163282
rect 364634 163144 365386 163282
rect 365554 163144 366214 163282
rect 366382 163144 367042 163282
rect 367210 163144 367870 163282
rect 368038 163144 368698 163282
rect 368866 163144 369526 163282
rect 369694 163144 370354 163282
rect 370522 163144 371274 163282
rect 371442 163144 372102 163282
rect 372270 163144 372930 163282
rect 373098 163144 373758 163282
rect 373926 163144 374586 163282
rect 374754 163144 375414 163282
rect 375582 163144 376242 163282
rect 376410 163144 377162 163282
rect 377330 163144 377990 163282
rect 378158 163144 378818 163282
rect 378986 163144 379646 163282
rect 379814 163144 380474 163282
rect 380642 163144 381302 163282
rect 381470 163144 382130 163282
rect 382298 163144 383050 163282
rect 383218 163144 383878 163282
rect 384046 163144 384706 163282
rect 384874 163144 385534 163282
rect 385702 163144 386362 163282
rect 386530 163144 387190 163282
rect 387358 163144 388018 163282
rect 388186 163144 388938 163282
rect 389106 163144 389766 163282
rect 389934 163144 390594 163282
rect 390762 163144 391422 163282
rect 391590 163144 392250 163282
rect 392418 163144 393078 163282
rect 393246 163144 393906 163282
rect 394074 163144 394826 163282
rect 394994 163144 395654 163282
rect 395822 163144 396482 163282
rect 396650 163144 397310 163282
rect 397478 163144 398138 163282
rect 398306 163144 398966 163282
rect 399134 163144 399794 163282
rect 399962 163144 400714 163282
rect 400882 163144 401542 163282
rect 401710 163144 402370 163282
rect 402538 163144 403198 163282
rect 403366 163144 404026 163282
rect 404194 163144 404854 163282
rect 405022 163144 405682 163282
rect 405850 163144 406602 163282
rect 406770 163144 407430 163282
rect 407598 163144 408258 163282
rect 408426 163144 409086 163282
rect 409254 163144 409914 163282
rect 410082 163144 410742 163282
rect 410910 163144 411570 163282
rect 411738 163144 412490 163282
rect 412658 163144 413318 163282
rect 413486 163144 414146 163282
rect 414314 163144 414974 163282
rect 415142 163144 415802 163282
rect 415970 163144 416630 163282
rect 416798 163144 417458 163282
rect 417626 163144 418378 163282
rect 418546 163144 419206 163282
rect 419374 163144 420034 163282
rect 420202 163144 420862 163282
rect 421030 163144 421690 163282
rect 421858 163144 422518 163282
rect 422686 163144 423346 163282
rect 423514 163144 424266 163282
rect 424434 163144 425094 163282
rect 425262 163144 425922 163282
rect 426090 163144 426750 163282
rect 426918 163144 427578 163282
rect 427746 163144 428406 163282
rect 428574 163144 429234 163282
rect 429402 163144 430154 163282
rect 430322 163144 430982 163282
rect 431150 163144 431810 163282
rect 431978 163144 432638 163282
rect 432806 163144 433466 163282
rect 433634 163144 434294 163282
rect 434462 163144 435122 163282
rect 435290 163144 436042 163282
rect 436210 163144 436870 163282
rect 437038 163144 437698 163282
rect 437866 163144 438526 163282
rect 438694 163144 439354 163282
rect 439522 163144 440182 163282
rect 440350 163144 441010 163282
rect 441178 163144 441930 163282
rect 442098 163144 442758 163282
rect 442926 163144 443586 163282
rect 443754 163144 444414 163282
rect 444582 163144 445242 163282
rect 445410 163144 446070 163282
rect 446238 163144 446898 163282
rect 447066 163144 447818 163282
rect 447986 163144 448646 163282
rect 448814 163144 449474 163282
rect 449642 163144 450302 163282
rect 450470 163144 451130 163282
rect 451298 163144 451958 163282
rect 452126 163144 452786 163282
rect 452954 163144 453706 163282
rect 453874 163144 454534 163282
rect 454702 163144 455362 163282
rect 455530 163144 456190 163282
rect 456358 163144 457018 163282
rect 457186 163144 457846 163282
rect 458014 163144 458674 163282
rect 458842 163144 459594 163282
rect 459762 163144 460422 163282
rect 460590 163144 461250 163282
rect 461418 163144 462078 163282
rect 462246 163144 462906 163282
rect 463074 163144 463734 163282
rect 463902 163144 464562 163282
rect 464730 163144 465482 163282
rect 465650 163144 466310 163282
rect 466478 163144 467138 163282
rect 467306 163144 467966 163282
rect 468134 163144 468794 163282
rect 468962 163144 469622 163282
rect 469790 163144 470450 163282
rect 470618 163144 471370 163282
rect 471538 163144 472198 163282
rect 472366 163144 473026 163282
rect 473194 163144 473854 163282
rect 474022 163144 474682 163282
rect 474850 163144 475510 163282
rect 475678 163144 476338 163282
rect 476506 163144 477258 163282
rect 477426 163144 478086 163282
rect 478254 163144 478914 163282
rect 479082 163144 479742 163282
rect 479910 163144 480570 163282
rect 480738 163144 481398 163282
rect 481566 163144 482226 163282
rect 482394 163144 483146 163282
rect 483314 163144 483974 163282
rect 484142 163144 484802 163282
rect 484970 163144 485630 163282
rect 485798 163144 486458 163282
rect 486626 163144 487286 163282
rect 487454 163144 488114 163282
rect 488282 163144 489034 163282
rect 489202 163144 489862 163282
rect 490030 163144 490690 163282
rect 490858 163144 491518 163282
rect 491686 163144 492346 163282
rect 492514 163144 493174 163282
rect 493342 163144 494002 163282
rect 494170 163144 494922 163282
rect 495090 163144 495750 163282
rect 495918 163144 496578 163282
rect 496746 163144 497406 163282
rect 497574 163144 498234 163282
rect 498402 163144 499062 163282
rect 499230 163144 499890 163282
rect 500058 163144 500810 163282
rect 500978 163144 501638 163282
rect 501806 163144 502466 163282
rect 502634 163144 503294 163282
rect 503462 163144 504122 163282
rect 504290 163144 504950 163282
rect 505118 163144 505778 163282
rect 505946 163144 506698 163282
rect 506866 163144 507526 163282
rect 507694 163144 508354 163282
rect 508522 163144 509182 163282
rect 509350 163144 510010 163282
rect 510178 163144 510838 163282
rect 511006 163144 511666 163282
rect 511834 163144 512586 163282
rect 512754 163144 513414 163282
rect 513582 163144 514242 163282
rect 514410 163144 515070 163282
rect 515238 163144 515898 163282
rect 516066 163144 516726 163282
rect 516894 163144 517554 163282
rect 517722 163144 518474 163282
rect 518642 163144 519302 163282
rect 519470 163144 520130 163282
rect 520298 163144 520958 163282
rect 521126 163144 521786 163282
rect 521954 163144 522614 163282
rect 522782 163144 523442 163282
rect 388 856 523552 163144
rect 388 711 32714 856
rect 32882 711 98218 856
rect 98386 711 163722 856
rect 163890 711 229226 856
rect 229394 711 294730 856
rect 294898 711 360234 856
rect 360402 711 425738 856
rect 425906 711 491242 856
rect 491410 711 523552 856
<< metal3 >>
rect 523200 163072 524400 163192
rect 523200 161576 524400 161696
rect 523200 160080 524400 160200
rect 523200 158584 524400 158704
rect 523200 157088 524400 157208
rect 523200 155592 524400 155712
rect 523200 154096 524400 154216
rect 523200 152600 524400 152720
rect 523200 151104 524400 151224
rect 523200 149608 524400 149728
rect 523200 148112 524400 148232
rect 523200 146616 524400 146736
rect 523200 145120 524400 145240
rect 523200 143624 524400 143744
rect 523200 142128 524400 142248
rect 523200 140496 524400 140616
rect 523200 139000 524400 139120
rect 523200 137504 524400 137624
rect 523200 136008 524400 136128
rect 523200 134512 524400 134632
rect 523200 133016 524400 133136
rect 523200 131520 524400 131640
rect 523200 130024 524400 130144
rect 523200 128528 524400 128648
rect 523200 127032 524400 127152
rect 523200 125536 524400 125656
rect 523200 124040 524400 124160
rect 523200 122544 524400 122664
rect 523200 121048 524400 121168
rect 523200 119552 524400 119672
rect 523200 118056 524400 118176
rect 523200 116424 524400 116544
rect 523200 114928 524400 115048
rect 523200 113432 524400 113552
rect 523200 111936 524400 112056
rect 523200 110440 524400 110560
rect 523200 108944 524400 109064
rect 523200 107448 524400 107568
rect 523200 105952 524400 106072
rect 523200 104456 524400 104576
rect 523200 102960 524400 103080
rect 523200 101464 524400 101584
rect 523200 99968 524400 100088
rect 523200 98472 524400 98592
rect 523200 96976 524400 97096
rect 523200 95480 524400 95600
rect 523200 93848 524400 93968
rect 523200 92352 524400 92472
rect 523200 90856 524400 90976
rect 523200 89360 524400 89480
rect 523200 87864 524400 87984
rect 523200 86368 524400 86488
rect 523200 84872 524400 84992
rect 523200 83376 524400 83496
rect 523200 81880 524400 82000
rect 523200 80384 524400 80504
rect 523200 78888 524400 79008
rect 523200 77392 524400 77512
rect 523200 75896 524400 76016
rect 523200 74400 524400 74520
rect 523200 72904 524400 73024
rect 523200 71408 524400 71528
rect 523200 69776 524400 69896
rect 523200 68280 524400 68400
rect 523200 66784 524400 66904
rect 523200 65288 524400 65408
rect 523200 63792 524400 63912
rect 523200 62296 524400 62416
rect 523200 60800 524400 60920
rect 523200 59304 524400 59424
rect 523200 57808 524400 57928
rect 523200 56312 524400 56432
rect 523200 54816 524400 54936
rect 523200 53320 524400 53440
rect 523200 51824 524400 51944
rect 523200 50328 524400 50448
rect 523200 48832 524400 48952
rect 523200 47200 524400 47320
rect 523200 45704 524400 45824
rect 523200 44208 524400 44328
rect 523200 42712 524400 42832
rect 523200 41216 524400 41336
rect 523200 39720 524400 39840
rect 523200 38224 524400 38344
rect 523200 36728 524400 36848
rect 523200 35232 524400 35352
rect 523200 33736 524400 33856
rect 523200 32240 524400 32360
rect 523200 30744 524400 30864
rect 523200 29248 524400 29368
rect 523200 27752 524400 27872
rect 523200 26256 524400 26376
rect 523200 24760 524400 24880
rect 523200 23128 524400 23248
rect 523200 21632 524400 21752
rect 523200 20136 524400 20256
rect 523200 18640 524400 18760
rect 523200 17144 524400 17264
rect 523200 15648 524400 15768
rect 523200 14152 524400 14272
rect 523200 12656 524400 12776
rect 523200 11160 524400 11280
rect 523200 9664 524400 9784
rect 523200 8168 524400 8288
rect 523200 6672 524400 6792
rect 523200 5176 524400 5296
rect 523200 3680 524400 3800
rect 523200 2184 524400 2304
rect 523200 688 524400 808
<< obsm3 >>
rect 2669 162992 523120 163165
rect 2669 161776 523200 162992
rect 2669 161496 523120 161776
rect 2669 160280 523200 161496
rect 2669 160000 523120 160280
rect 2669 158784 523200 160000
rect 2669 158504 523120 158784
rect 2669 157288 523200 158504
rect 2669 157008 523120 157288
rect 2669 155792 523200 157008
rect 2669 155512 523120 155792
rect 2669 154296 523200 155512
rect 2669 154016 523120 154296
rect 2669 152800 523200 154016
rect 2669 152520 523120 152800
rect 2669 151304 523200 152520
rect 2669 151024 523120 151304
rect 2669 149808 523200 151024
rect 2669 149528 523120 149808
rect 2669 148312 523200 149528
rect 2669 148032 523120 148312
rect 2669 146816 523200 148032
rect 2669 146536 523120 146816
rect 2669 145320 523200 146536
rect 2669 145040 523120 145320
rect 2669 143824 523200 145040
rect 2669 143544 523120 143824
rect 2669 142328 523200 143544
rect 2669 142048 523120 142328
rect 2669 140696 523200 142048
rect 2669 140416 523120 140696
rect 2669 139200 523200 140416
rect 2669 138920 523120 139200
rect 2669 137704 523200 138920
rect 2669 137424 523120 137704
rect 2669 136208 523200 137424
rect 2669 135928 523120 136208
rect 2669 134712 523200 135928
rect 2669 134432 523120 134712
rect 2669 133216 523200 134432
rect 2669 132936 523120 133216
rect 2669 131720 523200 132936
rect 2669 131440 523120 131720
rect 2669 130224 523200 131440
rect 2669 129944 523120 130224
rect 2669 128728 523200 129944
rect 2669 128448 523120 128728
rect 2669 127232 523200 128448
rect 2669 126952 523120 127232
rect 2669 125736 523200 126952
rect 2669 125456 523120 125736
rect 2669 124240 523200 125456
rect 2669 123960 523120 124240
rect 2669 122744 523200 123960
rect 2669 122464 523120 122744
rect 2669 121248 523200 122464
rect 2669 120968 523120 121248
rect 2669 119752 523200 120968
rect 2669 119472 523120 119752
rect 2669 118256 523200 119472
rect 2669 117976 523120 118256
rect 2669 116624 523200 117976
rect 2669 116344 523120 116624
rect 2669 115128 523200 116344
rect 2669 114848 523120 115128
rect 2669 113632 523200 114848
rect 2669 113352 523120 113632
rect 2669 112136 523200 113352
rect 2669 111856 523120 112136
rect 2669 110640 523200 111856
rect 2669 110360 523120 110640
rect 2669 109144 523200 110360
rect 2669 108864 523120 109144
rect 2669 107648 523200 108864
rect 2669 107368 523120 107648
rect 2669 106152 523200 107368
rect 2669 105872 523120 106152
rect 2669 104656 523200 105872
rect 2669 104376 523120 104656
rect 2669 103160 523200 104376
rect 2669 102880 523120 103160
rect 2669 101664 523200 102880
rect 2669 101384 523120 101664
rect 2669 100168 523200 101384
rect 2669 99888 523120 100168
rect 2669 98672 523200 99888
rect 2669 98392 523120 98672
rect 2669 97176 523200 98392
rect 2669 96896 523120 97176
rect 2669 95680 523200 96896
rect 2669 95400 523120 95680
rect 2669 94048 523200 95400
rect 2669 93768 523120 94048
rect 2669 92552 523200 93768
rect 2669 92272 523120 92552
rect 2669 91056 523200 92272
rect 2669 90776 523120 91056
rect 2669 89560 523200 90776
rect 2669 89280 523120 89560
rect 2669 88064 523200 89280
rect 2669 87784 523120 88064
rect 2669 86568 523200 87784
rect 2669 86288 523120 86568
rect 2669 85072 523200 86288
rect 2669 84792 523120 85072
rect 2669 83576 523200 84792
rect 2669 83296 523120 83576
rect 2669 82080 523200 83296
rect 2669 81800 523120 82080
rect 2669 80584 523200 81800
rect 2669 80304 523120 80584
rect 2669 79088 523200 80304
rect 2669 78808 523120 79088
rect 2669 77592 523200 78808
rect 2669 77312 523120 77592
rect 2669 76096 523200 77312
rect 2669 75816 523120 76096
rect 2669 74600 523200 75816
rect 2669 74320 523120 74600
rect 2669 73104 523200 74320
rect 2669 72824 523120 73104
rect 2669 71608 523200 72824
rect 2669 71328 523120 71608
rect 2669 69976 523200 71328
rect 2669 69696 523120 69976
rect 2669 68480 523200 69696
rect 2669 68200 523120 68480
rect 2669 66984 523200 68200
rect 2669 66704 523120 66984
rect 2669 65488 523200 66704
rect 2669 65208 523120 65488
rect 2669 63992 523200 65208
rect 2669 63712 523120 63992
rect 2669 62496 523200 63712
rect 2669 62216 523120 62496
rect 2669 61000 523200 62216
rect 2669 60720 523120 61000
rect 2669 59504 523200 60720
rect 2669 59224 523120 59504
rect 2669 58008 523200 59224
rect 2669 57728 523120 58008
rect 2669 56512 523200 57728
rect 2669 56232 523120 56512
rect 2669 55016 523200 56232
rect 2669 54736 523120 55016
rect 2669 53520 523200 54736
rect 2669 53240 523120 53520
rect 2669 52024 523200 53240
rect 2669 51744 523120 52024
rect 2669 50528 523200 51744
rect 2669 50248 523120 50528
rect 2669 49032 523200 50248
rect 2669 48752 523120 49032
rect 2669 47400 523200 48752
rect 2669 47120 523120 47400
rect 2669 45904 523200 47120
rect 2669 45624 523120 45904
rect 2669 44408 523200 45624
rect 2669 44128 523120 44408
rect 2669 42912 523200 44128
rect 2669 42632 523120 42912
rect 2669 41416 523200 42632
rect 2669 41136 523120 41416
rect 2669 39920 523200 41136
rect 2669 39640 523120 39920
rect 2669 38424 523200 39640
rect 2669 38144 523120 38424
rect 2669 36928 523200 38144
rect 2669 36648 523120 36928
rect 2669 35432 523200 36648
rect 2669 35152 523120 35432
rect 2669 33936 523200 35152
rect 2669 33656 523120 33936
rect 2669 32440 523200 33656
rect 2669 32160 523120 32440
rect 2669 30944 523200 32160
rect 2669 30664 523120 30944
rect 2669 29448 523200 30664
rect 2669 29168 523120 29448
rect 2669 27952 523200 29168
rect 2669 27672 523120 27952
rect 2669 26456 523200 27672
rect 2669 26176 523120 26456
rect 2669 24960 523200 26176
rect 2669 24680 523120 24960
rect 2669 23328 523200 24680
rect 2669 23048 523120 23328
rect 2669 21832 523200 23048
rect 2669 21552 523120 21832
rect 2669 20336 523200 21552
rect 2669 20056 523120 20336
rect 2669 18840 523200 20056
rect 2669 18560 523120 18840
rect 2669 17344 523200 18560
rect 2669 17064 523120 17344
rect 2669 15848 523200 17064
rect 2669 15568 523120 15848
rect 2669 14352 523200 15568
rect 2669 14072 523120 14352
rect 2669 12856 523200 14072
rect 2669 12576 523120 12856
rect 2669 11360 523200 12576
rect 2669 11080 523120 11360
rect 2669 9864 523200 11080
rect 2669 9584 523120 9864
rect 2669 8368 523200 9584
rect 2669 8088 523120 8368
rect 2669 6872 523200 8088
rect 2669 6592 523120 6872
rect 2669 5376 523200 6592
rect 2669 5096 523120 5376
rect 2669 3880 523200 5096
rect 2669 3600 523120 3880
rect 2669 2384 523200 3600
rect 2669 2104 523120 2384
rect 2669 888 523200 2104
rect 2669 715 523120 888
<< obsm4 >>
rect 1004 1531 518920 149812
<< metal5 >>
rect 1104 156856 522836 157496
rect 1104 143856 2200 144496
rect 109800 143856 120200 144496
rect 517800 143856 522836 144496
rect 1104 130856 2200 131496
rect 109800 130856 120200 131496
rect 517800 130856 522836 131496
rect 1104 117856 2200 118496
rect 109800 117856 120200 118496
rect 517800 117856 522836 118496
rect 1104 104856 2200 105496
rect 109800 104856 120200 105496
rect 517800 104856 522836 105496
rect 1104 91856 2200 92496
rect 109800 91856 120200 92496
rect 517800 91856 522836 92496
rect 1104 78856 2200 79496
rect 109800 78856 120200 79496
rect 517800 78856 522836 79496
rect 1104 65856 2200 66496
rect 109800 65856 120200 66496
rect 517800 65856 522836 66496
rect 1104 52856 2200 53496
rect 109800 52856 120200 53496
rect 517800 52856 522836 53496
rect 1104 39856 2200 40496
rect 109800 39856 120200 40496
rect 517800 39856 522836 40496
rect 1104 26856 2200 27496
rect 109800 26856 120200 27496
rect 517800 26856 522836 27496
rect 1104 13856 2200 14496
rect 109800 13856 120200 14496
rect 517800 13856 522836 14496
<< obsm5 >>
rect 1004 144816 518920 149812
rect 2520 143536 109480 144816
rect 120520 143536 517480 144816
rect 1004 131816 518920 143536
rect 2520 130536 109480 131816
rect 120520 130536 517480 131816
rect 1004 118816 518920 130536
rect 2520 117536 109480 118816
rect 120520 117536 517480 118816
rect 1004 105816 518920 117536
rect 2520 104536 109480 105816
rect 120520 104536 517480 105816
rect 1004 92816 518920 104536
rect 2520 91536 109480 92816
rect 120520 91536 517480 92816
rect 1004 79816 518920 91536
rect 2520 78536 109480 79816
rect 120520 78536 517480 79816
rect 1004 66816 518920 78536
rect 2520 65536 109480 66816
rect 120520 65536 517480 66816
rect 1004 53816 518920 65536
rect 2520 52536 109480 53816
rect 120520 52536 517480 53816
rect 1004 40816 518920 52536
rect 2520 39536 109480 40816
rect 120520 39536 517480 40816
rect 1004 27816 518920 39536
rect 2520 26536 109480 27816
rect 120520 26536 517480 27816
rect 1004 14816 518920 26536
rect 2520 13536 109480 14816
rect 120520 13536 517480 14816
rect 1004 2156 518920 13536
<< labels >>
rlabel metal5 s 1104 26856 2200 27496 6 VGND
port 1 nsew ground input
rlabel metal5 s 109800 26856 120200 27496 6 VGND
port 1 nsew ground input
rlabel metal5 s 517800 26856 522836 27496 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 52856 2200 53496 6 VGND
port 1 nsew ground input
rlabel metal5 s 109800 52856 120200 53496 6 VGND
port 1 nsew ground input
rlabel metal5 s 517800 52856 522836 53496 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 78856 2200 79496 6 VGND
port 1 nsew ground input
rlabel metal5 s 109800 78856 120200 79496 6 VGND
port 1 nsew ground input
rlabel metal5 s 517800 78856 522836 79496 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 104856 2200 105496 6 VGND
port 1 nsew ground input
rlabel metal5 s 109800 104856 120200 105496 6 VGND
port 1 nsew ground input
rlabel metal5 s 517800 104856 522836 105496 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 130856 2200 131496 6 VGND
port 1 nsew ground input
rlabel metal5 s 109800 130856 120200 131496 6 VGND
port 1 nsew ground input
rlabel metal5 s 517800 130856 522836 131496 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 156856 522836 157496 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 13856 2200 14496 6 VPWR
port 2 nsew power input
rlabel metal5 s 109800 13856 120200 14496 6 VPWR
port 2 nsew power input
rlabel metal5 s 517800 13856 522836 14496 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 39856 2200 40496 6 VPWR
port 2 nsew power input
rlabel metal5 s 109800 39856 120200 40496 6 VPWR
port 2 nsew power input
rlabel metal5 s 517800 39856 522836 40496 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 65856 2200 66496 6 VPWR
port 2 nsew power input
rlabel metal5 s 109800 65856 120200 66496 6 VPWR
port 2 nsew power input
rlabel metal5 s 517800 65856 522836 66496 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 91856 2200 92496 6 VPWR
port 2 nsew power input
rlabel metal5 s 109800 91856 120200 92496 6 VPWR
port 2 nsew power input
rlabel metal5 s 517800 91856 522836 92496 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 117856 2200 118496 6 VPWR
port 2 nsew power input
rlabel metal5 s 109800 117856 120200 118496 6 VPWR
port 2 nsew power input
rlabel metal5 s 517800 117856 522836 118496 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 143856 2200 144496 6 VPWR
port 2 nsew power input
rlabel metal5 s 109800 143856 120200 144496 6 VPWR
port 2 nsew power input
rlabel metal5 s 517800 143856 522836 144496 6 VPWR
port 2 nsew power input
rlabel metal2 s 294786 -400 294842 800 6 core_clk
port 3 nsew signal input
rlabel metal2 s 98274 -400 98330 800 6 core_rstn
port 4 nsew signal input
rlabel metal3 s 523200 63792 524400 63912 6 debug_in
port 5 nsew signal input
rlabel metal3 s 523200 65288 524400 65408 6 debug_mode
port 6 nsew signal output
rlabel metal3 s 523200 66784 524400 66904 6 debug_oeb
port 7 nsew signal output
rlabel metal3 s 523200 68280 524400 68400 6 debug_out
port 8 nsew signal output
rlabel metal3 s 523200 145120 524400 145240 6 flash_clk
port 9 nsew signal output
rlabel metal3 s 523200 143624 524400 143744 6 flash_csb
port 10 nsew signal output
rlabel metal3 s 523200 146616 524400 146736 6 flash_io0_di
port 11 nsew signal input
rlabel metal3 s 523200 148112 524400 148232 6 flash_io0_do
port 12 nsew signal output
rlabel metal3 s 523200 149608 524400 149728 6 flash_io0_oeb
port 13 nsew signal output
rlabel metal3 s 523200 151104 524400 151224 6 flash_io1_di
port 14 nsew signal input
rlabel metal3 s 523200 152600 524400 152720 6 flash_io1_do
port 15 nsew signal output
rlabel metal3 s 523200 154096 524400 154216 6 flash_io1_oeb
port 16 nsew signal output
rlabel metal3 s 523200 155592 524400 155712 6 flash_io2_di
port 17 nsew signal input
rlabel metal3 s 523200 157088 524400 157208 6 flash_io2_do
port 18 nsew signal output
rlabel metal3 s 523200 158584 524400 158704 6 flash_io2_oeb
port 19 nsew signal output
rlabel metal3 s 523200 160080 524400 160200 6 flash_io3_di
port 20 nsew signal input
rlabel metal3 s 523200 161576 524400 161696 6 flash_io3_do
port 21 nsew signal output
rlabel metal3 s 523200 163072 524400 163192 6 flash_io3_oeb
port 22 nsew signal output
rlabel metal2 s 32770 -400 32826 800 6 gpio_in_pad
port 23 nsew signal input
rlabel metal2 s 163778 -400 163834 800 6 gpio_inenb_pad
port 24 nsew signal output
rlabel metal2 s 229282 -400 229338 800 6 gpio_mode0_pad
port 25 nsew signal output
rlabel metal2 s 360290 -400 360346 800 6 gpio_mode1_pad
port 26 nsew signal output
rlabel metal2 s 425794 -400 425850 800 6 gpio_out_pad
port 27 nsew signal output
rlabel metal2 s 491298 -400 491354 800 6 gpio_outenb_pad
port 28 nsew signal output
rlabel metal3 s 523200 90856 524400 90976 6 hk_ack_i
port 29 nsew signal input
rlabel metal3 s 523200 93848 524400 93968 6 hk_cyc_o
port 30 nsew signal output
rlabel metal3 s 523200 95480 524400 95600 6 hk_dat_i[0]
port 31 nsew signal input
rlabel metal3 s 523200 110440 524400 110560 6 hk_dat_i[10]
port 32 nsew signal input
rlabel metal3 s 523200 111936 524400 112056 6 hk_dat_i[11]
port 33 nsew signal input
rlabel metal3 s 523200 113432 524400 113552 6 hk_dat_i[12]
port 34 nsew signal input
rlabel metal3 s 523200 114928 524400 115048 6 hk_dat_i[13]
port 35 nsew signal input
rlabel metal3 s 523200 116424 524400 116544 6 hk_dat_i[14]
port 36 nsew signal input
rlabel metal3 s 523200 118056 524400 118176 6 hk_dat_i[15]
port 37 nsew signal input
rlabel metal3 s 523200 119552 524400 119672 6 hk_dat_i[16]
port 38 nsew signal input
rlabel metal3 s 523200 121048 524400 121168 6 hk_dat_i[17]
port 39 nsew signal input
rlabel metal3 s 523200 122544 524400 122664 6 hk_dat_i[18]
port 40 nsew signal input
rlabel metal3 s 523200 124040 524400 124160 6 hk_dat_i[19]
port 41 nsew signal input
rlabel metal3 s 523200 96976 524400 97096 6 hk_dat_i[1]
port 42 nsew signal input
rlabel metal3 s 523200 125536 524400 125656 6 hk_dat_i[20]
port 43 nsew signal input
rlabel metal3 s 523200 127032 524400 127152 6 hk_dat_i[21]
port 44 nsew signal input
rlabel metal3 s 523200 128528 524400 128648 6 hk_dat_i[22]
port 45 nsew signal input
rlabel metal3 s 523200 130024 524400 130144 6 hk_dat_i[23]
port 46 nsew signal input
rlabel metal3 s 523200 131520 524400 131640 6 hk_dat_i[24]
port 47 nsew signal input
rlabel metal3 s 523200 133016 524400 133136 6 hk_dat_i[25]
port 48 nsew signal input
rlabel metal3 s 523200 134512 524400 134632 6 hk_dat_i[26]
port 49 nsew signal input
rlabel metal3 s 523200 136008 524400 136128 6 hk_dat_i[27]
port 50 nsew signal input
rlabel metal3 s 523200 137504 524400 137624 6 hk_dat_i[28]
port 51 nsew signal input
rlabel metal3 s 523200 139000 524400 139120 6 hk_dat_i[29]
port 52 nsew signal input
rlabel metal3 s 523200 98472 524400 98592 6 hk_dat_i[2]
port 53 nsew signal input
rlabel metal3 s 523200 140496 524400 140616 6 hk_dat_i[30]
port 54 nsew signal input
rlabel metal3 s 523200 142128 524400 142248 6 hk_dat_i[31]
port 55 nsew signal input
rlabel metal3 s 523200 99968 524400 100088 6 hk_dat_i[3]
port 56 nsew signal input
rlabel metal3 s 523200 101464 524400 101584 6 hk_dat_i[4]
port 57 nsew signal input
rlabel metal3 s 523200 102960 524400 103080 6 hk_dat_i[5]
port 58 nsew signal input
rlabel metal3 s 523200 104456 524400 104576 6 hk_dat_i[6]
port 59 nsew signal input
rlabel metal3 s 523200 105952 524400 106072 6 hk_dat_i[7]
port 60 nsew signal input
rlabel metal3 s 523200 107448 524400 107568 6 hk_dat_i[8]
port 61 nsew signal input
rlabel metal3 s 523200 108944 524400 109064 6 hk_dat_i[9]
port 62 nsew signal input
rlabel metal3 s 523200 92352 524400 92472 6 hk_stb_o
port 63 nsew signal output
rlabel metal2 s 521842 163200 521898 164400 6 irq[0]
port 64 nsew signal input
rlabel metal2 s 522670 163200 522726 164400 6 irq[1]
port 65 nsew signal input
rlabel metal2 s 523498 163200 523554 164400 6 irq[2]
port 66 nsew signal input
rlabel metal3 s 523200 74400 524400 74520 6 irq[3]
port 67 nsew signal input
rlabel metal3 s 523200 72904 524400 73024 6 irq[4]
port 68 nsew signal input
rlabel metal3 s 523200 71408 524400 71528 6 irq[5]
port 69 nsew signal input
rlabel metal2 s 386 163200 442 164400 6 la_iena[0]
port 70 nsew signal output
rlabel metal2 s 336830 163200 336886 164400 6 la_iena[100]
port 71 nsew signal output
rlabel metal2 s 340142 163200 340198 164400 6 la_iena[101]
port 72 nsew signal output
rlabel metal2 s 343546 163200 343602 164400 6 la_iena[102]
port 73 nsew signal output
rlabel metal2 s 346858 163200 346914 164400 6 la_iena[103]
port 74 nsew signal output
rlabel metal2 s 350262 163200 350318 164400 6 la_iena[104]
port 75 nsew signal output
rlabel metal2 s 353666 163200 353722 164400 6 la_iena[105]
port 76 nsew signal output
rlabel metal2 s 356978 163200 357034 164400 6 la_iena[106]
port 77 nsew signal output
rlabel metal2 s 360382 163200 360438 164400 6 la_iena[107]
port 78 nsew signal output
rlabel metal2 s 363694 163200 363750 164400 6 la_iena[108]
port 79 nsew signal output
rlabel metal2 s 367098 163200 367154 164400 6 la_iena[109]
port 80 nsew signal output
rlabel metal2 s 33966 163200 34022 164400 6 la_iena[10]
port 81 nsew signal output
rlabel metal2 s 370410 163200 370466 164400 6 la_iena[110]
port 82 nsew signal output
rlabel metal2 s 373814 163200 373870 164400 6 la_iena[111]
port 83 nsew signal output
rlabel metal2 s 377218 163200 377274 164400 6 la_iena[112]
port 84 nsew signal output
rlabel metal2 s 380530 163200 380586 164400 6 la_iena[113]
port 85 nsew signal output
rlabel metal2 s 383934 163200 383990 164400 6 la_iena[114]
port 86 nsew signal output
rlabel metal2 s 387246 163200 387302 164400 6 la_iena[115]
port 87 nsew signal output
rlabel metal2 s 390650 163200 390706 164400 6 la_iena[116]
port 88 nsew signal output
rlabel metal2 s 393962 163200 394018 164400 6 la_iena[117]
port 89 nsew signal output
rlabel metal2 s 397366 163200 397422 164400 6 la_iena[118]
port 90 nsew signal output
rlabel metal2 s 400770 163200 400826 164400 6 la_iena[119]
port 91 nsew signal output
rlabel metal2 s 37370 163200 37426 164400 6 la_iena[11]
port 92 nsew signal output
rlabel metal2 s 404082 163200 404138 164400 6 la_iena[120]
port 93 nsew signal output
rlabel metal2 s 407486 163200 407542 164400 6 la_iena[121]
port 94 nsew signal output
rlabel metal2 s 410798 163200 410854 164400 6 la_iena[122]
port 95 nsew signal output
rlabel metal2 s 414202 163200 414258 164400 6 la_iena[123]
port 96 nsew signal output
rlabel metal2 s 417514 163200 417570 164400 6 la_iena[124]
port 97 nsew signal output
rlabel metal2 s 420918 163200 420974 164400 6 la_iena[125]
port 98 nsew signal output
rlabel metal2 s 424322 163200 424378 164400 6 la_iena[126]
port 99 nsew signal output
rlabel metal2 s 427634 163200 427690 164400 6 la_iena[127]
port 100 nsew signal output
rlabel metal2 s 40682 163200 40738 164400 6 la_iena[12]
port 101 nsew signal output
rlabel metal2 s 44086 163200 44142 164400 6 la_iena[13]
port 102 nsew signal output
rlabel metal2 s 47490 163200 47546 164400 6 la_iena[14]
port 103 nsew signal output
rlabel metal2 s 50802 163200 50858 164400 6 la_iena[15]
port 104 nsew signal output
rlabel metal2 s 54206 163200 54262 164400 6 la_iena[16]
port 105 nsew signal output
rlabel metal2 s 57518 163200 57574 164400 6 la_iena[17]
port 106 nsew signal output
rlabel metal2 s 60922 163200 60978 164400 6 la_iena[18]
port 107 nsew signal output
rlabel metal2 s 64234 163200 64290 164400 6 la_iena[19]
port 108 nsew signal output
rlabel metal2 s 3698 163200 3754 164400 6 la_iena[1]
port 109 nsew signal output
rlabel metal2 s 67638 163200 67694 164400 6 la_iena[20]
port 110 nsew signal output
rlabel metal2 s 71042 163200 71098 164400 6 la_iena[21]
port 111 nsew signal output
rlabel metal2 s 74354 163200 74410 164400 6 la_iena[22]
port 112 nsew signal output
rlabel metal2 s 77758 163200 77814 164400 6 la_iena[23]
port 113 nsew signal output
rlabel metal2 s 81070 163200 81126 164400 6 la_iena[24]
port 114 nsew signal output
rlabel metal2 s 84474 163200 84530 164400 6 la_iena[25]
port 115 nsew signal output
rlabel metal2 s 87786 163200 87842 164400 6 la_iena[26]
port 116 nsew signal output
rlabel metal2 s 91190 163200 91246 164400 6 la_iena[27]
port 117 nsew signal output
rlabel metal2 s 94594 163200 94650 164400 6 la_iena[28]
port 118 nsew signal output
rlabel metal2 s 97906 163200 97962 164400 6 la_iena[29]
port 119 nsew signal output
rlabel metal2 s 7102 163200 7158 164400 6 la_iena[2]
port 120 nsew signal output
rlabel metal2 s 101310 163200 101366 164400 6 la_iena[30]
port 121 nsew signal output
rlabel metal2 s 104622 163200 104678 164400 6 la_iena[31]
port 122 nsew signal output
rlabel metal2 s 108026 163200 108082 164400 6 la_iena[32]
port 123 nsew signal output
rlabel metal2 s 111338 163200 111394 164400 6 la_iena[33]
port 124 nsew signal output
rlabel metal2 s 114742 163200 114798 164400 6 la_iena[34]
port 125 nsew signal output
rlabel metal2 s 118146 163200 118202 164400 6 la_iena[35]
port 126 nsew signal output
rlabel metal2 s 121458 163200 121514 164400 6 la_iena[36]
port 127 nsew signal output
rlabel metal2 s 124862 163200 124918 164400 6 la_iena[37]
port 128 nsew signal output
rlabel metal2 s 128174 163200 128230 164400 6 la_iena[38]
port 129 nsew signal output
rlabel metal2 s 131578 163200 131634 164400 6 la_iena[39]
port 130 nsew signal output
rlabel metal2 s 10414 163200 10470 164400 6 la_iena[3]
port 131 nsew signal output
rlabel metal2 s 134890 163200 134946 164400 6 la_iena[40]
port 132 nsew signal output
rlabel metal2 s 138294 163200 138350 164400 6 la_iena[41]
port 133 nsew signal output
rlabel metal2 s 141698 163200 141754 164400 6 la_iena[42]
port 134 nsew signal output
rlabel metal2 s 145010 163200 145066 164400 6 la_iena[43]
port 135 nsew signal output
rlabel metal2 s 148414 163200 148470 164400 6 la_iena[44]
port 136 nsew signal output
rlabel metal2 s 151726 163200 151782 164400 6 la_iena[45]
port 137 nsew signal output
rlabel metal2 s 155130 163200 155186 164400 6 la_iena[46]
port 138 nsew signal output
rlabel metal2 s 158442 163200 158498 164400 6 la_iena[47]
port 139 nsew signal output
rlabel metal2 s 161846 163200 161902 164400 6 la_iena[48]
port 140 nsew signal output
rlabel metal2 s 165250 163200 165306 164400 6 la_iena[49]
port 141 nsew signal output
rlabel metal2 s 13818 163200 13874 164400 6 la_iena[4]
port 142 nsew signal output
rlabel metal2 s 168562 163200 168618 164400 6 la_iena[50]
port 143 nsew signal output
rlabel metal2 s 171966 163200 172022 164400 6 la_iena[51]
port 144 nsew signal output
rlabel metal2 s 175278 163200 175334 164400 6 la_iena[52]
port 145 nsew signal output
rlabel metal2 s 178682 163200 178738 164400 6 la_iena[53]
port 146 nsew signal output
rlabel metal2 s 181994 163200 182050 164400 6 la_iena[54]
port 147 nsew signal output
rlabel metal2 s 185398 163200 185454 164400 6 la_iena[55]
port 148 nsew signal output
rlabel metal2 s 188802 163200 188858 164400 6 la_iena[56]
port 149 nsew signal output
rlabel metal2 s 192114 163200 192170 164400 6 la_iena[57]
port 150 nsew signal output
rlabel metal2 s 195518 163200 195574 164400 6 la_iena[58]
port 151 nsew signal output
rlabel metal2 s 198830 163200 198886 164400 6 la_iena[59]
port 152 nsew signal output
rlabel metal2 s 17130 163200 17186 164400 6 la_iena[5]
port 153 nsew signal output
rlabel metal2 s 202234 163200 202290 164400 6 la_iena[60]
port 154 nsew signal output
rlabel metal2 s 205546 163200 205602 164400 6 la_iena[61]
port 155 nsew signal output
rlabel metal2 s 208950 163200 209006 164400 6 la_iena[62]
port 156 nsew signal output
rlabel metal2 s 212354 163200 212410 164400 6 la_iena[63]
port 157 nsew signal output
rlabel metal2 s 215666 163200 215722 164400 6 la_iena[64]
port 158 nsew signal output
rlabel metal2 s 219070 163200 219126 164400 6 la_iena[65]
port 159 nsew signal output
rlabel metal2 s 222382 163200 222438 164400 6 la_iena[66]
port 160 nsew signal output
rlabel metal2 s 225786 163200 225842 164400 6 la_iena[67]
port 161 nsew signal output
rlabel metal2 s 229098 163200 229154 164400 6 la_iena[68]
port 162 nsew signal output
rlabel metal2 s 232502 163200 232558 164400 6 la_iena[69]
port 163 nsew signal output
rlabel metal2 s 20534 163200 20590 164400 6 la_iena[6]
port 164 nsew signal output
rlabel metal2 s 235906 163200 235962 164400 6 la_iena[70]
port 165 nsew signal output
rlabel metal2 s 239218 163200 239274 164400 6 la_iena[71]
port 166 nsew signal output
rlabel metal2 s 242622 163200 242678 164400 6 la_iena[72]
port 167 nsew signal output
rlabel metal2 s 245934 163200 245990 164400 6 la_iena[73]
port 168 nsew signal output
rlabel metal2 s 249338 163200 249394 164400 6 la_iena[74]
port 169 nsew signal output
rlabel metal2 s 252650 163200 252706 164400 6 la_iena[75]
port 170 nsew signal output
rlabel metal2 s 256054 163200 256110 164400 6 la_iena[76]
port 171 nsew signal output
rlabel metal2 s 259458 163200 259514 164400 6 la_iena[77]
port 172 nsew signal output
rlabel metal2 s 262770 163200 262826 164400 6 la_iena[78]
port 173 nsew signal output
rlabel metal2 s 266174 163200 266230 164400 6 la_iena[79]
port 174 nsew signal output
rlabel metal2 s 23938 163200 23994 164400 6 la_iena[7]
port 175 nsew signal output
rlabel metal2 s 269486 163200 269542 164400 6 la_iena[80]
port 176 nsew signal output
rlabel metal2 s 272890 163200 272946 164400 6 la_iena[81]
port 177 nsew signal output
rlabel metal2 s 276202 163200 276258 164400 6 la_iena[82]
port 178 nsew signal output
rlabel metal2 s 279606 163200 279662 164400 6 la_iena[83]
port 179 nsew signal output
rlabel metal2 s 283010 163200 283066 164400 6 la_iena[84]
port 180 nsew signal output
rlabel metal2 s 286322 163200 286378 164400 6 la_iena[85]
port 181 nsew signal output
rlabel metal2 s 289726 163200 289782 164400 6 la_iena[86]
port 182 nsew signal output
rlabel metal2 s 293038 163200 293094 164400 6 la_iena[87]
port 183 nsew signal output
rlabel metal2 s 296442 163200 296498 164400 6 la_iena[88]
port 184 nsew signal output
rlabel metal2 s 299754 163200 299810 164400 6 la_iena[89]
port 185 nsew signal output
rlabel metal2 s 27250 163200 27306 164400 6 la_iena[8]
port 186 nsew signal output
rlabel metal2 s 303158 163200 303214 164400 6 la_iena[90]
port 187 nsew signal output
rlabel metal2 s 306562 163200 306618 164400 6 la_iena[91]
port 188 nsew signal output
rlabel metal2 s 309874 163200 309930 164400 6 la_iena[92]
port 189 nsew signal output
rlabel metal2 s 313278 163200 313334 164400 6 la_iena[93]
port 190 nsew signal output
rlabel metal2 s 316590 163200 316646 164400 6 la_iena[94]
port 191 nsew signal output
rlabel metal2 s 319994 163200 320050 164400 6 la_iena[95]
port 192 nsew signal output
rlabel metal2 s 323306 163200 323362 164400 6 la_iena[96]
port 193 nsew signal output
rlabel metal2 s 326710 163200 326766 164400 6 la_iena[97]
port 194 nsew signal output
rlabel metal2 s 330114 163200 330170 164400 6 la_iena[98]
port 195 nsew signal output
rlabel metal2 s 333426 163200 333482 164400 6 la_iena[99]
port 196 nsew signal output
rlabel metal2 s 30654 163200 30710 164400 6 la_iena[9]
port 197 nsew signal output
rlabel metal2 s 1214 163200 1270 164400 6 la_input[0]
port 198 nsew signal input
rlabel metal2 s 337658 163200 337714 164400 6 la_input[100]
port 199 nsew signal input
rlabel metal2 s 340970 163200 341026 164400 6 la_input[101]
port 200 nsew signal input
rlabel metal2 s 344374 163200 344430 164400 6 la_input[102]
port 201 nsew signal input
rlabel metal2 s 347778 163200 347834 164400 6 la_input[103]
port 202 nsew signal input
rlabel metal2 s 351090 163200 351146 164400 6 la_input[104]
port 203 nsew signal input
rlabel metal2 s 354494 163200 354550 164400 6 la_input[105]
port 204 nsew signal input
rlabel metal2 s 357806 163200 357862 164400 6 la_input[106]
port 205 nsew signal input
rlabel metal2 s 361210 163200 361266 164400 6 la_input[107]
port 206 nsew signal input
rlabel metal2 s 364522 163200 364578 164400 6 la_input[108]
port 207 nsew signal input
rlabel metal2 s 367926 163200 367982 164400 6 la_input[109]
port 208 nsew signal input
rlabel metal2 s 34794 163200 34850 164400 6 la_input[10]
port 209 nsew signal input
rlabel metal2 s 371330 163200 371386 164400 6 la_input[110]
port 210 nsew signal input
rlabel metal2 s 374642 163200 374698 164400 6 la_input[111]
port 211 nsew signal input
rlabel metal2 s 378046 163200 378102 164400 6 la_input[112]
port 212 nsew signal input
rlabel metal2 s 381358 163200 381414 164400 6 la_input[113]
port 213 nsew signal input
rlabel metal2 s 384762 163200 384818 164400 6 la_input[114]
port 214 nsew signal input
rlabel metal2 s 388074 163200 388130 164400 6 la_input[115]
port 215 nsew signal input
rlabel metal2 s 391478 163200 391534 164400 6 la_input[116]
port 216 nsew signal input
rlabel metal2 s 394882 163200 394938 164400 6 la_input[117]
port 217 nsew signal input
rlabel metal2 s 398194 163200 398250 164400 6 la_input[118]
port 218 nsew signal input
rlabel metal2 s 401598 163200 401654 164400 6 la_input[119]
port 219 nsew signal input
rlabel metal2 s 38198 163200 38254 164400 6 la_input[11]
port 220 nsew signal input
rlabel metal2 s 404910 163200 404966 164400 6 la_input[120]
port 221 nsew signal input
rlabel metal2 s 408314 163200 408370 164400 6 la_input[121]
port 222 nsew signal input
rlabel metal2 s 411626 163200 411682 164400 6 la_input[122]
port 223 nsew signal input
rlabel metal2 s 415030 163200 415086 164400 6 la_input[123]
port 224 nsew signal input
rlabel metal2 s 418434 163200 418490 164400 6 la_input[124]
port 225 nsew signal input
rlabel metal2 s 421746 163200 421802 164400 6 la_input[125]
port 226 nsew signal input
rlabel metal2 s 425150 163200 425206 164400 6 la_input[126]
port 227 nsew signal input
rlabel metal2 s 428462 163200 428518 164400 6 la_input[127]
port 228 nsew signal input
rlabel metal2 s 41602 163200 41658 164400 6 la_input[12]
port 229 nsew signal input
rlabel metal2 s 44914 163200 44970 164400 6 la_input[13]
port 230 nsew signal input
rlabel metal2 s 48318 163200 48374 164400 6 la_input[14]
port 231 nsew signal input
rlabel metal2 s 51630 163200 51686 164400 6 la_input[15]
port 232 nsew signal input
rlabel metal2 s 55034 163200 55090 164400 6 la_input[16]
port 233 nsew signal input
rlabel metal2 s 58346 163200 58402 164400 6 la_input[17]
port 234 nsew signal input
rlabel metal2 s 61750 163200 61806 164400 6 la_input[18]
port 235 nsew signal input
rlabel metal2 s 65154 163200 65210 164400 6 la_input[19]
port 236 nsew signal input
rlabel metal2 s 4526 163200 4582 164400 6 la_input[1]
port 237 nsew signal input
rlabel metal2 s 68466 163200 68522 164400 6 la_input[20]
port 238 nsew signal input
rlabel metal2 s 71870 163200 71926 164400 6 la_input[21]
port 239 nsew signal input
rlabel metal2 s 75182 163200 75238 164400 6 la_input[22]
port 240 nsew signal input
rlabel metal2 s 78586 163200 78642 164400 6 la_input[23]
port 241 nsew signal input
rlabel metal2 s 81898 163200 81954 164400 6 la_input[24]
port 242 nsew signal input
rlabel metal2 s 85302 163200 85358 164400 6 la_input[25]
port 243 nsew signal input
rlabel metal2 s 88706 163200 88762 164400 6 la_input[26]
port 244 nsew signal input
rlabel metal2 s 92018 163200 92074 164400 6 la_input[27]
port 245 nsew signal input
rlabel metal2 s 95422 163200 95478 164400 6 la_input[28]
port 246 nsew signal input
rlabel metal2 s 98734 163200 98790 164400 6 la_input[29]
port 247 nsew signal input
rlabel metal2 s 7930 163200 7986 164400 6 la_input[2]
port 248 nsew signal input
rlabel metal2 s 102138 163200 102194 164400 6 la_input[30]
port 249 nsew signal input
rlabel metal2 s 105450 163200 105506 164400 6 la_input[31]
port 250 nsew signal input
rlabel metal2 s 108854 163200 108910 164400 6 la_input[32]
port 251 nsew signal input
rlabel metal2 s 112258 163200 112314 164400 6 la_input[33]
port 252 nsew signal input
rlabel metal2 s 115570 163200 115626 164400 6 la_input[34]
port 253 nsew signal input
rlabel metal2 s 118974 163200 119030 164400 6 la_input[35]
port 254 nsew signal input
rlabel metal2 s 122286 163200 122342 164400 6 la_input[36]
port 255 nsew signal input
rlabel metal2 s 125690 163200 125746 164400 6 la_input[37]
port 256 nsew signal input
rlabel metal2 s 129002 163200 129058 164400 6 la_input[38]
port 257 nsew signal input
rlabel metal2 s 132406 163200 132462 164400 6 la_input[39]
port 258 nsew signal input
rlabel metal2 s 11242 163200 11298 164400 6 la_input[3]
port 259 nsew signal input
rlabel metal2 s 135810 163200 135866 164400 6 la_input[40]
port 260 nsew signal input
rlabel metal2 s 139122 163200 139178 164400 6 la_input[41]
port 261 nsew signal input
rlabel metal2 s 142526 163200 142582 164400 6 la_input[42]
port 262 nsew signal input
rlabel metal2 s 145838 163200 145894 164400 6 la_input[43]
port 263 nsew signal input
rlabel metal2 s 149242 163200 149298 164400 6 la_input[44]
port 264 nsew signal input
rlabel metal2 s 152554 163200 152610 164400 6 la_input[45]
port 265 nsew signal input
rlabel metal2 s 155958 163200 156014 164400 6 la_input[46]
port 266 nsew signal input
rlabel metal2 s 159362 163200 159418 164400 6 la_input[47]
port 267 nsew signal input
rlabel metal2 s 162674 163200 162730 164400 6 la_input[48]
port 268 nsew signal input
rlabel metal2 s 166078 163200 166134 164400 6 la_input[49]
port 269 nsew signal input
rlabel metal2 s 14646 163200 14702 164400 6 la_input[4]
port 270 nsew signal input
rlabel metal2 s 169390 163200 169446 164400 6 la_input[50]
port 271 nsew signal input
rlabel metal2 s 172794 163200 172850 164400 6 la_input[51]
port 272 nsew signal input
rlabel metal2 s 176106 163200 176162 164400 6 la_input[52]
port 273 nsew signal input
rlabel metal2 s 179510 163200 179566 164400 6 la_input[53]
port 274 nsew signal input
rlabel metal2 s 182914 163200 182970 164400 6 la_input[54]
port 275 nsew signal input
rlabel metal2 s 186226 163200 186282 164400 6 la_input[55]
port 276 nsew signal input
rlabel metal2 s 189630 163200 189686 164400 6 la_input[56]
port 277 nsew signal input
rlabel metal2 s 192942 163200 192998 164400 6 la_input[57]
port 278 nsew signal input
rlabel metal2 s 196346 163200 196402 164400 6 la_input[58]
port 279 nsew signal input
rlabel metal2 s 199658 163200 199714 164400 6 la_input[59]
port 280 nsew signal input
rlabel metal2 s 18050 163200 18106 164400 6 la_input[5]
port 281 nsew signal input
rlabel metal2 s 203062 163200 203118 164400 6 la_input[60]
port 282 nsew signal input
rlabel metal2 s 206466 163200 206522 164400 6 la_input[61]
port 283 nsew signal input
rlabel metal2 s 209778 163200 209834 164400 6 la_input[62]
port 284 nsew signal input
rlabel metal2 s 213182 163200 213238 164400 6 la_input[63]
port 285 nsew signal input
rlabel metal2 s 216494 163200 216550 164400 6 la_input[64]
port 286 nsew signal input
rlabel metal2 s 219898 163200 219954 164400 6 la_input[65]
port 287 nsew signal input
rlabel metal2 s 223210 163200 223266 164400 6 la_input[66]
port 288 nsew signal input
rlabel metal2 s 226614 163200 226670 164400 6 la_input[67]
port 289 nsew signal input
rlabel metal2 s 230018 163200 230074 164400 6 la_input[68]
port 290 nsew signal input
rlabel metal2 s 233330 163200 233386 164400 6 la_input[69]
port 291 nsew signal input
rlabel metal2 s 21362 163200 21418 164400 6 la_input[6]
port 292 nsew signal input
rlabel metal2 s 236734 163200 236790 164400 6 la_input[70]
port 293 nsew signal input
rlabel metal2 s 240046 163200 240102 164400 6 la_input[71]
port 294 nsew signal input
rlabel metal2 s 243450 163200 243506 164400 6 la_input[72]
port 295 nsew signal input
rlabel metal2 s 246762 163200 246818 164400 6 la_input[73]
port 296 nsew signal input
rlabel metal2 s 250166 163200 250222 164400 6 la_input[74]
port 297 nsew signal input
rlabel metal2 s 253570 163200 253626 164400 6 la_input[75]
port 298 nsew signal input
rlabel metal2 s 256882 163200 256938 164400 6 la_input[76]
port 299 nsew signal input
rlabel metal2 s 260286 163200 260342 164400 6 la_input[77]
port 300 nsew signal input
rlabel metal2 s 263598 163200 263654 164400 6 la_input[78]
port 301 nsew signal input
rlabel metal2 s 267002 163200 267058 164400 6 la_input[79]
port 302 nsew signal input
rlabel metal2 s 24766 163200 24822 164400 6 la_input[7]
port 303 nsew signal input
rlabel metal2 s 270314 163200 270370 164400 6 la_input[80]
port 304 nsew signal input
rlabel metal2 s 273718 163200 273774 164400 6 la_input[81]
port 305 nsew signal input
rlabel metal2 s 277122 163200 277178 164400 6 la_input[82]
port 306 nsew signal input
rlabel metal2 s 280434 163200 280490 164400 6 la_input[83]
port 307 nsew signal input
rlabel metal2 s 283838 163200 283894 164400 6 la_input[84]
port 308 nsew signal input
rlabel metal2 s 287150 163200 287206 164400 6 la_input[85]
port 309 nsew signal input
rlabel metal2 s 290554 163200 290610 164400 6 la_input[86]
port 310 nsew signal input
rlabel metal2 s 293866 163200 293922 164400 6 la_input[87]
port 311 nsew signal input
rlabel metal2 s 297270 163200 297326 164400 6 la_input[88]
port 312 nsew signal input
rlabel metal2 s 300674 163200 300730 164400 6 la_input[89]
port 313 nsew signal input
rlabel metal2 s 28078 163200 28134 164400 6 la_input[8]
port 314 nsew signal input
rlabel metal2 s 303986 163200 304042 164400 6 la_input[90]
port 315 nsew signal input
rlabel metal2 s 307390 163200 307446 164400 6 la_input[91]
port 316 nsew signal input
rlabel metal2 s 310702 163200 310758 164400 6 la_input[92]
port 317 nsew signal input
rlabel metal2 s 314106 163200 314162 164400 6 la_input[93]
port 318 nsew signal input
rlabel metal2 s 317418 163200 317474 164400 6 la_input[94]
port 319 nsew signal input
rlabel metal2 s 320822 163200 320878 164400 6 la_input[95]
port 320 nsew signal input
rlabel metal2 s 324226 163200 324282 164400 6 la_input[96]
port 321 nsew signal input
rlabel metal2 s 327538 163200 327594 164400 6 la_input[97]
port 322 nsew signal input
rlabel metal2 s 330942 163200 330998 164400 6 la_input[98]
port 323 nsew signal input
rlabel metal2 s 334254 163200 334310 164400 6 la_input[99]
port 324 nsew signal input
rlabel metal2 s 31482 163200 31538 164400 6 la_input[9]
port 325 nsew signal input
rlabel metal2 s 2042 163200 2098 164400 6 la_oenb[0]
port 326 nsew signal output
rlabel metal2 s 338486 163200 338542 164400 6 la_oenb[100]
port 327 nsew signal output
rlabel metal2 s 341890 163200 341946 164400 6 la_oenb[101]
port 328 nsew signal output
rlabel metal2 s 345202 163200 345258 164400 6 la_oenb[102]
port 329 nsew signal output
rlabel metal2 s 348606 163200 348662 164400 6 la_oenb[103]
port 330 nsew signal output
rlabel metal2 s 351918 163200 351974 164400 6 la_oenb[104]
port 331 nsew signal output
rlabel metal2 s 355322 163200 355378 164400 6 la_oenb[105]
port 332 nsew signal output
rlabel metal2 s 358634 163200 358690 164400 6 la_oenb[106]
port 333 nsew signal output
rlabel metal2 s 362038 163200 362094 164400 6 la_oenb[107]
port 334 nsew signal output
rlabel metal2 s 365442 163200 365498 164400 6 la_oenb[108]
port 335 nsew signal output
rlabel metal2 s 368754 163200 368810 164400 6 la_oenb[109]
port 336 nsew signal output
rlabel metal2 s 35714 163200 35770 164400 6 la_oenb[10]
port 337 nsew signal output
rlabel metal2 s 372158 163200 372214 164400 6 la_oenb[110]
port 338 nsew signal output
rlabel metal2 s 375470 163200 375526 164400 6 la_oenb[111]
port 339 nsew signal output
rlabel metal2 s 378874 163200 378930 164400 6 la_oenb[112]
port 340 nsew signal output
rlabel metal2 s 382186 163200 382242 164400 6 la_oenb[113]
port 341 nsew signal output
rlabel metal2 s 385590 163200 385646 164400 6 la_oenb[114]
port 342 nsew signal output
rlabel metal2 s 388994 163200 389050 164400 6 la_oenb[115]
port 343 nsew signal output
rlabel metal2 s 392306 163200 392362 164400 6 la_oenb[116]
port 344 nsew signal output
rlabel metal2 s 395710 163200 395766 164400 6 la_oenb[117]
port 345 nsew signal output
rlabel metal2 s 399022 163200 399078 164400 6 la_oenb[118]
port 346 nsew signal output
rlabel metal2 s 402426 163200 402482 164400 6 la_oenb[119]
port 347 nsew signal output
rlabel metal2 s 39026 163200 39082 164400 6 la_oenb[11]
port 348 nsew signal output
rlabel metal2 s 405738 163200 405794 164400 6 la_oenb[120]
port 349 nsew signal output
rlabel metal2 s 409142 163200 409198 164400 6 la_oenb[121]
port 350 nsew signal output
rlabel metal2 s 412546 163200 412602 164400 6 la_oenb[122]
port 351 nsew signal output
rlabel metal2 s 415858 163200 415914 164400 6 la_oenb[123]
port 352 nsew signal output
rlabel metal2 s 419262 163200 419318 164400 6 la_oenb[124]
port 353 nsew signal output
rlabel metal2 s 422574 163200 422630 164400 6 la_oenb[125]
port 354 nsew signal output
rlabel metal2 s 425978 163200 426034 164400 6 la_oenb[126]
port 355 nsew signal output
rlabel metal2 s 429290 163200 429346 164400 6 la_oenb[127]
port 356 nsew signal output
rlabel metal2 s 42430 163200 42486 164400 6 la_oenb[12]
port 357 nsew signal output
rlabel metal2 s 45742 163200 45798 164400 6 la_oenb[13]
port 358 nsew signal output
rlabel metal2 s 49146 163200 49202 164400 6 la_oenb[14]
port 359 nsew signal output
rlabel metal2 s 52458 163200 52514 164400 6 la_oenb[15]
port 360 nsew signal output
rlabel metal2 s 55862 163200 55918 164400 6 la_oenb[16]
port 361 nsew signal output
rlabel metal2 s 59266 163200 59322 164400 6 la_oenb[17]
port 362 nsew signal output
rlabel metal2 s 62578 163200 62634 164400 6 la_oenb[18]
port 363 nsew signal output
rlabel metal2 s 65982 163200 66038 164400 6 la_oenb[19]
port 364 nsew signal output
rlabel metal2 s 5354 163200 5410 164400 6 la_oenb[1]
port 365 nsew signal output
rlabel metal2 s 69294 163200 69350 164400 6 la_oenb[20]
port 366 nsew signal output
rlabel metal2 s 72698 163200 72754 164400 6 la_oenb[21]
port 367 nsew signal output
rlabel metal2 s 76010 163200 76066 164400 6 la_oenb[22]
port 368 nsew signal output
rlabel metal2 s 79414 163200 79470 164400 6 la_oenb[23]
port 369 nsew signal output
rlabel metal2 s 82818 163200 82874 164400 6 la_oenb[24]
port 370 nsew signal output
rlabel metal2 s 86130 163200 86186 164400 6 la_oenb[25]
port 371 nsew signal output
rlabel metal2 s 89534 163200 89590 164400 6 la_oenb[26]
port 372 nsew signal output
rlabel metal2 s 92846 163200 92902 164400 6 la_oenb[27]
port 373 nsew signal output
rlabel metal2 s 96250 163200 96306 164400 6 la_oenb[28]
port 374 nsew signal output
rlabel metal2 s 99562 163200 99618 164400 6 la_oenb[29]
port 375 nsew signal output
rlabel metal2 s 8758 163200 8814 164400 6 la_oenb[2]
port 376 nsew signal output
rlabel metal2 s 102966 163200 103022 164400 6 la_oenb[30]
port 377 nsew signal output
rlabel metal2 s 106370 163200 106426 164400 6 la_oenb[31]
port 378 nsew signal output
rlabel metal2 s 109682 163200 109738 164400 6 la_oenb[32]
port 379 nsew signal output
rlabel metal2 s 113086 163200 113142 164400 6 la_oenb[33]
port 380 nsew signal output
rlabel metal2 s 116398 163200 116454 164400 6 la_oenb[34]
port 381 nsew signal output
rlabel metal2 s 119802 163200 119858 164400 6 la_oenb[35]
port 382 nsew signal output
rlabel metal2 s 123114 163200 123170 164400 6 la_oenb[36]
port 383 nsew signal output
rlabel metal2 s 126518 163200 126574 164400 6 la_oenb[37]
port 384 nsew signal output
rlabel metal2 s 129922 163200 129978 164400 6 la_oenb[38]
port 385 nsew signal output
rlabel metal2 s 133234 163200 133290 164400 6 la_oenb[39]
port 386 nsew signal output
rlabel metal2 s 12162 163200 12218 164400 6 la_oenb[3]
port 387 nsew signal output
rlabel metal2 s 136638 163200 136694 164400 6 la_oenb[40]
port 388 nsew signal output
rlabel metal2 s 139950 163200 140006 164400 6 la_oenb[41]
port 389 nsew signal output
rlabel metal2 s 143354 163200 143410 164400 6 la_oenb[42]
port 390 nsew signal output
rlabel metal2 s 146666 163200 146722 164400 6 la_oenb[43]
port 391 nsew signal output
rlabel metal2 s 150070 163200 150126 164400 6 la_oenb[44]
port 392 nsew signal output
rlabel metal2 s 153474 163200 153530 164400 6 la_oenb[45]
port 393 nsew signal output
rlabel metal2 s 156786 163200 156842 164400 6 la_oenb[46]
port 394 nsew signal output
rlabel metal2 s 160190 163200 160246 164400 6 la_oenb[47]
port 395 nsew signal output
rlabel metal2 s 163502 163200 163558 164400 6 la_oenb[48]
port 396 nsew signal output
rlabel metal2 s 166906 163200 166962 164400 6 la_oenb[49]
port 397 nsew signal output
rlabel metal2 s 15474 163200 15530 164400 6 la_oenb[4]
port 398 nsew signal output
rlabel metal2 s 170218 163200 170274 164400 6 la_oenb[50]
port 399 nsew signal output
rlabel metal2 s 173622 163200 173678 164400 6 la_oenb[51]
port 400 nsew signal output
rlabel metal2 s 177026 163200 177082 164400 6 la_oenb[52]
port 401 nsew signal output
rlabel metal2 s 180338 163200 180394 164400 6 la_oenb[53]
port 402 nsew signal output
rlabel metal2 s 183742 163200 183798 164400 6 la_oenb[54]
port 403 nsew signal output
rlabel metal2 s 187054 163200 187110 164400 6 la_oenb[55]
port 404 nsew signal output
rlabel metal2 s 190458 163200 190514 164400 6 la_oenb[56]
port 405 nsew signal output
rlabel metal2 s 193770 163200 193826 164400 6 la_oenb[57]
port 406 nsew signal output
rlabel metal2 s 197174 163200 197230 164400 6 la_oenb[58]
port 407 nsew signal output
rlabel metal2 s 200578 163200 200634 164400 6 la_oenb[59]
port 408 nsew signal output
rlabel metal2 s 18878 163200 18934 164400 6 la_oenb[5]
port 409 nsew signal output
rlabel metal2 s 203890 163200 203946 164400 6 la_oenb[60]
port 410 nsew signal output
rlabel metal2 s 207294 163200 207350 164400 6 la_oenb[61]
port 411 nsew signal output
rlabel metal2 s 210606 163200 210662 164400 6 la_oenb[62]
port 412 nsew signal output
rlabel metal2 s 214010 163200 214066 164400 6 la_oenb[63]
port 413 nsew signal output
rlabel metal2 s 217322 163200 217378 164400 6 la_oenb[64]
port 414 nsew signal output
rlabel metal2 s 220726 163200 220782 164400 6 la_oenb[65]
port 415 nsew signal output
rlabel metal2 s 224130 163200 224186 164400 6 la_oenb[66]
port 416 nsew signal output
rlabel metal2 s 227442 163200 227498 164400 6 la_oenb[67]
port 417 nsew signal output
rlabel metal2 s 230846 163200 230902 164400 6 la_oenb[68]
port 418 nsew signal output
rlabel metal2 s 234158 163200 234214 164400 6 la_oenb[69]
port 419 nsew signal output
rlabel metal2 s 22190 163200 22246 164400 6 la_oenb[6]
port 420 nsew signal output
rlabel metal2 s 237562 163200 237618 164400 6 la_oenb[70]
port 421 nsew signal output
rlabel metal2 s 240874 163200 240930 164400 6 la_oenb[71]
port 422 nsew signal output
rlabel metal2 s 244278 163200 244334 164400 6 la_oenb[72]
port 423 nsew signal output
rlabel metal2 s 247682 163200 247738 164400 6 la_oenb[73]
port 424 nsew signal output
rlabel metal2 s 250994 163200 251050 164400 6 la_oenb[74]
port 425 nsew signal output
rlabel metal2 s 254398 163200 254454 164400 6 la_oenb[75]
port 426 nsew signal output
rlabel metal2 s 257710 163200 257766 164400 6 la_oenb[76]
port 427 nsew signal output
rlabel metal2 s 261114 163200 261170 164400 6 la_oenb[77]
port 428 nsew signal output
rlabel metal2 s 264426 163200 264482 164400 6 la_oenb[78]
port 429 nsew signal output
rlabel metal2 s 267830 163200 267886 164400 6 la_oenb[79]
port 430 nsew signal output
rlabel metal2 s 25594 163200 25650 164400 6 la_oenb[7]
port 431 nsew signal output
rlabel metal2 s 271234 163200 271290 164400 6 la_oenb[80]
port 432 nsew signal output
rlabel metal2 s 274546 163200 274602 164400 6 la_oenb[81]
port 433 nsew signal output
rlabel metal2 s 277950 163200 278006 164400 6 la_oenb[82]
port 434 nsew signal output
rlabel metal2 s 281262 163200 281318 164400 6 la_oenb[83]
port 435 nsew signal output
rlabel metal2 s 284666 163200 284722 164400 6 la_oenb[84]
port 436 nsew signal output
rlabel metal2 s 287978 163200 288034 164400 6 la_oenb[85]
port 437 nsew signal output
rlabel metal2 s 291382 163200 291438 164400 6 la_oenb[86]
port 438 nsew signal output
rlabel metal2 s 294786 163200 294842 164400 6 la_oenb[87]
port 439 nsew signal output
rlabel metal2 s 298098 163200 298154 164400 6 la_oenb[88]
port 440 nsew signal output
rlabel metal2 s 301502 163200 301558 164400 6 la_oenb[89]
port 441 nsew signal output
rlabel metal2 s 28906 163200 28962 164400 6 la_oenb[8]
port 442 nsew signal output
rlabel metal2 s 304814 163200 304870 164400 6 la_oenb[90]
port 443 nsew signal output
rlabel metal2 s 308218 163200 308274 164400 6 la_oenb[91]
port 444 nsew signal output
rlabel metal2 s 311530 163200 311586 164400 6 la_oenb[92]
port 445 nsew signal output
rlabel metal2 s 314934 163200 314990 164400 6 la_oenb[93]
port 446 nsew signal output
rlabel metal2 s 318338 163200 318394 164400 6 la_oenb[94]
port 447 nsew signal output
rlabel metal2 s 321650 163200 321706 164400 6 la_oenb[95]
port 448 nsew signal output
rlabel metal2 s 325054 163200 325110 164400 6 la_oenb[96]
port 449 nsew signal output
rlabel metal2 s 328366 163200 328422 164400 6 la_oenb[97]
port 450 nsew signal output
rlabel metal2 s 331770 163200 331826 164400 6 la_oenb[98]
port 451 nsew signal output
rlabel metal2 s 335082 163200 335138 164400 6 la_oenb[99]
port 452 nsew signal output
rlabel metal2 s 32310 163200 32366 164400 6 la_oenb[9]
port 453 nsew signal output
rlabel metal2 s 2870 163200 2926 164400 6 la_output[0]
port 454 nsew signal output
rlabel metal2 s 339314 163200 339370 164400 6 la_output[100]
port 455 nsew signal output
rlabel metal2 s 342718 163200 342774 164400 6 la_output[101]
port 456 nsew signal output
rlabel metal2 s 346030 163200 346086 164400 6 la_output[102]
port 457 nsew signal output
rlabel metal2 s 349434 163200 349490 164400 6 la_output[103]
port 458 nsew signal output
rlabel metal2 s 352746 163200 352802 164400 6 la_output[104]
port 459 nsew signal output
rlabel metal2 s 356150 163200 356206 164400 6 la_output[105]
port 460 nsew signal output
rlabel metal2 s 359554 163200 359610 164400 6 la_output[106]
port 461 nsew signal output
rlabel metal2 s 362866 163200 362922 164400 6 la_output[107]
port 462 nsew signal output
rlabel metal2 s 366270 163200 366326 164400 6 la_output[108]
port 463 nsew signal output
rlabel metal2 s 369582 163200 369638 164400 6 la_output[109]
port 464 nsew signal output
rlabel metal2 s 36542 163200 36598 164400 6 la_output[10]
port 465 nsew signal output
rlabel metal2 s 372986 163200 373042 164400 6 la_output[110]
port 466 nsew signal output
rlabel metal2 s 376298 163200 376354 164400 6 la_output[111]
port 467 nsew signal output
rlabel metal2 s 379702 163200 379758 164400 6 la_output[112]
port 468 nsew signal output
rlabel metal2 s 383106 163200 383162 164400 6 la_output[113]
port 469 nsew signal output
rlabel metal2 s 386418 163200 386474 164400 6 la_output[114]
port 470 nsew signal output
rlabel metal2 s 389822 163200 389878 164400 6 la_output[115]
port 471 nsew signal output
rlabel metal2 s 393134 163200 393190 164400 6 la_output[116]
port 472 nsew signal output
rlabel metal2 s 396538 163200 396594 164400 6 la_output[117]
port 473 nsew signal output
rlabel metal2 s 399850 163200 399906 164400 6 la_output[118]
port 474 nsew signal output
rlabel metal2 s 403254 163200 403310 164400 6 la_output[119]
port 475 nsew signal output
rlabel metal2 s 39854 163200 39910 164400 6 la_output[11]
port 476 nsew signal output
rlabel metal2 s 406658 163200 406714 164400 6 la_output[120]
port 477 nsew signal output
rlabel metal2 s 409970 163200 410026 164400 6 la_output[121]
port 478 nsew signal output
rlabel metal2 s 413374 163200 413430 164400 6 la_output[122]
port 479 nsew signal output
rlabel metal2 s 416686 163200 416742 164400 6 la_output[123]
port 480 nsew signal output
rlabel metal2 s 420090 163200 420146 164400 6 la_output[124]
port 481 nsew signal output
rlabel metal2 s 423402 163200 423458 164400 6 la_output[125]
port 482 nsew signal output
rlabel metal2 s 426806 163200 426862 164400 6 la_output[126]
port 483 nsew signal output
rlabel metal2 s 430210 163200 430266 164400 6 la_output[127]
port 484 nsew signal output
rlabel metal2 s 43258 163200 43314 164400 6 la_output[12]
port 485 nsew signal output
rlabel metal2 s 46570 163200 46626 164400 6 la_output[13]
port 486 nsew signal output
rlabel metal2 s 49974 163200 50030 164400 6 la_output[14]
port 487 nsew signal output
rlabel metal2 s 53378 163200 53434 164400 6 la_output[15]
port 488 nsew signal output
rlabel metal2 s 56690 163200 56746 164400 6 la_output[16]
port 489 nsew signal output
rlabel metal2 s 60094 163200 60150 164400 6 la_output[17]
port 490 nsew signal output
rlabel metal2 s 63406 163200 63462 164400 6 la_output[18]
port 491 nsew signal output
rlabel metal2 s 66810 163200 66866 164400 6 la_output[19]
port 492 nsew signal output
rlabel metal2 s 6274 163200 6330 164400 6 la_output[1]
port 493 nsew signal output
rlabel metal2 s 70122 163200 70178 164400 6 la_output[20]
port 494 nsew signal output
rlabel metal2 s 73526 163200 73582 164400 6 la_output[21]
port 495 nsew signal output
rlabel metal2 s 76930 163200 76986 164400 6 la_output[22]
port 496 nsew signal output
rlabel metal2 s 80242 163200 80298 164400 6 la_output[23]
port 497 nsew signal output
rlabel metal2 s 83646 163200 83702 164400 6 la_output[24]
port 498 nsew signal output
rlabel metal2 s 86958 163200 87014 164400 6 la_output[25]
port 499 nsew signal output
rlabel metal2 s 90362 163200 90418 164400 6 la_output[26]
port 500 nsew signal output
rlabel metal2 s 93674 163200 93730 164400 6 la_output[27]
port 501 nsew signal output
rlabel metal2 s 97078 163200 97134 164400 6 la_output[28]
port 502 nsew signal output
rlabel metal2 s 100482 163200 100538 164400 6 la_output[29]
port 503 nsew signal output
rlabel metal2 s 9586 163200 9642 164400 6 la_output[2]
port 504 nsew signal output
rlabel metal2 s 103794 163200 103850 164400 6 la_output[30]
port 505 nsew signal output
rlabel metal2 s 107198 163200 107254 164400 6 la_output[31]
port 506 nsew signal output
rlabel metal2 s 110510 163200 110566 164400 6 la_output[32]
port 507 nsew signal output
rlabel metal2 s 113914 163200 113970 164400 6 la_output[33]
port 508 nsew signal output
rlabel metal2 s 117226 163200 117282 164400 6 la_output[34]
port 509 nsew signal output
rlabel metal2 s 120630 163200 120686 164400 6 la_output[35]
port 510 nsew signal output
rlabel metal2 s 124034 163200 124090 164400 6 la_output[36]
port 511 nsew signal output
rlabel metal2 s 127346 163200 127402 164400 6 la_output[37]
port 512 nsew signal output
rlabel metal2 s 130750 163200 130806 164400 6 la_output[38]
port 513 nsew signal output
rlabel metal2 s 134062 163200 134118 164400 6 la_output[39]
port 514 nsew signal output
rlabel metal2 s 12990 163200 13046 164400 6 la_output[3]
port 515 nsew signal output
rlabel metal2 s 137466 163200 137522 164400 6 la_output[40]
port 516 nsew signal output
rlabel metal2 s 140778 163200 140834 164400 6 la_output[41]
port 517 nsew signal output
rlabel metal2 s 144182 163200 144238 164400 6 la_output[42]
port 518 nsew signal output
rlabel metal2 s 147586 163200 147642 164400 6 la_output[43]
port 519 nsew signal output
rlabel metal2 s 150898 163200 150954 164400 6 la_output[44]
port 520 nsew signal output
rlabel metal2 s 154302 163200 154358 164400 6 la_output[45]
port 521 nsew signal output
rlabel metal2 s 157614 163200 157670 164400 6 la_output[46]
port 522 nsew signal output
rlabel metal2 s 161018 163200 161074 164400 6 la_output[47]
port 523 nsew signal output
rlabel metal2 s 164330 163200 164386 164400 6 la_output[48]
port 524 nsew signal output
rlabel metal2 s 167734 163200 167790 164400 6 la_output[49]
port 525 nsew signal output
rlabel metal2 s 16302 163200 16358 164400 6 la_output[4]
port 526 nsew signal output
rlabel metal2 s 171138 163200 171194 164400 6 la_output[50]
port 527 nsew signal output
rlabel metal2 s 174450 163200 174506 164400 6 la_output[51]
port 528 nsew signal output
rlabel metal2 s 177854 163200 177910 164400 6 la_output[52]
port 529 nsew signal output
rlabel metal2 s 181166 163200 181222 164400 6 la_output[53]
port 530 nsew signal output
rlabel metal2 s 184570 163200 184626 164400 6 la_output[54]
port 531 nsew signal output
rlabel metal2 s 187882 163200 187938 164400 6 la_output[55]
port 532 nsew signal output
rlabel metal2 s 191286 163200 191342 164400 6 la_output[56]
port 533 nsew signal output
rlabel metal2 s 194690 163200 194746 164400 6 la_output[57]
port 534 nsew signal output
rlabel metal2 s 198002 163200 198058 164400 6 la_output[58]
port 535 nsew signal output
rlabel metal2 s 201406 163200 201462 164400 6 la_output[59]
port 536 nsew signal output
rlabel metal2 s 19706 163200 19762 164400 6 la_output[5]
port 537 nsew signal output
rlabel metal2 s 204718 163200 204774 164400 6 la_output[60]
port 538 nsew signal output
rlabel metal2 s 208122 163200 208178 164400 6 la_output[61]
port 539 nsew signal output
rlabel metal2 s 211434 163200 211490 164400 6 la_output[62]
port 540 nsew signal output
rlabel metal2 s 214838 163200 214894 164400 6 la_output[63]
port 541 nsew signal output
rlabel metal2 s 218242 163200 218298 164400 6 la_output[64]
port 542 nsew signal output
rlabel metal2 s 221554 163200 221610 164400 6 la_output[65]
port 543 nsew signal output
rlabel metal2 s 224958 163200 225014 164400 6 la_output[66]
port 544 nsew signal output
rlabel metal2 s 228270 163200 228326 164400 6 la_output[67]
port 545 nsew signal output
rlabel metal2 s 231674 163200 231730 164400 6 la_output[68]
port 546 nsew signal output
rlabel metal2 s 234986 163200 235042 164400 6 la_output[69]
port 547 nsew signal output
rlabel metal2 s 23018 163200 23074 164400 6 la_output[6]
port 548 nsew signal output
rlabel metal2 s 238390 163200 238446 164400 6 la_output[70]
port 549 nsew signal output
rlabel metal2 s 241794 163200 241850 164400 6 la_output[71]
port 550 nsew signal output
rlabel metal2 s 245106 163200 245162 164400 6 la_output[72]
port 551 nsew signal output
rlabel metal2 s 248510 163200 248566 164400 6 la_output[73]
port 552 nsew signal output
rlabel metal2 s 251822 163200 251878 164400 6 la_output[74]
port 553 nsew signal output
rlabel metal2 s 255226 163200 255282 164400 6 la_output[75]
port 554 nsew signal output
rlabel metal2 s 258538 163200 258594 164400 6 la_output[76]
port 555 nsew signal output
rlabel metal2 s 261942 163200 261998 164400 6 la_output[77]
port 556 nsew signal output
rlabel metal2 s 265346 163200 265402 164400 6 la_output[78]
port 557 nsew signal output
rlabel metal2 s 268658 163200 268714 164400 6 la_output[79]
port 558 nsew signal output
rlabel metal2 s 26422 163200 26478 164400 6 la_output[7]
port 559 nsew signal output
rlabel metal2 s 272062 163200 272118 164400 6 la_output[80]
port 560 nsew signal output
rlabel metal2 s 275374 163200 275430 164400 6 la_output[81]
port 561 nsew signal output
rlabel metal2 s 278778 163200 278834 164400 6 la_output[82]
port 562 nsew signal output
rlabel metal2 s 282090 163200 282146 164400 6 la_output[83]
port 563 nsew signal output
rlabel metal2 s 285494 163200 285550 164400 6 la_output[84]
port 564 nsew signal output
rlabel metal2 s 288898 163200 288954 164400 6 la_output[85]
port 565 nsew signal output
rlabel metal2 s 292210 163200 292266 164400 6 la_output[86]
port 566 nsew signal output
rlabel metal2 s 295614 163200 295670 164400 6 la_output[87]
port 567 nsew signal output
rlabel metal2 s 298926 163200 298982 164400 6 la_output[88]
port 568 nsew signal output
rlabel metal2 s 302330 163200 302386 164400 6 la_output[89]
port 569 nsew signal output
rlabel metal2 s 29826 163200 29882 164400 6 la_output[8]
port 570 nsew signal output
rlabel metal2 s 305642 163200 305698 164400 6 la_output[90]
port 571 nsew signal output
rlabel metal2 s 309046 163200 309102 164400 6 la_output[91]
port 572 nsew signal output
rlabel metal2 s 312450 163200 312506 164400 6 la_output[92]
port 573 nsew signal output
rlabel metal2 s 315762 163200 315818 164400 6 la_output[93]
port 574 nsew signal output
rlabel metal2 s 319166 163200 319222 164400 6 la_output[94]
port 575 nsew signal output
rlabel metal2 s 322478 163200 322534 164400 6 la_output[95]
port 576 nsew signal output
rlabel metal2 s 325882 163200 325938 164400 6 la_output[96]
port 577 nsew signal output
rlabel metal2 s 329194 163200 329250 164400 6 la_output[97]
port 578 nsew signal output
rlabel metal2 s 332598 163200 332654 164400 6 la_output[98]
port 579 nsew signal output
rlabel metal2 s 336002 163200 336058 164400 6 la_output[99]
port 580 nsew signal output
rlabel metal2 s 33138 163200 33194 164400 6 la_output[9]
port 581 nsew signal output
rlabel metal2 s 431038 163200 431094 164400 6 mprj_ack_i
port 582 nsew signal input
rlabel metal2 s 435178 163200 435234 164400 6 mprj_adr_o[0]
port 583 nsew signal output
rlabel metal2 s 463790 163200 463846 164400 6 mprj_adr_o[10]
port 584 nsew signal output
rlabel metal2 s 466366 163200 466422 164400 6 mprj_adr_o[11]
port 585 nsew signal output
rlabel metal2 s 468850 163200 468906 164400 6 mprj_adr_o[12]
port 586 nsew signal output
rlabel metal2 s 471426 163200 471482 164400 6 mprj_adr_o[13]
port 587 nsew signal output
rlabel metal2 s 473910 163200 473966 164400 6 mprj_adr_o[14]
port 588 nsew signal output
rlabel metal2 s 476394 163200 476450 164400 6 mprj_adr_o[15]
port 589 nsew signal output
rlabel metal2 s 478970 163200 479026 164400 6 mprj_adr_o[16]
port 590 nsew signal output
rlabel metal2 s 481454 163200 481510 164400 6 mprj_adr_o[17]
port 591 nsew signal output
rlabel metal2 s 484030 163200 484086 164400 6 mprj_adr_o[18]
port 592 nsew signal output
rlabel metal2 s 486514 163200 486570 164400 6 mprj_adr_o[19]
port 593 nsew signal output
rlabel metal2 s 438582 163200 438638 164400 6 mprj_adr_o[1]
port 594 nsew signal output
rlabel metal2 s 489090 163200 489146 164400 6 mprj_adr_o[20]
port 595 nsew signal output
rlabel metal2 s 491574 163200 491630 164400 6 mprj_adr_o[21]
port 596 nsew signal output
rlabel metal2 s 494058 163200 494114 164400 6 mprj_adr_o[22]
port 597 nsew signal output
rlabel metal2 s 496634 163200 496690 164400 6 mprj_adr_o[23]
port 598 nsew signal output
rlabel metal2 s 499118 163200 499174 164400 6 mprj_adr_o[24]
port 599 nsew signal output
rlabel metal2 s 501694 163200 501750 164400 6 mprj_adr_o[25]
port 600 nsew signal output
rlabel metal2 s 504178 163200 504234 164400 6 mprj_adr_o[26]
port 601 nsew signal output
rlabel metal2 s 506754 163200 506810 164400 6 mprj_adr_o[27]
port 602 nsew signal output
rlabel metal2 s 509238 163200 509294 164400 6 mprj_adr_o[28]
port 603 nsew signal output
rlabel metal2 s 511722 163200 511778 164400 6 mprj_adr_o[29]
port 604 nsew signal output
rlabel metal2 s 441986 163200 442042 164400 6 mprj_adr_o[2]
port 605 nsew signal output
rlabel metal2 s 514298 163200 514354 164400 6 mprj_adr_o[30]
port 606 nsew signal output
rlabel metal2 s 516782 163200 516838 164400 6 mprj_adr_o[31]
port 607 nsew signal output
rlabel metal2 s 445298 163200 445354 164400 6 mprj_adr_o[3]
port 608 nsew signal output
rlabel metal2 s 448702 163200 448758 164400 6 mprj_adr_o[4]
port 609 nsew signal output
rlabel metal2 s 451186 163200 451242 164400 6 mprj_adr_o[5]
port 610 nsew signal output
rlabel metal2 s 453762 163200 453818 164400 6 mprj_adr_o[6]
port 611 nsew signal output
rlabel metal2 s 456246 163200 456302 164400 6 mprj_adr_o[7]
port 612 nsew signal output
rlabel metal2 s 458730 163200 458786 164400 6 mprj_adr_o[8]
port 613 nsew signal output
rlabel metal2 s 461306 163200 461362 164400 6 mprj_adr_o[9]
port 614 nsew signal output
rlabel metal2 s 431866 163200 431922 164400 6 mprj_cyc_o
port 615 nsew signal output
rlabel metal2 s 436098 163200 436154 164400 6 mprj_dat_i[0]
port 616 nsew signal input
rlabel metal2 s 464618 163200 464674 164400 6 mprj_dat_i[10]
port 617 nsew signal input
rlabel metal2 s 467194 163200 467250 164400 6 mprj_dat_i[11]
port 618 nsew signal input
rlabel metal2 s 469678 163200 469734 164400 6 mprj_dat_i[12]
port 619 nsew signal input
rlabel metal2 s 472254 163200 472310 164400 6 mprj_dat_i[13]
port 620 nsew signal input
rlabel metal2 s 474738 163200 474794 164400 6 mprj_dat_i[14]
port 621 nsew signal input
rlabel metal2 s 477314 163200 477370 164400 6 mprj_dat_i[15]
port 622 nsew signal input
rlabel metal2 s 479798 163200 479854 164400 6 mprj_dat_i[16]
port 623 nsew signal input
rlabel metal2 s 482282 163200 482338 164400 6 mprj_dat_i[17]
port 624 nsew signal input
rlabel metal2 s 484858 163200 484914 164400 6 mprj_dat_i[18]
port 625 nsew signal input
rlabel metal2 s 487342 163200 487398 164400 6 mprj_dat_i[19]
port 626 nsew signal input
rlabel metal2 s 439410 163200 439466 164400 6 mprj_dat_i[1]
port 627 nsew signal input
rlabel metal2 s 489918 163200 489974 164400 6 mprj_dat_i[20]
port 628 nsew signal input
rlabel metal2 s 492402 163200 492458 164400 6 mprj_dat_i[21]
port 629 nsew signal input
rlabel metal2 s 494978 163200 495034 164400 6 mprj_dat_i[22]
port 630 nsew signal input
rlabel metal2 s 497462 163200 497518 164400 6 mprj_dat_i[23]
port 631 nsew signal input
rlabel metal2 s 499946 163200 500002 164400 6 mprj_dat_i[24]
port 632 nsew signal input
rlabel metal2 s 502522 163200 502578 164400 6 mprj_dat_i[25]
port 633 nsew signal input
rlabel metal2 s 505006 163200 505062 164400 6 mprj_dat_i[26]
port 634 nsew signal input
rlabel metal2 s 507582 163200 507638 164400 6 mprj_dat_i[27]
port 635 nsew signal input
rlabel metal2 s 510066 163200 510122 164400 6 mprj_dat_i[28]
port 636 nsew signal input
rlabel metal2 s 512642 163200 512698 164400 6 mprj_dat_i[29]
port 637 nsew signal input
rlabel metal2 s 442814 163200 442870 164400 6 mprj_dat_i[2]
port 638 nsew signal input
rlabel metal2 s 515126 163200 515182 164400 6 mprj_dat_i[30]
port 639 nsew signal input
rlabel metal2 s 517610 163200 517666 164400 6 mprj_dat_i[31]
port 640 nsew signal input
rlabel metal2 s 446126 163200 446182 164400 6 mprj_dat_i[3]
port 641 nsew signal input
rlabel metal2 s 449530 163200 449586 164400 6 mprj_dat_i[4]
port 642 nsew signal input
rlabel metal2 s 452014 163200 452070 164400 6 mprj_dat_i[5]
port 643 nsew signal input
rlabel metal2 s 454590 163200 454646 164400 6 mprj_dat_i[6]
port 644 nsew signal input
rlabel metal2 s 457074 163200 457130 164400 6 mprj_dat_i[7]
port 645 nsew signal input
rlabel metal2 s 459650 163200 459706 164400 6 mprj_dat_i[8]
port 646 nsew signal input
rlabel metal2 s 462134 163200 462190 164400 6 mprj_dat_i[9]
port 647 nsew signal input
rlabel metal2 s 436926 163200 436982 164400 6 mprj_dat_o[0]
port 648 nsew signal output
rlabel metal2 s 465538 163200 465594 164400 6 mprj_dat_o[10]
port 649 nsew signal output
rlabel metal2 s 468022 163200 468078 164400 6 mprj_dat_o[11]
port 650 nsew signal output
rlabel metal2 s 470506 163200 470562 164400 6 mprj_dat_o[12]
port 651 nsew signal output
rlabel metal2 s 473082 163200 473138 164400 6 mprj_dat_o[13]
port 652 nsew signal output
rlabel metal2 s 475566 163200 475622 164400 6 mprj_dat_o[14]
port 653 nsew signal output
rlabel metal2 s 478142 163200 478198 164400 6 mprj_dat_o[15]
port 654 nsew signal output
rlabel metal2 s 480626 163200 480682 164400 6 mprj_dat_o[16]
port 655 nsew signal output
rlabel metal2 s 483202 163200 483258 164400 6 mprj_dat_o[17]
port 656 nsew signal output
rlabel metal2 s 485686 163200 485742 164400 6 mprj_dat_o[18]
port 657 nsew signal output
rlabel metal2 s 488170 163200 488226 164400 6 mprj_dat_o[19]
port 658 nsew signal output
rlabel metal2 s 440238 163200 440294 164400 6 mprj_dat_o[1]
port 659 nsew signal output
rlabel metal2 s 490746 163200 490802 164400 6 mprj_dat_o[20]
port 660 nsew signal output
rlabel metal2 s 493230 163200 493286 164400 6 mprj_dat_o[21]
port 661 nsew signal output
rlabel metal2 s 495806 163200 495862 164400 6 mprj_dat_o[22]
port 662 nsew signal output
rlabel metal2 s 498290 163200 498346 164400 6 mprj_dat_o[23]
port 663 nsew signal output
rlabel metal2 s 500866 163200 500922 164400 6 mprj_dat_o[24]
port 664 nsew signal output
rlabel metal2 s 503350 163200 503406 164400 6 mprj_dat_o[25]
port 665 nsew signal output
rlabel metal2 s 505834 163200 505890 164400 6 mprj_dat_o[26]
port 666 nsew signal output
rlabel metal2 s 508410 163200 508466 164400 6 mprj_dat_o[27]
port 667 nsew signal output
rlabel metal2 s 510894 163200 510950 164400 6 mprj_dat_o[28]
port 668 nsew signal output
rlabel metal2 s 513470 163200 513526 164400 6 mprj_dat_o[29]
port 669 nsew signal output
rlabel metal2 s 443642 163200 443698 164400 6 mprj_dat_o[2]
port 670 nsew signal output
rlabel metal2 s 515954 163200 516010 164400 6 mprj_dat_o[30]
port 671 nsew signal output
rlabel metal2 s 518530 163200 518586 164400 6 mprj_dat_o[31]
port 672 nsew signal output
rlabel metal2 s 446954 163200 447010 164400 6 mprj_dat_o[3]
port 673 nsew signal output
rlabel metal2 s 450358 163200 450414 164400 6 mprj_dat_o[4]
port 674 nsew signal output
rlabel metal2 s 452842 163200 452898 164400 6 mprj_dat_o[5]
port 675 nsew signal output
rlabel metal2 s 455418 163200 455474 164400 6 mprj_dat_o[6]
port 676 nsew signal output
rlabel metal2 s 457902 163200 457958 164400 6 mprj_dat_o[7]
port 677 nsew signal output
rlabel metal2 s 460478 163200 460534 164400 6 mprj_dat_o[8]
port 678 nsew signal output
rlabel metal2 s 462962 163200 463018 164400 6 mprj_dat_o[9]
port 679 nsew signal output
rlabel metal2 s 437754 163200 437810 164400 6 mprj_sel_o[0]
port 680 nsew signal output
rlabel metal2 s 441066 163200 441122 164400 6 mprj_sel_o[1]
port 681 nsew signal output
rlabel metal2 s 444470 163200 444526 164400 6 mprj_sel_o[2]
port 682 nsew signal output
rlabel metal2 s 447874 163200 447930 164400 6 mprj_sel_o[3]
port 683 nsew signal output
rlabel metal2 s 432694 163200 432750 164400 6 mprj_stb_o
port 684 nsew signal output
rlabel metal2 s 433522 163200 433578 164400 6 mprj_wb_iena
port 685 nsew signal output
rlabel metal2 s 434350 163200 434406 164400 6 mprj_we_o
port 686 nsew signal output
rlabel metal3 s 523200 89360 524400 89480 6 qspi_enabled
port 687 nsew signal output
rlabel metal3 s 523200 83376 524400 83496 6 ser_rx
port 688 nsew signal input
rlabel metal3 s 523200 84872 524400 84992 6 ser_tx
port 689 nsew signal output
rlabel metal3 s 523200 80384 524400 80504 6 spi_csb
port 690 nsew signal output
rlabel metal3 s 523200 86368 524400 86488 6 spi_enabled
port 691 nsew signal output
rlabel metal3 s 523200 78888 524400 79008 6 spi_sck
port 692 nsew signal output
rlabel metal3 s 523200 81880 524400 82000 6 spi_sdi
port 693 nsew signal input
rlabel metal3 s 523200 77392 524400 77512 6 spi_sdo
port 694 nsew signal output
rlabel metal3 s 523200 75896 524400 76016 6 spi_sdoenb
port 695 nsew signal output
rlabel metal3 s 523200 2184 524400 2304 6 sram_ro_addr[0]
port 696 nsew signal input
rlabel metal3 s 523200 3680 524400 3800 6 sram_ro_addr[1]
port 697 nsew signal input
rlabel metal3 s 523200 5176 524400 5296 6 sram_ro_addr[2]
port 698 nsew signal input
rlabel metal3 s 523200 6672 524400 6792 6 sram_ro_addr[3]
port 699 nsew signal input
rlabel metal3 s 523200 8168 524400 8288 6 sram_ro_addr[4]
port 700 nsew signal input
rlabel metal3 s 523200 9664 524400 9784 6 sram_ro_addr[5]
port 701 nsew signal input
rlabel metal3 s 523200 11160 524400 11280 6 sram_ro_addr[6]
port 702 nsew signal input
rlabel metal3 s 523200 12656 524400 12776 6 sram_ro_addr[7]
port 703 nsew signal input
rlabel metal3 s 523200 14152 524400 14272 6 sram_ro_clk
port 704 nsew signal input
rlabel metal3 s 523200 688 524400 808 6 sram_ro_csb
port 705 nsew signal input
rlabel metal3 s 523200 15648 524400 15768 6 sram_ro_data[0]
port 706 nsew signal output
rlabel metal3 s 523200 30744 524400 30864 6 sram_ro_data[10]
port 707 nsew signal output
rlabel metal3 s 523200 32240 524400 32360 6 sram_ro_data[11]
port 708 nsew signal output
rlabel metal3 s 523200 33736 524400 33856 6 sram_ro_data[12]
port 709 nsew signal output
rlabel metal3 s 523200 35232 524400 35352 6 sram_ro_data[13]
port 710 nsew signal output
rlabel metal3 s 523200 36728 524400 36848 6 sram_ro_data[14]
port 711 nsew signal output
rlabel metal3 s 523200 38224 524400 38344 6 sram_ro_data[15]
port 712 nsew signal output
rlabel metal3 s 523200 39720 524400 39840 6 sram_ro_data[16]
port 713 nsew signal output
rlabel metal3 s 523200 41216 524400 41336 6 sram_ro_data[17]
port 714 nsew signal output
rlabel metal3 s 523200 42712 524400 42832 6 sram_ro_data[18]
port 715 nsew signal output
rlabel metal3 s 523200 44208 524400 44328 6 sram_ro_data[19]
port 716 nsew signal output
rlabel metal3 s 523200 17144 524400 17264 6 sram_ro_data[1]
port 717 nsew signal output
rlabel metal3 s 523200 45704 524400 45824 6 sram_ro_data[20]
port 718 nsew signal output
rlabel metal3 s 523200 47200 524400 47320 6 sram_ro_data[21]
port 719 nsew signal output
rlabel metal3 s 523200 48832 524400 48952 6 sram_ro_data[22]
port 720 nsew signal output
rlabel metal3 s 523200 50328 524400 50448 6 sram_ro_data[23]
port 721 nsew signal output
rlabel metal3 s 523200 51824 524400 51944 6 sram_ro_data[24]
port 722 nsew signal output
rlabel metal3 s 523200 53320 524400 53440 6 sram_ro_data[25]
port 723 nsew signal output
rlabel metal3 s 523200 54816 524400 54936 6 sram_ro_data[26]
port 724 nsew signal output
rlabel metal3 s 523200 56312 524400 56432 6 sram_ro_data[27]
port 725 nsew signal output
rlabel metal3 s 523200 57808 524400 57928 6 sram_ro_data[28]
port 726 nsew signal output
rlabel metal3 s 523200 59304 524400 59424 6 sram_ro_data[29]
port 727 nsew signal output
rlabel metal3 s 523200 18640 524400 18760 6 sram_ro_data[2]
port 728 nsew signal output
rlabel metal3 s 523200 60800 524400 60920 6 sram_ro_data[30]
port 729 nsew signal output
rlabel metal3 s 523200 62296 524400 62416 6 sram_ro_data[31]
port 730 nsew signal output
rlabel metal3 s 523200 20136 524400 20256 6 sram_ro_data[3]
port 731 nsew signal output
rlabel metal3 s 523200 21632 524400 21752 6 sram_ro_data[4]
port 732 nsew signal output
rlabel metal3 s 523200 23128 524400 23248 6 sram_ro_data[5]
port 733 nsew signal output
rlabel metal3 s 523200 24760 524400 24880 6 sram_ro_data[6]
port 734 nsew signal output
rlabel metal3 s 523200 26256 524400 26376 6 sram_ro_data[7]
port 735 nsew signal output
rlabel metal3 s 523200 27752 524400 27872 6 sram_ro_data[8]
port 736 nsew signal output
rlabel metal3 s 523200 29248 524400 29368 6 sram_ro_data[9]
port 737 nsew signal output
rlabel metal3 s 523200 69776 524400 69896 6 trap
port 738 nsew signal output
rlabel metal3 s 523200 87864 524400 87984 6 uart_enabled
port 739 nsew signal output
rlabel metal2 s 519358 163200 519414 164400 6 user_irq_ena[0]
port 740 nsew signal output
rlabel metal2 s 520186 163200 520242 164400 6 user_irq_ena[1]
port 741 nsew signal output
rlabel metal2 s 521014 163200 521070 164400 6 user_irq_ena[2]
port 742 nsew signal output
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 524000 164000
string LEFview TRUE
string GDS_FILE ../gds/mgmt_core_wrapper.gds
string GDS_END 183921168
string GDS_START 182803602
<< end >>

