// This is the unpowered netlist.
module RAM128 (CLK,
    EN0,
    A0,
    Di0,
    Do0,
    WE0);
 input CLK;
 input EN0;
 input [6:0] A0;
 input [31:0] Di0;
 output [31:0] Do0;
 input [3:0] WE0;

 wire \A0BUF[0].X ;
 wire \A0BUF[1].X ;
 wire \A0BUF[2].X ;
 wire \A0BUF[3].X ;
 wire \A0BUF[4].X ;
 wire \A0BUF[5].X ;
 wire \A0BUF[6].X ;
 wire \BLOCK[0].RAM32.A0BUF[0].X ;
 wire \BLOCK[0].RAM32.A0BUF[1].X ;
 wire \BLOCK[0].RAM32.A0BUF[2].X ;
 wire \BLOCK[0].RAM32.A0BUF[3].X ;
 wire \BLOCK[0].RAM32.A0BUF[4].X ;
 wire \BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].A ;
 wire \BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ;
 wire \BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ;
 wire \BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ;
 wire \BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ;
 wire \BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ;
 wire \BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ;
 wire \BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ;
 wire \BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ;
 wire \BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].A ;
 wire \BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].TE_B ;
 wire \BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ;
 wire \BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ;
 wire \BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ;
 wire \BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ;
 wire \BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ;
 wire \BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ;
 wire \BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ;
 wire \BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ;
 wire \BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].A ;
 wire \BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].TE_B ;
 wire \BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ;
 wire \BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ;
 wire \BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ;
 wire \BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ;
 wire \BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ;
 wire \BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ;
 wire \BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ;
 wire \BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ;
 wire \BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].A ;
 wire \BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].TE_B ;
 wire \BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ;
 wire \BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ;
 wire \BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ;
 wire \BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ;
 wire \BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ;
 wire \BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ;
 wire \BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ;
 wire \BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ;
 wire \BLOCK[0].RAM32.CLK ;
 wire \BLOCK[0].RAM32.CLKBUF.X ;
 wire \BLOCK[0].RAM32.DEC0.EN ;
 wire \BLOCK[0].RAM32.DIBUF[0].A ;
 wire \BLOCK[0].RAM32.DIBUF[0].X ;
 wire \BLOCK[0].RAM32.DIBUF[10].A ;
 wire \BLOCK[0].RAM32.DIBUF[10].X ;
 wire \BLOCK[0].RAM32.DIBUF[11].A ;
 wire \BLOCK[0].RAM32.DIBUF[11].X ;
 wire \BLOCK[0].RAM32.DIBUF[12].A ;
 wire \BLOCK[0].RAM32.DIBUF[12].X ;
 wire \BLOCK[0].RAM32.DIBUF[13].A ;
 wire \BLOCK[0].RAM32.DIBUF[13].X ;
 wire \BLOCK[0].RAM32.DIBUF[14].A ;
 wire \BLOCK[0].RAM32.DIBUF[14].X ;
 wire \BLOCK[0].RAM32.DIBUF[15].A ;
 wire \BLOCK[0].RAM32.DIBUF[15].X ;
 wire \BLOCK[0].RAM32.DIBUF[16].A ;
 wire \BLOCK[0].RAM32.DIBUF[16].X ;
 wire \BLOCK[0].RAM32.DIBUF[17].A ;
 wire \BLOCK[0].RAM32.DIBUF[17].X ;
 wire \BLOCK[0].RAM32.DIBUF[18].A ;
 wire \BLOCK[0].RAM32.DIBUF[18].X ;
 wire \BLOCK[0].RAM32.DIBUF[19].A ;
 wire \BLOCK[0].RAM32.DIBUF[19].X ;
 wire \BLOCK[0].RAM32.DIBUF[1].A ;
 wire \BLOCK[0].RAM32.DIBUF[1].X ;
 wire \BLOCK[0].RAM32.DIBUF[20].A ;
 wire \BLOCK[0].RAM32.DIBUF[20].X ;
 wire \BLOCK[0].RAM32.DIBUF[21].A ;
 wire \BLOCK[0].RAM32.DIBUF[21].X ;
 wire \BLOCK[0].RAM32.DIBUF[22].A ;
 wire \BLOCK[0].RAM32.DIBUF[22].X ;
 wire \BLOCK[0].RAM32.DIBUF[23].A ;
 wire \BLOCK[0].RAM32.DIBUF[23].X ;
 wire \BLOCK[0].RAM32.DIBUF[24].A ;
 wire \BLOCK[0].RAM32.DIBUF[24].X ;
 wire \BLOCK[0].RAM32.DIBUF[25].A ;
 wire \BLOCK[0].RAM32.DIBUF[25].X ;
 wire \BLOCK[0].RAM32.DIBUF[26].A ;
 wire \BLOCK[0].RAM32.DIBUF[26].X ;
 wire \BLOCK[0].RAM32.DIBUF[27].A ;
 wire \BLOCK[0].RAM32.DIBUF[27].X ;
 wire \BLOCK[0].RAM32.DIBUF[28].A ;
 wire \BLOCK[0].RAM32.DIBUF[28].X ;
 wire \BLOCK[0].RAM32.DIBUF[29].A ;
 wire \BLOCK[0].RAM32.DIBUF[29].X ;
 wire \BLOCK[0].RAM32.DIBUF[2].A ;
 wire \BLOCK[0].RAM32.DIBUF[2].X ;
 wire \BLOCK[0].RAM32.DIBUF[30].A ;
 wire \BLOCK[0].RAM32.DIBUF[30].X ;
 wire \BLOCK[0].RAM32.DIBUF[31].A ;
 wire \BLOCK[0].RAM32.DIBUF[31].X ;
 wire \BLOCK[0].RAM32.DIBUF[3].A ;
 wire \BLOCK[0].RAM32.DIBUF[3].X ;
 wire \BLOCK[0].RAM32.DIBUF[4].A ;
 wire \BLOCK[0].RAM32.DIBUF[4].X ;
 wire \BLOCK[0].RAM32.DIBUF[5].A ;
 wire \BLOCK[0].RAM32.DIBUF[5].X ;
 wire \BLOCK[0].RAM32.DIBUF[6].A ;
 wire \BLOCK[0].RAM32.DIBUF[6].X ;
 wire \BLOCK[0].RAM32.DIBUF[7].A ;
 wire \BLOCK[0].RAM32.DIBUF[7].X ;
 wire \BLOCK[0].RAM32.DIBUF[8].A ;
 wire \BLOCK[0].RAM32.DIBUF[8].X ;
 wire \BLOCK[0].RAM32.DIBUF[9].A ;
 wire \BLOCK[0].RAM32.DIBUF[9].X ;
 wire \BLOCK[0].RAM32.Do0[0] ;
 wire \BLOCK[0].RAM32.Do0[10] ;
 wire \BLOCK[0].RAM32.Do0[11] ;
 wire \BLOCK[0].RAM32.Do0[12] ;
 wire \BLOCK[0].RAM32.Do0[13] ;
 wire \BLOCK[0].RAM32.Do0[14] ;
 wire \BLOCK[0].RAM32.Do0[15] ;
 wire \BLOCK[0].RAM32.Do0[16] ;
 wire \BLOCK[0].RAM32.Do0[17] ;
 wire \BLOCK[0].RAM32.Do0[18] ;
 wire \BLOCK[0].RAM32.Do0[19] ;
 wire \BLOCK[0].RAM32.Do0[1] ;
 wire \BLOCK[0].RAM32.Do0[20] ;
 wire \BLOCK[0].RAM32.Do0[21] ;
 wire \BLOCK[0].RAM32.Do0[22] ;
 wire \BLOCK[0].RAM32.Do0[23] ;
 wire \BLOCK[0].RAM32.Do0[24] ;
 wire \BLOCK[0].RAM32.Do0[25] ;
 wire \BLOCK[0].RAM32.Do0[26] ;
 wire \BLOCK[0].RAM32.Do0[27] ;
 wire \BLOCK[0].RAM32.Do0[28] ;
 wire \BLOCK[0].RAM32.Do0[29] ;
 wire \BLOCK[0].RAM32.Do0[2] ;
 wire \BLOCK[0].RAM32.Do0[30] ;
 wire \BLOCK[0].RAM32.Do0[31] ;
 wire \BLOCK[0].RAM32.Do0[3] ;
 wire \BLOCK[0].RAM32.Do0[4] ;
 wire \BLOCK[0].RAM32.Do0[5] ;
 wire \BLOCK[0].RAM32.Do0[6] ;
 wire \BLOCK[0].RAM32.Do0[7] ;
 wire \BLOCK[0].RAM32.Do0[8] ;
 wire \BLOCK[0].RAM32.Do0[9] ;
 wire \BLOCK[0].RAM32.Do0_REG.CLKBUF[0] ;
 wire \BLOCK[0].RAM32.Do0_REG.CLKBUF[1] ;
 wire \BLOCK[0].RAM32.Do0_REG.CLKBUF[2] ;
 wire \BLOCK[0].RAM32.Do0_REG.CLKBUF[3] ;
 wire \BLOCK[0].RAM32.Do0_REG.CLK_buf ;
 wire \BLOCK[0].RAM32.EN0 ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.CLKBUF.X ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.EN ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[0].A ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[0].X ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[1].A ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[1].X ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[2].A ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[2].X ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[3].A ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[3].X ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.CLKBUF.X ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.EN ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[0].X ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[1].X ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[2].X ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[3].X ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.CLKBUF.X ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.EN ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.EN_buf ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[0].X ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[1].X ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[2].X ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[3].X ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.CLKBUF.X ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.EN ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.EN_buf ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[0].X ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[1].X ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[2].X ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[3].X ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.SEL0 ;
 wire \BLOCK[0].RAM32.WEBUF[0].A ;
 wire \BLOCK[0].RAM32.WEBUF[1].A ;
 wire \BLOCK[0].RAM32.WEBUF[2].A ;
 wire \BLOCK[0].RAM32.WEBUF[3].A ;
 wire \BLOCK[1].RAM32.A0BUF[0].X ;
 wire \BLOCK[1].RAM32.A0BUF[1].X ;
 wire \BLOCK[1].RAM32.A0BUF[2].X ;
 wire \BLOCK[1].RAM32.A0BUF[3].X ;
 wire \BLOCK[1].RAM32.A0BUF[4].X ;
 wire \BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].A ;
 wire \BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ;
 wire \BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ;
 wire \BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ;
 wire \BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ;
 wire \BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ;
 wire \BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ;
 wire \BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ;
 wire \BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ;
 wire \BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].A ;
 wire \BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].TE_B ;
 wire \BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ;
 wire \BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ;
 wire \BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ;
 wire \BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ;
 wire \BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ;
 wire \BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ;
 wire \BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ;
 wire \BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ;
 wire \BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].A ;
 wire \BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].TE_B ;
 wire \BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ;
 wire \BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ;
 wire \BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ;
 wire \BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ;
 wire \BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ;
 wire \BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ;
 wire \BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ;
 wire \BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ;
 wire \BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].A ;
 wire \BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].TE_B ;
 wire \BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ;
 wire \BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ;
 wire \BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ;
 wire \BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ;
 wire \BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ;
 wire \BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ;
 wire \BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ;
 wire \BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ;
 wire \BLOCK[1].RAM32.CLKBUF.X ;
 wire \BLOCK[1].RAM32.DEC0.EN ;
 wire \BLOCK[1].RAM32.DIBUF[0].X ;
 wire \BLOCK[1].RAM32.DIBUF[10].X ;
 wire \BLOCK[1].RAM32.DIBUF[11].X ;
 wire \BLOCK[1].RAM32.DIBUF[12].X ;
 wire \BLOCK[1].RAM32.DIBUF[13].X ;
 wire \BLOCK[1].RAM32.DIBUF[14].X ;
 wire \BLOCK[1].RAM32.DIBUF[15].X ;
 wire \BLOCK[1].RAM32.DIBUF[16].X ;
 wire \BLOCK[1].RAM32.DIBUF[17].X ;
 wire \BLOCK[1].RAM32.DIBUF[18].X ;
 wire \BLOCK[1].RAM32.DIBUF[19].X ;
 wire \BLOCK[1].RAM32.DIBUF[1].X ;
 wire \BLOCK[1].RAM32.DIBUF[20].X ;
 wire \BLOCK[1].RAM32.DIBUF[21].X ;
 wire \BLOCK[1].RAM32.DIBUF[22].X ;
 wire \BLOCK[1].RAM32.DIBUF[23].X ;
 wire \BLOCK[1].RAM32.DIBUF[24].X ;
 wire \BLOCK[1].RAM32.DIBUF[25].X ;
 wire \BLOCK[1].RAM32.DIBUF[26].X ;
 wire \BLOCK[1].RAM32.DIBUF[27].X ;
 wire \BLOCK[1].RAM32.DIBUF[28].X ;
 wire \BLOCK[1].RAM32.DIBUF[29].X ;
 wire \BLOCK[1].RAM32.DIBUF[2].X ;
 wire \BLOCK[1].RAM32.DIBUF[30].X ;
 wire \BLOCK[1].RAM32.DIBUF[31].X ;
 wire \BLOCK[1].RAM32.DIBUF[3].X ;
 wire \BLOCK[1].RAM32.DIBUF[4].X ;
 wire \BLOCK[1].RAM32.DIBUF[5].X ;
 wire \BLOCK[1].RAM32.DIBUF[6].X ;
 wire \BLOCK[1].RAM32.DIBUF[7].X ;
 wire \BLOCK[1].RAM32.DIBUF[8].X ;
 wire \BLOCK[1].RAM32.DIBUF[9].X ;
 wire \BLOCK[1].RAM32.Do0[0] ;
 wire \BLOCK[1].RAM32.Do0[10] ;
 wire \BLOCK[1].RAM32.Do0[11] ;
 wire \BLOCK[1].RAM32.Do0[12] ;
 wire \BLOCK[1].RAM32.Do0[13] ;
 wire \BLOCK[1].RAM32.Do0[14] ;
 wire \BLOCK[1].RAM32.Do0[15] ;
 wire \BLOCK[1].RAM32.Do0[16] ;
 wire \BLOCK[1].RAM32.Do0[17] ;
 wire \BLOCK[1].RAM32.Do0[18] ;
 wire \BLOCK[1].RAM32.Do0[19] ;
 wire \BLOCK[1].RAM32.Do0[1] ;
 wire \BLOCK[1].RAM32.Do0[20] ;
 wire \BLOCK[1].RAM32.Do0[21] ;
 wire \BLOCK[1].RAM32.Do0[22] ;
 wire \BLOCK[1].RAM32.Do0[23] ;
 wire \BLOCK[1].RAM32.Do0[24] ;
 wire \BLOCK[1].RAM32.Do0[25] ;
 wire \BLOCK[1].RAM32.Do0[26] ;
 wire \BLOCK[1].RAM32.Do0[27] ;
 wire \BLOCK[1].RAM32.Do0[28] ;
 wire \BLOCK[1].RAM32.Do0[29] ;
 wire \BLOCK[1].RAM32.Do0[2] ;
 wire \BLOCK[1].RAM32.Do0[30] ;
 wire \BLOCK[1].RAM32.Do0[31] ;
 wire \BLOCK[1].RAM32.Do0[3] ;
 wire \BLOCK[1].RAM32.Do0[4] ;
 wire \BLOCK[1].RAM32.Do0[5] ;
 wire \BLOCK[1].RAM32.Do0[6] ;
 wire \BLOCK[1].RAM32.Do0[7] ;
 wire \BLOCK[1].RAM32.Do0[8] ;
 wire \BLOCK[1].RAM32.Do0[9] ;
 wire \BLOCK[1].RAM32.Do0_REG.CLKBUF[0] ;
 wire \BLOCK[1].RAM32.Do0_REG.CLKBUF[1] ;
 wire \BLOCK[1].RAM32.Do0_REG.CLKBUF[2] ;
 wire \BLOCK[1].RAM32.Do0_REG.CLKBUF[3] ;
 wire \BLOCK[1].RAM32.Do0_REG.CLK_buf ;
 wire \BLOCK[1].RAM32.EN0 ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.CLKBUF.X ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.EN ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[0].A ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[0].X ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[1].A ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[1].X ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[2].A ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[2].X ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[3].A ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[3].X ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.CLKBUF.X ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.EN ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[0].X ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[1].X ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[2].X ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[3].X ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.CLKBUF.X ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.EN ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.EN_buf ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[0].X ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[1].X ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[2].X ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[3].X ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.CLKBUF.X ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.EN ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.EN_buf ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[0].X ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[1].X ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[2].X ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[3].X ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.SEL0 ;
 wire \BLOCK[2].RAM32.A0BUF[0].X ;
 wire \BLOCK[2].RAM32.A0BUF[1].X ;
 wire \BLOCK[2].RAM32.A0BUF[2].X ;
 wire \BLOCK[2].RAM32.A0BUF[3].X ;
 wire \BLOCK[2].RAM32.A0BUF[4].X ;
 wire \BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].A ;
 wire \BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ;
 wire \BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ;
 wire \BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ;
 wire \BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ;
 wire \BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ;
 wire \BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ;
 wire \BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ;
 wire \BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ;
 wire \BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].A ;
 wire \BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].TE_B ;
 wire \BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ;
 wire \BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ;
 wire \BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ;
 wire \BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ;
 wire \BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ;
 wire \BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ;
 wire \BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ;
 wire \BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ;
 wire \BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].A ;
 wire \BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].TE_B ;
 wire \BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ;
 wire \BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ;
 wire \BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ;
 wire \BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ;
 wire \BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ;
 wire \BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ;
 wire \BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ;
 wire \BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ;
 wire \BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].A ;
 wire \BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].TE_B ;
 wire \BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ;
 wire \BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ;
 wire \BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ;
 wire \BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ;
 wire \BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ;
 wire \BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ;
 wire \BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ;
 wire \BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ;
 wire \BLOCK[2].RAM32.CLKBUF.X ;
 wire \BLOCK[2].RAM32.DEC0.EN ;
 wire \BLOCK[2].RAM32.DIBUF[0].X ;
 wire \BLOCK[2].RAM32.DIBUF[10].X ;
 wire \BLOCK[2].RAM32.DIBUF[11].X ;
 wire \BLOCK[2].RAM32.DIBUF[12].X ;
 wire \BLOCK[2].RAM32.DIBUF[13].X ;
 wire \BLOCK[2].RAM32.DIBUF[14].X ;
 wire \BLOCK[2].RAM32.DIBUF[15].X ;
 wire \BLOCK[2].RAM32.DIBUF[16].X ;
 wire \BLOCK[2].RAM32.DIBUF[17].X ;
 wire \BLOCK[2].RAM32.DIBUF[18].X ;
 wire \BLOCK[2].RAM32.DIBUF[19].X ;
 wire \BLOCK[2].RAM32.DIBUF[1].X ;
 wire \BLOCK[2].RAM32.DIBUF[20].X ;
 wire \BLOCK[2].RAM32.DIBUF[21].X ;
 wire \BLOCK[2].RAM32.DIBUF[22].X ;
 wire \BLOCK[2].RAM32.DIBUF[23].X ;
 wire \BLOCK[2].RAM32.DIBUF[24].X ;
 wire \BLOCK[2].RAM32.DIBUF[25].X ;
 wire \BLOCK[2].RAM32.DIBUF[26].X ;
 wire \BLOCK[2].RAM32.DIBUF[27].X ;
 wire \BLOCK[2].RAM32.DIBUF[28].X ;
 wire \BLOCK[2].RAM32.DIBUF[29].X ;
 wire \BLOCK[2].RAM32.DIBUF[2].X ;
 wire \BLOCK[2].RAM32.DIBUF[30].X ;
 wire \BLOCK[2].RAM32.DIBUF[31].X ;
 wire \BLOCK[2].RAM32.DIBUF[3].X ;
 wire \BLOCK[2].RAM32.DIBUF[4].X ;
 wire \BLOCK[2].RAM32.DIBUF[5].X ;
 wire \BLOCK[2].RAM32.DIBUF[6].X ;
 wire \BLOCK[2].RAM32.DIBUF[7].X ;
 wire \BLOCK[2].RAM32.DIBUF[8].X ;
 wire \BLOCK[2].RAM32.DIBUF[9].X ;
 wire \BLOCK[2].RAM32.Do0[0] ;
 wire \BLOCK[2].RAM32.Do0[10] ;
 wire \BLOCK[2].RAM32.Do0[11] ;
 wire \BLOCK[2].RAM32.Do0[12] ;
 wire \BLOCK[2].RAM32.Do0[13] ;
 wire \BLOCK[2].RAM32.Do0[14] ;
 wire \BLOCK[2].RAM32.Do0[15] ;
 wire \BLOCK[2].RAM32.Do0[16] ;
 wire \BLOCK[2].RAM32.Do0[17] ;
 wire \BLOCK[2].RAM32.Do0[18] ;
 wire \BLOCK[2].RAM32.Do0[19] ;
 wire \BLOCK[2].RAM32.Do0[1] ;
 wire \BLOCK[2].RAM32.Do0[20] ;
 wire \BLOCK[2].RAM32.Do0[21] ;
 wire \BLOCK[2].RAM32.Do0[22] ;
 wire \BLOCK[2].RAM32.Do0[23] ;
 wire \BLOCK[2].RAM32.Do0[24] ;
 wire \BLOCK[2].RAM32.Do0[25] ;
 wire \BLOCK[2].RAM32.Do0[26] ;
 wire \BLOCK[2].RAM32.Do0[27] ;
 wire \BLOCK[2].RAM32.Do0[28] ;
 wire \BLOCK[2].RAM32.Do0[29] ;
 wire \BLOCK[2].RAM32.Do0[2] ;
 wire \BLOCK[2].RAM32.Do0[30] ;
 wire \BLOCK[2].RAM32.Do0[31] ;
 wire \BLOCK[2].RAM32.Do0[3] ;
 wire \BLOCK[2].RAM32.Do0[4] ;
 wire \BLOCK[2].RAM32.Do0[5] ;
 wire \BLOCK[2].RAM32.Do0[6] ;
 wire \BLOCK[2].RAM32.Do0[7] ;
 wire \BLOCK[2].RAM32.Do0[8] ;
 wire \BLOCK[2].RAM32.Do0[9] ;
 wire \BLOCK[2].RAM32.Do0_REG.CLKBUF[0] ;
 wire \BLOCK[2].RAM32.Do0_REG.CLKBUF[1] ;
 wire \BLOCK[2].RAM32.Do0_REG.CLKBUF[2] ;
 wire \BLOCK[2].RAM32.Do0_REG.CLKBUF[3] ;
 wire \BLOCK[2].RAM32.Do0_REG.CLK_buf ;
 wire \BLOCK[2].RAM32.EN0 ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.CLKBUF.X ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.EN ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[0].A ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[0].X ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[1].A ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[1].X ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[2].A ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[2].X ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[3].A ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[3].X ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.CLKBUF.X ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.EN ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[0].X ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[1].X ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[2].X ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[3].X ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.CLKBUF.X ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.EN ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.EN_buf ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[0].X ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[1].X ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[2].X ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[3].X ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.CLKBUF.X ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.EN ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.EN_buf ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[0].X ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[1].X ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[2].X ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[3].X ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.SEL0 ;
 wire \BLOCK[3].RAM32.A0BUF[0].X ;
 wire \BLOCK[3].RAM32.A0BUF[1].X ;
 wire \BLOCK[3].RAM32.A0BUF[2].X ;
 wire \BLOCK[3].RAM32.A0BUF[3].X ;
 wire \BLOCK[3].RAM32.A0BUF[4].X ;
 wire \BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].A ;
 wire \BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].TE_B ;
 wire \BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ;
 wire \BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ;
 wire \BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ;
 wire \BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ;
 wire \BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ;
 wire \BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ;
 wire \BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ;
 wire \BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ;
 wire \BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].A ;
 wire \BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].TE_B ;
 wire \BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ;
 wire \BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ;
 wire \BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ;
 wire \BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ;
 wire \BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ;
 wire \BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ;
 wire \BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ;
 wire \BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ;
 wire \BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].A ;
 wire \BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].TE_B ;
 wire \BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ;
 wire \BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ;
 wire \BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ;
 wire \BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ;
 wire \BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ;
 wire \BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ;
 wire \BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ;
 wire \BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ;
 wire \BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].A ;
 wire \BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].TE_B ;
 wire \BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ;
 wire \BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ;
 wire \BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ;
 wire \BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ;
 wire \BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ;
 wire \BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ;
 wire \BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ;
 wire \BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ;
 wire \BLOCK[3].RAM32.CLKBUF.X ;
 wire \BLOCK[3].RAM32.DEC0.EN ;
 wire \BLOCK[3].RAM32.DIBUF[0].X ;
 wire \BLOCK[3].RAM32.DIBUF[10].X ;
 wire \BLOCK[3].RAM32.DIBUF[11].X ;
 wire \BLOCK[3].RAM32.DIBUF[12].X ;
 wire \BLOCK[3].RAM32.DIBUF[13].X ;
 wire \BLOCK[3].RAM32.DIBUF[14].X ;
 wire \BLOCK[3].RAM32.DIBUF[15].X ;
 wire \BLOCK[3].RAM32.DIBUF[16].X ;
 wire \BLOCK[3].RAM32.DIBUF[17].X ;
 wire \BLOCK[3].RAM32.DIBUF[18].X ;
 wire \BLOCK[3].RAM32.DIBUF[19].X ;
 wire \BLOCK[3].RAM32.DIBUF[1].X ;
 wire \BLOCK[3].RAM32.DIBUF[20].X ;
 wire \BLOCK[3].RAM32.DIBUF[21].X ;
 wire \BLOCK[3].RAM32.DIBUF[22].X ;
 wire \BLOCK[3].RAM32.DIBUF[23].X ;
 wire \BLOCK[3].RAM32.DIBUF[24].X ;
 wire \BLOCK[3].RAM32.DIBUF[25].X ;
 wire \BLOCK[3].RAM32.DIBUF[26].X ;
 wire \BLOCK[3].RAM32.DIBUF[27].X ;
 wire \BLOCK[3].RAM32.DIBUF[28].X ;
 wire \BLOCK[3].RAM32.DIBUF[29].X ;
 wire \BLOCK[3].RAM32.DIBUF[2].X ;
 wire \BLOCK[3].RAM32.DIBUF[30].X ;
 wire \BLOCK[3].RAM32.DIBUF[31].X ;
 wire \BLOCK[3].RAM32.DIBUF[3].X ;
 wire \BLOCK[3].RAM32.DIBUF[4].X ;
 wire \BLOCK[3].RAM32.DIBUF[5].X ;
 wire \BLOCK[3].RAM32.DIBUF[6].X ;
 wire \BLOCK[3].RAM32.DIBUF[7].X ;
 wire \BLOCK[3].RAM32.DIBUF[8].X ;
 wire \BLOCK[3].RAM32.DIBUF[9].X ;
 wire \BLOCK[3].RAM32.Do0[0] ;
 wire \BLOCK[3].RAM32.Do0[10] ;
 wire \BLOCK[3].RAM32.Do0[11] ;
 wire \BLOCK[3].RAM32.Do0[12] ;
 wire \BLOCK[3].RAM32.Do0[13] ;
 wire \BLOCK[3].RAM32.Do0[14] ;
 wire \BLOCK[3].RAM32.Do0[15] ;
 wire \BLOCK[3].RAM32.Do0[16] ;
 wire \BLOCK[3].RAM32.Do0[17] ;
 wire \BLOCK[3].RAM32.Do0[18] ;
 wire \BLOCK[3].RAM32.Do0[19] ;
 wire \BLOCK[3].RAM32.Do0[1] ;
 wire \BLOCK[3].RAM32.Do0[20] ;
 wire \BLOCK[3].RAM32.Do0[21] ;
 wire \BLOCK[3].RAM32.Do0[22] ;
 wire \BLOCK[3].RAM32.Do0[23] ;
 wire \BLOCK[3].RAM32.Do0[24] ;
 wire \BLOCK[3].RAM32.Do0[25] ;
 wire \BLOCK[3].RAM32.Do0[26] ;
 wire \BLOCK[3].RAM32.Do0[27] ;
 wire \BLOCK[3].RAM32.Do0[28] ;
 wire \BLOCK[3].RAM32.Do0[29] ;
 wire \BLOCK[3].RAM32.Do0[2] ;
 wire \BLOCK[3].RAM32.Do0[30] ;
 wire \BLOCK[3].RAM32.Do0[31] ;
 wire \BLOCK[3].RAM32.Do0[3] ;
 wire \BLOCK[3].RAM32.Do0[4] ;
 wire \BLOCK[3].RAM32.Do0[5] ;
 wire \BLOCK[3].RAM32.Do0[6] ;
 wire \BLOCK[3].RAM32.Do0[7] ;
 wire \BLOCK[3].RAM32.Do0[8] ;
 wire \BLOCK[3].RAM32.Do0[9] ;
 wire \BLOCK[3].RAM32.Do0_REG.CLKBUF[0] ;
 wire \BLOCK[3].RAM32.Do0_REG.CLKBUF[1] ;
 wire \BLOCK[3].RAM32.Do0_REG.CLKBUF[2] ;
 wire \BLOCK[3].RAM32.Do0_REG.CLKBUF[3] ;
 wire \BLOCK[3].RAM32.Do0_REG.CLK_buf ;
 wire \BLOCK[3].RAM32.EN0 ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.CLKBUF.X ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.EN ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.EN_buf ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[0].A ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[0].X ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[1].A ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[1].X ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[2].A ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[2].X ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[3].A ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[3].X ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.CLKBUF.X ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.EN ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.EN_buf ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[0].X ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[1].X ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[2].X ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[3].X ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.CLKBUF.X ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.EN ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.EN_buf ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[0].X ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[1].X ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[2].X ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[3].X ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.CLKBUF.X ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.EN ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.EN_buf ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[0].X ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[1].X ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[2].X ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[3].X ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CLK_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ;
 wire \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.SEL0 ;
 wire \DEC0.EN ;
 wire \Do0MUX.SEL0[0] ;
 wire \Do0MUX.SEL0[1] ;
 wire \Do0MUX.SEL0[2] ;
 wire \Do0MUX.SEL0[3] ;
 wire \Do0MUX.SEL1[0] ;
 wire \Do0MUX.SEL1[1] ;
 wire \Do0MUX.SEL1[2] ;
 wire \Do0MUX.SEL1[3] ;

 sky130_fd_sc_hd__clkbuf_2 \A0BUF[0].__cell__  (.A(A0[0]),
    .X(\A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \A0BUF[1].__cell__  (.A(A0[1]),
    .X(\A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \A0BUF[2].__cell__  (.A(A0[2]),
    .X(\A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \A0BUF[3].__cell__  (.A(A0[3]),
    .X(\A0BUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \A0BUF[4].__cell__  (.A(A0[4]),
    .X(\A0BUF[4].X ));
 sky130_fd_sc_hd__clkbuf_2 \A0BUF[5].__cell__  (.A(A0[5]),
    .X(\A0BUF[5].X ));
 sky130_fd_sc_hd__clkbuf_2 \A0BUF[6].__cell__  (.A(A0[6]),
    .X(\A0BUF[6].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.A0BUF[0].__cell__  (.A(\A0BUF[0].X ),
    .X(\BLOCK[0].RAM32.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.A0BUF[1].__cell__  (.A(\A0BUF[1].X ),
    .X(\BLOCK[0].RAM32.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.A0BUF[2].__cell__  (.A(\A0BUF[2].X ),
    .X(\BLOCK[0].RAM32.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.A0BUF[3].__cell__  (.A(\A0BUF[3].X ),
    .X(\BLOCK[0].RAM32.A0BUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.A0BUF[4].__cell__  (.A(\A0BUF[4].X ),
    .X(\BLOCK[0].RAM32.A0BUF[4].X ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].__cell__  (.A(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].__cell__  (.A(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].__cell__  (.A(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].__cell__  (.A(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].__cell__  (.A(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].__cell__  (.A(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].__cell__  (.A(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].__cell__  (.A(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].__cell__  (.A(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].__cell__  (.A(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].__cell__  (.A(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].__cell__  (.A(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].__cell__  (.A(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].__cell__  (.A(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].__cell__  (.A(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].__cell__  (.A(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].__cell__  (.A(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].__cell__  (.A(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].__cell__  (.A(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].__cell__  (.A(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].__cell__  (.A(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].__cell__  (.A(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].__cell__  (.A(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].__cell__  (.A(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].__cell__  (.A(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].__cell__  (.A(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].__cell__  (.A(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].__cell__  (.A(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].__cell__  (.A(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].__cell__  (.A(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].__cell__  (.A(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].__cell__  (.A(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.CLKBUF.__cell__  (.A(\BLOCK[0].RAM32.CLK ),
    .X(\BLOCK[0].RAM32.CLKBUF.X ));
 sky130_fd_sc_hd__nor3b_2 \BLOCK[0].RAM32.DEC0.AND0  (.A(\BLOCK[0].RAM32.A0BUF[3].X ),
    .B(\BLOCK[0].RAM32.A0BUF[4].X ),
    .C_N(\BLOCK[0].RAM32.DEC0.EN ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and3b_2 \BLOCK[0].RAM32.DEC0.AND1  (.A_N(\BLOCK[0].RAM32.A0BUF[4].X ),
    .B(\BLOCK[0].RAM32.A0BUF[3].X ),
    .C(\BLOCK[0].RAM32.DEC0.EN ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and3b_2 \BLOCK[0].RAM32.DEC0.AND2  (.A_N(\BLOCK[0].RAM32.A0BUF[3].X ),
    .B(\BLOCK[0].RAM32.A0BUF[4].X ),
    .C(\BLOCK[0].RAM32.DEC0.EN ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and3_2 \BLOCK[0].RAM32.DEC0.AND3  (.A(\BLOCK[0].RAM32.A0BUF[4].X ),
    .B(\BLOCK[0].RAM32.A0BUF[3].X ),
    .C(\BLOCK[0].RAM32.DEC0.EN ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[0].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[0].A ),
    .X(\BLOCK[0].RAM32.DIBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[10].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[10].A ),
    .X(\BLOCK[0].RAM32.DIBUF[10].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[11].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[11].A ),
    .X(\BLOCK[0].RAM32.DIBUF[11].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[12].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[12].A ),
    .X(\BLOCK[0].RAM32.DIBUF[12].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[13].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[13].A ),
    .X(\BLOCK[0].RAM32.DIBUF[13].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[14].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[14].A ),
    .X(\BLOCK[0].RAM32.DIBUF[14].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[15].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[15].A ),
    .X(\BLOCK[0].RAM32.DIBUF[15].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[16].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[16].A ),
    .X(\BLOCK[0].RAM32.DIBUF[16].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[17].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[17].A ),
    .X(\BLOCK[0].RAM32.DIBUF[17].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[18].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[18].A ),
    .X(\BLOCK[0].RAM32.DIBUF[18].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[19].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[19].A ),
    .X(\BLOCK[0].RAM32.DIBUF[19].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[1].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[1].A ),
    .X(\BLOCK[0].RAM32.DIBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[20].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[20].A ),
    .X(\BLOCK[0].RAM32.DIBUF[20].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[21].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[21].A ),
    .X(\BLOCK[0].RAM32.DIBUF[21].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[22].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[22].A ),
    .X(\BLOCK[0].RAM32.DIBUF[22].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[23].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[23].A ),
    .X(\BLOCK[0].RAM32.DIBUF[23].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[24].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[24].A ),
    .X(\BLOCK[0].RAM32.DIBUF[24].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[25].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[25].A ),
    .X(\BLOCK[0].RAM32.DIBUF[25].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[26].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[26].A ),
    .X(\BLOCK[0].RAM32.DIBUF[26].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[27].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[27].A ),
    .X(\BLOCK[0].RAM32.DIBUF[27].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[28].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[28].A ),
    .X(\BLOCK[0].RAM32.DIBUF[28].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[29].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[29].A ),
    .X(\BLOCK[0].RAM32.DIBUF[29].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[2].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[2].A ),
    .X(\BLOCK[0].RAM32.DIBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[30].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[30].A ),
    .X(\BLOCK[0].RAM32.DIBUF[30].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[31].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[31].A ),
    .X(\BLOCK[0].RAM32.DIBUF[31].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[3].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[3].A ),
    .X(\BLOCK[0].RAM32.DIBUF[3].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[4].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[4].A ),
    .X(\BLOCK[0].RAM32.DIBUF[4].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[5].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[5].A ),
    .X(\BLOCK[0].RAM32.DIBUF[5].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[6].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[6].A ),
    .X(\BLOCK[0].RAM32.DIBUF[6].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[7].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[7].A ),
    .X(\BLOCK[0].RAM32.DIBUF[7].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[8].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[8].A ),
    .X(\BLOCK[0].RAM32.DIBUF[8].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[0].RAM32.DIBUF[9].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[9].A ),
    .X(\BLOCK[0].RAM32.DIBUF[9].X ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.Do0_REG.Do_CLKBUF[0]  (.A(\BLOCK[0].RAM32.Do0_REG.CLK_buf ),
    .X(\BLOCK[0].RAM32.Do0_REG.CLKBUF[0] ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.Do0_REG.Do_CLKBUF[1]  (.A(\BLOCK[0].RAM32.Do0_REG.CLK_buf ),
    .X(\BLOCK[0].RAM32.Do0_REG.CLKBUF[1] ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.Do0_REG.Do_CLKBUF[2]  (.A(\BLOCK[0].RAM32.Do0_REG.CLK_buf ),
    .X(\BLOCK[0].RAM32.Do0_REG.CLKBUF[2] ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.Do0_REG.Do_CLKBUF[3]  (.A(\BLOCK[0].RAM32.Do0_REG.CLK_buf ),
    .X(\BLOCK[0].RAM32.Do0_REG.CLKBUF[3] ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ),
    .Q(\BLOCK[0].RAM32.Do0[0] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ),
    .Q(\BLOCK[0].RAM32.Do0[1] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ),
    .Q(\BLOCK[0].RAM32.Do0[2] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ),
    .Q(\BLOCK[0].RAM32.Do0[3] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ),
    .Q(\BLOCK[0].RAM32.Do0[4] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ),
    .Q(\BLOCK[0].RAM32.Do0[5] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ),
    .Q(\BLOCK[0].RAM32.Do0[6] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ),
    .Q(\BLOCK[0].RAM32.Do0[7] ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[0]  (.DIODE(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[1]  (.DIODE(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[2]  (.DIODE(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[3]  (.DIODE(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[4]  (.DIODE(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[5]  (.DIODE(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[6]  (.DIODE(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[7]  (.DIODE(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[0]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ),
    .Q(\BLOCK[0].RAM32.Do0[8] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[1]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ),
    .Q(\BLOCK[0].RAM32.Do0[9] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[2]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ),
    .Q(\BLOCK[0].RAM32.Do0[10] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[3]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ),
    .Q(\BLOCK[0].RAM32.Do0[11] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[4]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ),
    .Q(\BLOCK[0].RAM32.Do0[12] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[5]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ),
    .Q(\BLOCK[0].RAM32.Do0[13] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[6]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ),
    .Q(\BLOCK[0].RAM32.Do0[14] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[7]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ),
    .Q(\BLOCK[0].RAM32.Do0[15] ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[0]  (.DIODE(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[1]  (.DIODE(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[2]  (.DIODE(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[3]  (.DIODE(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[4]  (.DIODE(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[5]  (.DIODE(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[6]  (.DIODE(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[7]  (.DIODE(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[0]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ),
    .Q(\BLOCK[0].RAM32.Do0[16] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[1]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ),
    .Q(\BLOCK[0].RAM32.Do0[17] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[2]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ),
    .Q(\BLOCK[0].RAM32.Do0[18] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[3]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ),
    .Q(\BLOCK[0].RAM32.Do0[19] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[4]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ),
    .Q(\BLOCK[0].RAM32.Do0[20] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[5]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ),
    .Q(\BLOCK[0].RAM32.Do0[21] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[6]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ),
    .Q(\BLOCK[0].RAM32.Do0[22] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[7]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ),
    .Q(\BLOCK[0].RAM32.Do0[23] ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[0]  (.DIODE(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[1]  (.DIODE(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[2]  (.DIODE(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[3]  (.DIODE(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[4]  (.DIODE(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[5]  (.DIODE(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[6]  (.DIODE(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[7]  (.DIODE(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[0]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ),
    .Q(\BLOCK[0].RAM32.Do0[24] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[1]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ),
    .Q(\BLOCK[0].RAM32.Do0[25] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[2]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ),
    .Q(\BLOCK[0].RAM32.Do0[26] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[3]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ),
    .Q(\BLOCK[0].RAM32.Do0[27] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[4]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ),
    .Q(\BLOCK[0].RAM32.Do0[28] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[5]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ),
    .Q(\BLOCK[0].RAM32.Do0[29] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[6]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ),
    .Q(\BLOCK[0].RAM32.Do0[30] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[0].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[7]  (.CLK(\BLOCK[0].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ),
    .Q(\BLOCK[0].RAM32.Do0[31] ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.Do0_REG.Root_CLKBUF  (.A(\BLOCK[0].RAM32.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.EN0BUF.__cell__  (.A(\BLOCK[0].RAM32.EN0 ),
    .X(\BLOCK[0].RAM32.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.FBUFENBUF0[0].__cell__  (.A(\BLOCK[0].RAM32.EN0 ),
    .X(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.FBUFENBUF0[1].__cell__  (.A(\BLOCK[0].RAM32.EN0 ),
    .X(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.FBUFENBUF0[2].__cell__  (.A(\BLOCK[0].RAM32.EN0 ),
    .X(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.FBUFENBUF0[3].__cell__  (.A(\BLOCK[0].RAM32.EN0 ),
    .X(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\BLOCK[0].RAM32.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\BLOCK[0].RAM32.A0BUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\BLOCK[0].RAM32.A0BUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\BLOCK[0].RAM32.A0BUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.AND0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.AND1  (.A_N(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.AND2  (.A_N(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.AND3  (.A_N(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.AND4  (.A_N(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.AND5  (.A_N(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.AND6  (.A_N(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.AND7  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.ENBUF  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.EN ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[0].A ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[1].__cell__  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[1].A ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[2].__cell__  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[2].A ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[3].__cell__  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[3].A ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\BLOCK[0].RAM32.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\BLOCK[0].RAM32.A0BUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\BLOCK[0].RAM32.A0BUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\BLOCK[0].RAM32.A0BUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.AND0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.AND1  (.A_N(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.AND2  (.A_N(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.AND3  (.A_N(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.AND4  (.A_N(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.AND5  (.A_N(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.AND6  (.A_N(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.AND7  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.ENBUF  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.EN ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[0].A ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[1].__cell__  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[1].A ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[2].__cell__  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[2].A ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[3].__cell__  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[3].A ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[2].RAM8.CLKBUF.__cell__  (.A(\BLOCK[0].RAM32.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.ABUF[0]  (.A(\BLOCK[0].RAM32.A0BUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.ABUF[1]  (.A(\BLOCK[0].RAM32.A0BUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.ABUF[2]  (.A(\BLOCK[0].RAM32.A0BUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.AND0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D_N(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.AND1  (.A_N(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.AND2  (.A_N(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .D(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.AND3  (.A_N(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.AND4  (.A_N(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .B_N(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.AND5  (.A_N(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.AND6  (.A_N(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.AND7  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.ENBUF  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.EN ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[0].__cell__  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[0].A ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[1].__cell__  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[1].A ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[2].__cell__  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[2].A ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[3].__cell__  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[3].A ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[3].RAM8.CLKBUF.__cell__  (.A(\BLOCK[0].RAM32.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.ABUF[0]  (.A(\BLOCK[0].RAM32.A0BUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.ABUF[1]  (.A(\BLOCK[0].RAM32.A0BUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.ABUF[2]  (.A(\BLOCK[0].RAM32.A0BUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.AND0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D_N(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.AND1  (.A_N(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.AND2  (.A_N(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .D(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.AND3  (.A_N(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.AND4  (.A_N(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .B_N(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.AND5  (.A_N(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.AND6  (.A_N(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.AND7  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.ENBUF  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.EN ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[0].__cell__  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[0].A ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[1].__cell__  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[1].A ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[2].__cell__  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[2].A ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[3].__cell__  (.A(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[3].A ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[0].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[0].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.CLKBUF  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.SEL0BUF  (.A(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.SEL0 ),
    .X(\BLOCK[0].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \BLOCK[0].RAM32.TIE0[0].__cell__  (.LO(\BLOCK[0].RAM32.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__conb_1 \BLOCK[0].RAM32.TIE0[1].__cell__  (.LO(\BLOCK[0].RAM32.BYTE[1].FLOATBUF0[10].A ));
 sky130_fd_sc_hd__conb_1 \BLOCK[0].RAM32.TIE0[2].__cell__  (.LO(\BLOCK[0].RAM32.BYTE[2].FLOATBUF0[16].A ));
 sky130_fd_sc_hd__conb_1 \BLOCK[0].RAM32.TIE0[3].__cell__  (.LO(\BLOCK[0].RAM32.BYTE[3].FLOATBUF0[24].A ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.WEBUF[0].__cell__  (.A(\BLOCK[0].RAM32.WEBUF[0].A ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.WEBUF[1].__cell__  (.A(\BLOCK[0].RAM32.WEBUF[1].A ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[1].A ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.WEBUF[2].__cell__  (.A(\BLOCK[0].RAM32.WEBUF[2].A ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[2].A ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[0].RAM32.WEBUF[3].__cell__  (.A(\BLOCK[0].RAM32.WEBUF[3].A ),
    .X(\BLOCK[0].RAM32.SLICE[0].RAM8.WEBUF[3].A ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.A0BUF[0].__cell__  (.A(\A0BUF[0].X ),
    .X(\BLOCK[1].RAM32.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.A0BUF[1].__cell__  (.A(\A0BUF[1].X ),
    .X(\BLOCK[1].RAM32.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.A0BUF[2].__cell__  (.A(\A0BUF[2].X ),
    .X(\BLOCK[1].RAM32.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.A0BUF[3].__cell__  (.A(\A0BUF[3].X ),
    .X(\BLOCK[1].RAM32.A0BUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.A0BUF[4].__cell__  (.A(\A0BUF[4].X ),
    .X(\BLOCK[1].RAM32.A0BUF[4].X ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].__cell__  (.A(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].__cell__  (.A(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].__cell__  (.A(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].__cell__  (.A(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].__cell__  (.A(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].__cell__  (.A(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].__cell__  (.A(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].__cell__  (.A(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].__cell__  (.A(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].__cell__  (.A(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].__cell__  (.A(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].__cell__  (.A(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].__cell__  (.A(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].__cell__  (.A(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].__cell__  (.A(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].__cell__  (.A(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].__cell__  (.A(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].__cell__  (.A(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].__cell__  (.A(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].__cell__  (.A(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].__cell__  (.A(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].__cell__  (.A(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].__cell__  (.A(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].__cell__  (.A(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].__cell__  (.A(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].__cell__  (.A(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].__cell__  (.A(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].__cell__  (.A(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].__cell__  (.A(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].__cell__  (.A(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].__cell__  (.A(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].__cell__  (.A(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.CLKBUF.__cell__  (.A(\BLOCK[0].RAM32.CLK ),
    .X(\BLOCK[1].RAM32.CLKBUF.X ));
 sky130_fd_sc_hd__nor3b_2 \BLOCK[1].RAM32.DEC0.AND0  (.A(\BLOCK[1].RAM32.A0BUF[3].X ),
    .B(\BLOCK[1].RAM32.A0BUF[4].X ),
    .C_N(\BLOCK[1].RAM32.DEC0.EN ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and3b_2 \BLOCK[1].RAM32.DEC0.AND1  (.A_N(\BLOCK[1].RAM32.A0BUF[4].X ),
    .B(\BLOCK[1].RAM32.A0BUF[3].X ),
    .C(\BLOCK[1].RAM32.DEC0.EN ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and3b_2 \BLOCK[1].RAM32.DEC0.AND2  (.A_N(\BLOCK[1].RAM32.A0BUF[3].X ),
    .B(\BLOCK[1].RAM32.A0BUF[4].X ),
    .C(\BLOCK[1].RAM32.DEC0.EN ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and3_2 \BLOCK[1].RAM32.DEC0.AND3  (.A(\BLOCK[1].RAM32.A0BUF[4].X ),
    .B(\BLOCK[1].RAM32.A0BUF[3].X ),
    .C(\BLOCK[1].RAM32.DEC0.EN ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[0].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[0].A ),
    .X(\BLOCK[1].RAM32.DIBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[10].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[10].A ),
    .X(\BLOCK[1].RAM32.DIBUF[10].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[11].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[11].A ),
    .X(\BLOCK[1].RAM32.DIBUF[11].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[12].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[12].A ),
    .X(\BLOCK[1].RAM32.DIBUF[12].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[13].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[13].A ),
    .X(\BLOCK[1].RAM32.DIBUF[13].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[14].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[14].A ),
    .X(\BLOCK[1].RAM32.DIBUF[14].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[15].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[15].A ),
    .X(\BLOCK[1].RAM32.DIBUF[15].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[16].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[16].A ),
    .X(\BLOCK[1].RAM32.DIBUF[16].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[17].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[17].A ),
    .X(\BLOCK[1].RAM32.DIBUF[17].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[18].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[18].A ),
    .X(\BLOCK[1].RAM32.DIBUF[18].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[19].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[19].A ),
    .X(\BLOCK[1].RAM32.DIBUF[19].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[1].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[1].A ),
    .X(\BLOCK[1].RAM32.DIBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[20].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[20].A ),
    .X(\BLOCK[1].RAM32.DIBUF[20].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[21].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[21].A ),
    .X(\BLOCK[1].RAM32.DIBUF[21].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[22].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[22].A ),
    .X(\BLOCK[1].RAM32.DIBUF[22].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[23].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[23].A ),
    .X(\BLOCK[1].RAM32.DIBUF[23].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[24].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[24].A ),
    .X(\BLOCK[1].RAM32.DIBUF[24].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[25].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[25].A ),
    .X(\BLOCK[1].RAM32.DIBUF[25].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[26].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[26].A ),
    .X(\BLOCK[1].RAM32.DIBUF[26].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[27].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[27].A ),
    .X(\BLOCK[1].RAM32.DIBUF[27].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[28].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[28].A ),
    .X(\BLOCK[1].RAM32.DIBUF[28].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[29].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[29].A ),
    .X(\BLOCK[1].RAM32.DIBUF[29].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[2].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[2].A ),
    .X(\BLOCK[1].RAM32.DIBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[30].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[30].A ),
    .X(\BLOCK[1].RAM32.DIBUF[30].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[31].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[31].A ),
    .X(\BLOCK[1].RAM32.DIBUF[31].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[3].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[3].A ),
    .X(\BLOCK[1].RAM32.DIBUF[3].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[4].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[4].A ),
    .X(\BLOCK[1].RAM32.DIBUF[4].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[5].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[5].A ),
    .X(\BLOCK[1].RAM32.DIBUF[5].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[6].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[6].A ),
    .X(\BLOCK[1].RAM32.DIBUF[6].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[7].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[7].A ),
    .X(\BLOCK[1].RAM32.DIBUF[7].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[8].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[8].A ),
    .X(\BLOCK[1].RAM32.DIBUF[8].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[1].RAM32.DIBUF[9].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[9].A ),
    .X(\BLOCK[1].RAM32.DIBUF[9].X ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.Do0_REG.Do_CLKBUF[0]  (.A(\BLOCK[1].RAM32.Do0_REG.CLK_buf ),
    .X(\BLOCK[1].RAM32.Do0_REG.CLKBUF[0] ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.Do0_REG.Do_CLKBUF[1]  (.A(\BLOCK[1].RAM32.Do0_REG.CLK_buf ),
    .X(\BLOCK[1].RAM32.Do0_REG.CLKBUF[1] ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.Do0_REG.Do_CLKBUF[2]  (.A(\BLOCK[1].RAM32.Do0_REG.CLK_buf ),
    .X(\BLOCK[1].RAM32.Do0_REG.CLKBUF[2] ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.Do0_REG.Do_CLKBUF[3]  (.A(\BLOCK[1].RAM32.Do0_REG.CLK_buf ),
    .X(\BLOCK[1].RAM32.Do0_REG.CLKBUF[3] ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ),
    .Q(\BLOCK[1].RAM32.Do0[0] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ),
    .Q(\BLOCK[1].RAM32.Do0[1] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ),
    .Q(\BLOCK[1].RAM32.Do0[2] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ),
    .Q(\BLOCK[1].RAM32.Do0[3] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ),
    .Q(\BLOCK[1].RAM32.Do0[4] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ),
    .Q(\BLOCK[1].RAM32.Do0[5] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ),
    .Q(\BLOCK[1].RAM32.Do0[6] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ),
    .Q(\BLOCK[1].RAM32.Do0[7] ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[0]  (.DIODE(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[1]  (.DIODE(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[2]  (.DIODE(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[3]  (.DIODE(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[4]  (.DIODE(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[5]  (.DIODE(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[6]  (.DIODE(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[7]  (.DIODE(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[0]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ),
    .Q(\BLOCK[1].RAM32.Do0[8] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[1]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ),
    .Q(\BLOCK[1].RAM32.Do0[9] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[2]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ),
    .Q(\BLOCK[1].RAM32.Do0[10] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[3]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ),
    .Q(\BLOCK[1].RAM32.Do0[11] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[4]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ),
    .Q(\BLOCK[1].RAM32.Do0[12] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[5]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ),
    .Q(\BLOCK[1].RAM32.Do0[13] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[6]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ),
    .Q(\BLOCK[1].RAM32.Do0[14] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[7]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ),
    .Q(\BLOCK[1].RAM32.Do0[15] ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[0]  (.DIODE(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[1]  (.DIODE(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[2]  (.DIODE(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[3]  (.DIODE(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[4]  (.DIODE(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[5]  (.DIODE(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[6]  (.DIODE(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[7]  (.DIODE(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[0]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ),
    .Q(\BLOCK[1].RAM32.Do0[16] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[1]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ),
    .Q(\BLOCK[1].RAM32.Do0[17] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[2]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ),
    .Q(\BLOCK[1].RAM32.Do0[18] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[3]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ),
    .Q(\BLOCK[1].RAM32.Do0[19] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[4]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ),
    .Q(\BLOCK[1].RAM32.Do0[20] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[5]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ),
    .Q(\BLOCK[1].RAM32.Do0[21] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[6]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ),
    .Q(\BLOCK[1].RAM32.Do0[22] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[7]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ),
    .Q(\BLOCK[1].RAM32.Do0[23] ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[0]  (.DIODE(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[1]  (.DIODE(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[2]  (.DIODE(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[3]  (.DIODE(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[4]  (.DIODE(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[5]  (.DIODE(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[6]  (.DIODE(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[7]  (.DIODE(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[0]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ),
    .Q(\BLOCK[1].RAM32.Do0[24] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[1]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ),
    .Q(\BLOCK[1].RAM32.Do0[25] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[2]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ),
    .Q(\BLOCK[1].RAM32.Do0[26] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[3]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ),
    .Q(\BLOCK[1].RAM32.Do0[27] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[4]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ),
    .Q(\BLOCK[1].RAM32.Do0[28] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[5]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ),
    .Q(\BLOCK[1].RAM32.Do0[29] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[6]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ),
    .Q(\BLOCK[1].RAM32.Do0[30] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[1].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[7]  (.CLK(\BLOCK[1].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ),
    .Q(\BLOCK[1].RAM32.Do0[31] ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.Do0_REG.Root_CLKBUF  (.A(\BLOCK[1].RAM32.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.EN0BUF.__cell__  (.A(\BLOCK[1].RAM32.EN0 ),
    .X(\BLOCK[1].RAM32.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.FBUFENBUF0[0].__cell__  (.A(\BLOCK[1].RAM32.EN0 ),
    .X(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.FBUFENBUF0[1].__cell__  (.A(\BLOCK[1].RAM32.EN0 ),
    .X(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.FBUFENBUF0[2].__cell__  (.A(\BLOCK[1].RAM32.EN0 ),
    .X(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.FBUFENBUF0[3].__cell__  (.A(\BLOCK[1].RAM32.EN0 ),
    .X(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\BLOCK[1].RAM32.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\BLOCK[1].RAM32.A0BUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\BLOCK[1].RAM32.A0BUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\BLOCK[1].RAM32.A0BUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.AND0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.AND1  (.A_N(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.AND2  (.A_N(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.AND3  (.A_N(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.AND4  (.A_N(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.AND5  (.A_N(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.AND6  (.A_N(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.AND7  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.ENBUF  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.EN ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[0].A ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[1].__cell__  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[1].A ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[2].__cell__  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[2].A ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[3].__cell__  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[3].A ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\BLOCK[1].RAM32.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\BLOCK[1].RAM32.A0BUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\BLOCK[1].RAM32.A0BUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\BLOCK[1].RAM32.A0BUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.AND0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.AND1  (.A_N(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.AND2  (.A_N(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.AND3  (.A_N(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.AND4  (.A_N(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.AND5  (.A_N(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.AND6  (.A_N(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.AND7  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.ENBUF  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.EN ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[0].A ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[1].__cell__  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[1].A ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[2].__cell__  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[2].A ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[3].__cell__  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[3].A ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[2].RAM8.CLKBUF.__cell__  (.A(\BLOCK[1].RAM32.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.ABUF[0]  (.A(\BLOCK[1].RAM32.A0BUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.ABUF[1]  (.A(\BLOCK[1].RAM32.A0BUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.ABUF[2]  (.A(\BLOCK[1].RAM32.A0BUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.AND0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D_N(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.AND1  (.A_N(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.AND2  (.A_N(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .D(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.AND3  (.A_N(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.AND4  (.A_N(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .B_N(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.AND5  (.A_N(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.AND6  (.A_N(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.AND7  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.ENBUF  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.EN ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[0].__cell__  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[0].A ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[1].__cell__  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[1].A ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[2].__cell__  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[2].A ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[3].__cell__  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[3].A ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[3].RAM8.CLKBUF.__cell__  (.A(\BLOCK[1].RAM32.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.ABUF[0]  (.A(\BLOCK[1].RAM32.A0BUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.ABUF[1]  (.A(\BLOCK[1].RAM32.A0BUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.ABUF[2]  (.A(\BLOCK[1].RAM32.A0BUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.AND0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D_N(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.AND1  (.A_N(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.AND2  (.A_N(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .D(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.AND3  (.A_N(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.AND4  (.A_N(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .B_N(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.AND5  (.A_N(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.AND6  (.A_N(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.AND7  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.ENBUF  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.EN ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[0].__cell__  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[0].A ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[1].__cell__  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[1].A ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[2].__cell__  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[2].A ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[3].__cell__  (.A(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[3].A ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[1].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[1].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.CLKBUF  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.SEL0BUF  (.A(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.SEL0 ),
    .X(\BLOCK[1].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \BLOCK[1].RAM32.TIE0[0].__cell__  (.LO(\BLOCK[1].RAM32.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__conb_1 \BLOCK[1].RAM32.TIE0[1].__cell__  (.LO(\BLOCK[1].RAM32.BYTE[1].FLOATBUF0[10].A ));
 sky130_fd_sc_hd__conb_1 \BLOCK[1].RAM32.TIE0[2].__cell__  (.LO(\BLOCK[1].RAM32.BYTE[2].FLOATBUF0[16].A ));
 sky130_fd_sc_hd__conb_1 \BLOCK[1].RAM32.TIE0[3].__cell__  (.LO(\BLOCK[1].RAM32.BYTE[3].FLOATBUF0[24].A ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.WEBUF[0].__cell__  (.A(\BLOCK[0].RAM32.WEBUF[0].A ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.WEBUF[1].__cell__  (.A(\BLOCK[0].RAM32.WEBUF[1].A ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[1].A ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.WEBUF[2].__cell__  (.A(\BLOCK[0].RAM32.WEBUF[2].A ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[2].A ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[1].RAM32.WEBUF[3].__cell__  (.A(\BLOCK[0].RAM32.WEBUF[3].A ),
    .X(\BLOCK[1].RAM32.SLICE[0].RAM8.WEBUF[3].A ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.A0BUF[0].__cell__  (.A(\A0BUF[0].X ),
    .X(\BLOCK[2].RAM32.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.A0BUF[1].__cell__  (.A(\A0BUF[1].X ),
    .X(\BLOCK[2].RAM32.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.A0BUF[2].__cell__  (.A(\A0BUF[2].X ),
    .X(\BLOCK[2].RAM32.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.A0BUF[3].__cell__  (.A(\A0BUF[3].X ),
    .X(\BLOCK[2].RAM32.A0BUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.A0BUF[4].__cell__  (.A(\A0BUF[4].X ),
    .X(\BLOCK[2].RAM32.A0BUF[4].X ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].__cell__  (.A(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].__cell__  (.A(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].__cell__  (.A(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].__cell__  (.A(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].__cell__  (.A(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].__cell__  (.A(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].__cell__  (.A(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].__cell__  (.A(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].__cell__  (.A(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].__cell__  (.A(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].__cell__  (.A(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].__cell__  (.A(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].__cell__  (.A(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].__cell__  (.A(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].__cell__  (.A(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].__cell__  (.A(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].__cell__  (.A(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].__cell__  (.A(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].__cell__  (.A(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].__cell__  (.A(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].__cell__  (.A(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].__cell__  (.A(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].__cell__  (.A(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].__cell__  (.A(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].__cell__  (.A(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].__cell__  (.A(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].__cell__  (.A(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].__cell__  (.A(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].__cell__  (.A(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].__cell__  (.A(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].__cell__  (.A(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].__cell__  (.A(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.CLKBUF.__cell__  (.A(\BLOCK[0].RAM32.CLK ),
    .X(\BLOCK[2].RAM32.CLKBUF.X ));
 sky130_fd_sc_hd__nor3b_2 \BLOCK[2].RAM32.DEC0.AND0  (.A(\BLOCK[2].RAM32.A0BUF[3].X ),
    .B(\BLOCK[2].RAM32.A0BUF[4].X ),
    .C_N(\BLOCK[2].RAM32.DEC0.EN ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and3b_2 \BLOCK[2].RAM32.DEC0.AND1  (.A_N(\BLOCK[2].RAM32.A0BUF[4].X ),
    .B(\BLOCK[2].RAM32.A0BUF[3].X ),
    .C(\BLOCK[2].RAM32.DEC0.EN ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and3b_2 \BLOCK[2].RAM32.DEC0.AND2  (.A_N(\BLOCK[2].RAM32.A0BUF[3].X ),
    .B(\BLOCK[2].RAM32.A0BUF[4].X ),
    .C(\BLOCK[2].RAM32.DEC0.EN ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and3_2 \BLOCK[2].RAM32.DEC0.AND3  (.A(\BLOCK[2].RAM32.A0BUF[4].X ),
    .B(\BLOCK[2].RAM32.A0BUF[3].X ),
    .C(\BLOCK[2].RAM32.DEC0.EN ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[0].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[0].A ),
    .X(\BLOCK[2].RAM32.DIBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[10].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[10].A ),
    .X(\BLOCK[2].RAM32.DIBUF[10].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[11].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[11].A ),
    .X(\BLOCK[2].RAM32.DIBUF[11].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[12].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[12].A ),
    .X(\BLOCK[2].RAM32.DIBUF[12].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[13].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[13].A ),
    .X(\BLOCK[2].RAM32.DIBUF[13].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[14].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[14].A ),
    .X(\BLOCK[2].RAM32.DIBUF[14].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[15].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[15].A ),
    .X(\BLOCK[2].RAM32.DIBUF[15].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[16].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[16].A ),
    .X(\BLOCK[2].RAM32.DIBUF[16].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[17].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[17].A ),
    .X(\BLOCK[2].RAM32.DIBUF[17].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[18].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[18].A ),
    .X(\BLOCK[2].RAM32.DIBUF[18].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[19].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[19].A ),
    .X(\BLOCK[2].RAM32.DIBUF[19].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[1].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[1].A ),
    .X(\BLOCK[2].RAM32.DIBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[20].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[20].A ),
    .X(\BLOCK[2].RAM32.DIBUF[20].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[21].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[21].A ),
    .X(\BLOCK[2].RAM32.DIBUF[21].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[22].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[22].A ),
    .X(\BLOCK[2].RAM32.DIBUF[22].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[23].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[23].A ),
    .X(\BLOCK[2].RAM32.DIBUF[23].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[24].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[24].A ),
    .X(\BLOCK[2].RAM32.DIBUF[24].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[25].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[25].A ),
    .X(\BLOCK[2].RAM32.DIBUF[25].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[26].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[26].A ),
    .X(\BLOCK[2].RAM32.DIBUF[26].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[27].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[27].A ),
    .X(\BLOCK[2].RAM32.DIBUF[27].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[28].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[28].A ),
    .X(\BLOCK[2].RAM32.DIBUF[28].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[29].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[29].A ),
    .X(\BLOCK[2].RAM32.DIBUF[29].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[2].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[2].A ),
    .X(\BLOCK[2].RAM32.DIBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[30].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[30].A ),
    .X(\BLOCK[2].RAM32.DIBUF[30].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[31].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[31].A ),
    .X(\BLOCK[2].RAM32.DIBUF[31].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[3].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[3].A ),
    .X(\BLOCK[2].RAM32.DIBUF[3].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[4].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[4].A ),
    .X(\BLOCK[2].RAM32.DIBUF[4].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[5].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[5].A ),
    .X(\BLOCK[2].RAM32.DIBUF[5].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[6].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[6].A ),
    .X(\BLOCK[2].RAM32.DIBUF[6].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[7].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[7].A ),
    .X(\BLOCK[2].RAM32.DIBUF[7].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[8].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[8].A ),
    .X(\BLOCK[2].RAM32.DIBUF[8].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[2].RAM32.DIBUF[9].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[9].A ),
    .X(\BLOCK[2].RAM32.DIBUF[9].X ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.Do0_REG.Do_CLKBUF[0]  (.A(\BLOCK[2].RAM32.Do0_REG.CLK_buf ),
    .X(\BLOCK[2].RAM32.Do0_REG.CLKBUF[0] ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.Do0_REG.Do_CLKBUF[1]  (.A(\BLOCK[2].RAM32.Do0_REG.CLK_buf ),
    .X(\BLOCK[2].RAM32.Do0_REG.CLKBUF[1] ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.Do0_REG.Do_CLKBUF[2]  (.A(\BLOCK[2].RAM32.Do0_REG.CLK_buf ),
    .X(\BLOCK[2].RAM32.Do0_REG.CLKBUF[2] ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.Do0_REG.Do_CLKBUF[3]  (.A(\BLOCK[2].RAM32.Do0_REG.CLK_buf ),
    .X(\BLOCK[2].RAM32.Do0_REG.CLKBUF[3] ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ),
    .Q(\BLOCK[2].RAM32.Do0[0] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ),
    .Q(\BLOCK[2].RAM32.Do0[1] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ),
    .Q(\BLOCK[2].RAM32.Do0[2] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ),
    .Q(\BLOCK[2].RAM32.Do0[3] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ),
    .Q(\BLOCK[2].RAM32.Do0[4] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ),
    .Q(\BLOCK[2].RAM32.Do0[5] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ),
    .Q(\BLOCK[2].RAM32.Do0[6] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ),
    .Q(\BLOCK[2].RAM32.Do0[7] ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[0]  (.DIODE(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[1]  (.DIODE(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[2]  (.DIODE(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[3]  (.DIODE(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[4]  (.DIODE(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[5]  (.DIODE(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[6]  (.DIODE(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[7]  (.DIODE(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[0]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ),
    .Q(\BLOCK[2].RAM32.Do0[8] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[1]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ),
    .Q(\BLOCK[2].RAM32.Do0[9] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[2]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ),
    .Q(\BLOCK[2].RAM32.Do0[10] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[3]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ),
    .Q(\BLOCK[2].RAM32.Do0[11] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[4]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ),
    .Q(\BLOCK[2].RAM32.Do0[12] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[5]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ),
    .Q(\BLOCK[2].RAM32.Do0[13] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[6]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ),
    .Q(\BLOCK[2].RAM32.Do0[14] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[7]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ),
    .Q(\BLOCK[2].RAM32.Do0[15] ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[0]  (.DIODE(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[1]  (.DIODE(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[2]  (.DIODE(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[3]  (.DIODE(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[4]  (.DIODE(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[5]  (.DIODE(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[6]  (.DIODE(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[7]  (.DIODE(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[0]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ),
    .Q(\BLOCK[2].RAM32.Do0[16] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[1]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ),
    .Q(\BLOCK[2].RAM32.Do0[17] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[2]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ),
    .Q(\BLOCK[2].RAM32.Do0[18] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[3]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ),
    .Q(\BLOCK[2].RAM32.Do0[19] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[4]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ),
    .Q(\BLOCK[2].RAM32.Do0[20] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[5]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ),
    .Q(\BLOCK[2].RAM32.Do0[21] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[6]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ),
    .Q(\BLOCK[2].RAM32.Do0[22] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[7]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ),
    .Q(\BLOCK[2].RAM32.Do0[23] ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[0]  (.DIODE(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[1]  (.DIODE(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[2]  (.DIODE(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[3]  (.DIODE(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[4]  (.DIODE(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[5]  (.DIODE(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[6]  (.DIODE(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[7]  (.DIODE(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[0]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ),
    .Q(\BLOCK[2].RAM32.Do0[24] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[1]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ),
    .Q(\BLOCK[2].RAM32.Do0[25] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[2]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ),
    .Q(\BLOCK[2].RAM32.Do0[26] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[3]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ),
    .Q(\BLOCK[2].RAM32.Do0[27] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[4]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ),
    .Q(\BLOCK[2].RAM32.Do0[28] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[5]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ),
    .Q(\BLOCK[2].RAM32.Do0[29] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[6]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ),
    .Q(\BLOCK[2].RAM32.Do0[30] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[2].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[7]  (.CLK(\BLOCK[2].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ),
    .Q(\BLOCK[2].RAM32.Do0[31] ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.Do0_REG.Root_CLKBUF  (.A(\BLOCK[2].RAM32.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.EN0BUF.__cell__  (.A(\BLOCK[2].RAM32.EN0 ),
    .X(\BLOCK[2].RAM32.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.FBUFENBUF0[0].__cell__  (.A(\BLOCK[2].RAM32.EN0 ),
    .X(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.FBUFENBUF0[1].__cell__  (.A(\BLOCK[2].RAM32.EN0 ),
    .X(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.FBUFENBUF0[2].__cell__  (.A(\BLOCK[2].RAM32.EN0 ),
    .X(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.FBUFENBUF0[3].__cell__  (.A(\BLOCK[2].RAM32.EN0 ),
    .X(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\BLOCK[2].RAM32.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\BLOCK[2].RAM32.A0BUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\BLOCK[2].RAM32.A0BUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\BLOCK[2].RAM32.A0BUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.AND0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.AND1  (.A_N(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.AND2  (.A_N(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.AND3  (.A_N(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.AND4  (.A_N(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.AND5  (.A_N(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.AND6  (.A_N(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.AND7  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.ENBUF  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.EN ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[0].A ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[1].__cell__  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[1].A ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[2].__cell__  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[2].A ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[3].__cell__  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[3].A ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\BLOCK[2].RAM32.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\BLOCK[2].RAM32.A0BUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\BLOCK[2].RAM32.A0BUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\BLOCK[2].RAM32.A0BUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.AND0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.AND1  (.A_N(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.AND2  (.A_N(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.AND3  (.A_N(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.AND4  (.A_N(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.AND5  (.A_N(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.AND6  (.A_N(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.AND7  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.ENBUF  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.EN ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[0].A ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[1].__cell__  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[1].A ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[2].__cell__  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[2].A ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[3].__cell__  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[3].A ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[2].RAM8.CLKBUF.__cell__  (.A(\BLOCK[2].RAM32.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.ABUF[0]  (.A(\BLOCK[2].RAM32.A0BUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.ABUF[1]  (.A(\BLOCK[2].RAM32.A0BUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.ABUF[2]  (.A(\BLOCK[2].RAM32.A0BUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.AND0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D_N(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.AND1  (.A_N(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.AND2  (.A_N(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .D(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.AND3  (.A_N(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.AND4  (.A_N(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .B_N(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.AND5  (.A_N(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.AND6  (.A_N(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.AND7  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.ENBUF  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.EN ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[0].__cell__  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[0].A ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[1].__cell__  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[1].A ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[2].__cell__  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[2].A ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[3].__cell__  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[3].A ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[3].RAM8.CLKBUF.__cell__  (.A(\BLOCK[2].RAM32.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.ABUF[0]  (.A(\BLOCK[2].RAM32.A0BUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.ABUF[1]  (.A(\BLOCK[2].RAM32.A0BUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.ABUF[2]  (.A(\BLOCK[2].RAM32.A0BUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.AND0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D_N(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.AND1  (.A_N(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.AND2  (.A_N(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .D(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.AND3  (.A_N(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.AND4  (.A_N(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .B_N(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.AND5  (.A_N(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.AND6  (.A_N(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.AND7  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.ENBUF  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.EN ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[0].__cell__  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[0].A ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[1].__cell__  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[1].A ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[2].__cell__  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[2].A ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[3].__cell__  (.A(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[3].A ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[2].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[2].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.CLKBUF  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.SEL0BUF  (.A(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.SEL0 ),
    .X(\BLOCK[2].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \BLOCK[2].RAM32.TIE0[0].__cell__  (.LO(\BLOCK[2].RAM32.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__conb_1 \BLOCK[2].RAM32.TIE0[1].__cell__  (.LO(\BLOCK[2].RAM32.BYTE[1].FLOATBUF0[10].A ));
 sky130_fd_sc_hd__conb_1 \BLOCK[2].RAM32.TIE0[2].__cell__  (.LO(\BLOCK[2].RAM32.BYTE[2].FLOATBUF0[16].A ));
 sky130_fd_sc_hd__conb_1 \BLOCK[2].RAM32.TIE0[3].__cell__  (.LO(\BLOCK[2].RAM32.BYTE[3].FLOATBUF0[24].A ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.WEBUF[0].__cell__  (.A(\BLOCK[0].RAM32.WEBUF[0].A ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.WEBUF[1].__cell__  (.A(\BLOCK[0].RAM32.WEBUF[1].A ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[1].A ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.WEBUF[2].__cell__  (.A(\BLOCK[0].RAM32.WEBUF[2].A ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[2].A ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[2].RAM32.WEBUF[3].__cell__  (.A(\BLOCK[0].RAM32.WEBUF[3].A ),
    .X(\BLOCK[2].RAM32.SLICE[0].RAM8.WEBUF[3].A ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.A0BUF[0].__cell__  (.A(\A0BUF[0].X ),
    .X(\BLOCK[3].RAM32.A0BUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.A0BUF[1].__cell__  (.A(\A0BUF[1].X ),
    .X(\BLOCK[3].RAM32.A0BUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.A0BUF[2].__cell__  (.A(\A0BUF[2].X ),
    .X(\BLOCK[3].RAM32.A0BUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.A0BUF[3].__cell__  (.A(\A0BUF[3].X ),
    .X(\BLOCK[3].RAM32.A0BUF[3].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.A0BUF[4].__cell__  (.A(\A0BUF[4].X ),
    .X(\BLOCK[3].RAM32.A0BUF[4].X ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].__cell__  (.A(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].__cell__  (.A(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].__cell__  (.A(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].__cell__  (.A(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].__cell__  (.A(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].__cell__  (.A(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].__cell__  (.A(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].__cell__  (.A(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].__cell__  (.A(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].__cell__  (.A(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].__cell__  (.A(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].__cell__  (.A(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].__cell__  (.A(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].__cell__  (.A(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].__cell__  (.A(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].__cell__  (.A(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].__cell__  (.A(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].__cell__  (.A(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].__cell__  (.A(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].__cell__  (.A(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].__cell__  (.A(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].__cell__  (.A(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].__cell__  (.A(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].__cell__  (.A(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].__cell__  (.A(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].__cell__  (.A(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].__cell__  (.A(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].__cell__  (.A(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].__cell__  (.A(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].__cell__  (.A(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].__cell__  (.A(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].__cell__  (.A(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].A ),
    .TE_B(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].TE_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.CLKBUF.__cell__  (.A(\BLOCK[0].RAM32.CLK ),
    .X(\BLOCK[3].RAM32.CLKBUF.X ));
 sky130_fd_sc_hd__nor3b_2 \BLOCK[3].RAM32.DEC0.AND0  (.A(\BLOCK[3].RAM32.A0BUF[3].X ),
    .B(\BLOCK[3].RAM32.A0BUF[4].X ),
    .C_N(\BLOCK[3].RAM32.DEC0.EN ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and3b_2 \BLOCK[3].RAM32.DEC0.AND1  (.A_N(\BLOCK[3].RAM32.A0BUF[4].X ),
    .B(\BLOCK[3].RAM32.A0BUF[3].X ),
    .C(\BLOCK[3].RAM32.DEC0.EN ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and3b_2 \BLOCK[3].RAM32.DEC0.AND2  (.A_N(\BLOCK[3].RAM32.A0BUF[3].X ),
    .B(\BLOCK[3].RAM32.A0BUF[4].X ),
    .C(\BLOCK[3].RAM32.DEC0.EN ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__and3_2 \BLOCK[3].RAM32.DEC0.AND3  (.A(\BLOCK[3].RAM32.A0BUF[4].X ),
    .B(\BLOCK[3].RAM32.A0BUF[3].X ),
    .C(\BLOCK[3].RAM32.DEC0.EN ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[0].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[0].A ),
    .X(\BLOCK[3].RAM32.DIBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[10].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[10].A ),
    .X(\BLOCK[3].RAM32.DIBUF[10].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[11].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[11].A ),
    .X(\BLOCK[3].RAM32.DIBUF[11].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[12].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[12].A ),
    .X(\BLOCK[3].RAM32.DIBUF[12].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[13].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[13].A ),
    .X(\BLOCK[3].RAM32.DIBUF[13].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[14].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[14].A ),
    .X(\BLOCK[3].RAM32.DIBUF[14].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[15].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[15].A ),
    .X(\BLOCK[3].RAM32.DIBUF[15].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[16].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[16].A ),
    .X(\BLOCK[3].RAM32.DIBUF[16].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[17].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[17].A ),
    .X(\BLOCK[3].RAM32.DIBUF[17].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[18].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[18].A ),
    .X(\BLOCK[3].RAM32.DIBUF[18].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[19].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[19].A ),
    .X(\BLOCK[3].RAM32.DIBUF[19].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[1].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[1].A ),
    .X(\BLOCK[3].RAM32.DIBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[20].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[20].A ),
    .X(\BLOCK[3].RAM32.DIBUF[20].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[21].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[21].A ),
    .X(\BLOCK[3].RAM32.DIBUF[21].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[22].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[22].A ),
    .X(\BLOCK[3].RAM32.DIBUF[22].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[23].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[23].A ),
    .X(\BLOCK[3].RAM32.DIBUF[23].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[24].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[24].A ),
    .X(\BLOCK[3].RAM32.DIBUF[24].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[25].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[25].A ),
    .X(\BLOCK[3].RAM32.DIBUF[25].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[26].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[26].A ),
    .X(\BLOCK[3].RAM32.DIBUF[26].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[27].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[27].A ),
    .X(\BLOCK[3].RAM32.DIBUF[27].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[28].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[28].A ),
    .X(\BLOCK[3].RAM32.DIBUF[28].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[29].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[29].A ),
    .X(\BLOCK[3].RAM32.DIBUF[29].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[2].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[2].A ),
    .X(\BLOCK[3].RAM32.DIBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[30].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[30].A ),
    .X(\BLOCK[3].RAM32.DIBUF[30].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[31].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[31].A ),
    .X(\BLOCK[3].RAM32.DIBUF[31].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[3].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[3].A ),
    .X(\BLOCK[3].RAM32.DIBUF[3].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[4].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[4].A ),
    .X(\BLOCK[3].RAM32.DIBUF[4].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[5].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[5].A ),
    .X(\BLOCK[3].RAM32.DIBUF[5].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[6].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[6].A ),
    .X(\BLOCK[3].RAM32.DIBUF[6].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[7].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[7].A ),
    .X(\BLOCK[3].RAM32.DIBUF[7].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[8].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[8].A ),
    .X(\BLOCK[3].RAM32.DIBUF[8].X ));
 sky130_fd_sc_hd__clkbuf_16 \BLOCK[3].RAM32.DIBUF[9].__cell__  (.A(\BLOCK[0].RAM32.DIBUF[9].A ),
    .X(\BLOCK[3].RAM32.DIBUF[9].X ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.Do0_REG.Do_CLKBUF[0]  (.A(\BLOCK[3].RAM32.Do0_REG.CLK_buf ),
    .X(\BLOCK[3].RAM32.Do0_REG.CLKBUF[0] ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.Do0_REG.Do_CLKBUF[1]  (.A(\BLOCK[3].RAM32.Do0_REG.CLK_buf ),
    .X(\BLOCK[3].RAM32.Do0_REG.CLKBUF[1] ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.Do0_REG.Do_CLKBUF[2]  (.A(\BLOCK[3].RAM32.Do0_REG.CLK_buf ),
    .X(\BLOCK[3].RAM32.Do0_REG.CLKBUF[2] ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.Do0_REG.Do_CLKBUF[3]  (.A(\BLOCK[3].RAM32.Do0_REG.CLK_buf ),
    .X(\BLOCK[3].RAM32.Do0_REG.CLKBUF[3] ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[0]  (.DIODE(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[1]  (.DIODE(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[2]  (.DIODE(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[3]  (.DIODE(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[4]  (.DIODE(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[5]  (.DIODE(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[6]  (.DIODE(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[0].DIODE[7]  (.DIODE(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[0]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ),
    .Q(\BLOCK[3].RAM32.Do0[0] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[1]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ),
    .Q(\BLOCK[3].RAM32.Do0[1] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[2]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ),
    .Q(\BLOCK[3].RAM32.Do0[2] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[3]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ),
    .Q(\BLOCK[3].RAM32.Do0[3] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[4]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ),
    .Q(\BLOCK[3].RAM32.Do0[4] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[5]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ),
    .Q(\BLOCK[3].RAM32.Do0[5] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[6]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ),
    .Q(\BLOCK[3].RAM32.Do0[6] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[0].Do_FF[7]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[0] ),
    .D(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ),
    .Q(\BLOCK[3].RAM32.Do0[7] ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[0]  (.DIODE(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[1]  (.DIODE(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[2]  (.DIODE(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[3]  (.DIODE(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[4]  (.DIODE(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[5]  (.DIODE(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[6]  (.DIODE(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[1].DIODE[7]  (.DIODE(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[0]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ),
    .Q(\BLOCK[3].RAM32.Do0[8] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[1]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ),
    .Q(\BLOCK[3].RAM32.Do0[9] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[2]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ),
    .Q(\BLOCK[3].RAM32.Do0[10] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[3]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ),
    .Q(\BLOCK[3].RAM32.Do0[11] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[4]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ),
    .Q(\BLOCK[3].RAM32.Do0[12] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[5]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ),
    .Q(\BLOCK[3].RAM32.Do0[13] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[6]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ),
    .Q(\BLOCK[3].RAM32.Do0[14] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[1].Do_FF[7]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[1] ),
    .D(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ),
    .Q(\BLOCK[3].RAM32.Do0[15] ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[0]  (.DIODE(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[1]  (.DIODE(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[2]  (.DIODE(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[3]  (.DIODE(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[4]  (.DIODE(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[5]  (.DIODE(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[6]  (.DIODE(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[2].DIODE[7]  (.DIODE(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[0]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ),
    .Q(\BLOCK[3].RAM32.Do0[16] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[1]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ),
    .Q(\BLOCK[3].RAM32.Do0[17] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[2]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ),
    .Q(\BLOCK[3].RAM32.Do0[18] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[3]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ),
    .Q(\BLOCK[3].RAM32.Do0[19] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[4]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ),
    .Q(\BLOCK[3].RAM32.Do0[20] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[5]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ),
    .Q(\BLOCK[3].RAM32.Do0[21] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[6]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ),
    .Q(\BLOCK[3].RAM32.Do0[22] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[2].Do_FF[7]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[2] ),
    .D(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ),
    .Q(\BLOCK[3].RAM32.Do0[23] ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[0]  (.DIODE(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[1]  (.DIODE(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[2]  (.DIODE(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[3]  (.DIODE(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[4]  (.DIODE(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[5]  (.DIODE(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[6]  (.DIODE(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[3].DIODE[7]  (.DIODE(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[0]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ),
    .Q(\BLOCK[3].RAM32.Do0[24] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[1]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ),
    .Q(\BLOCK[3].RAM32.Do0[25] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[2]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ),
    .Q(\BLOCK[3].RAM32.Do0[26] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[3]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ),
    .Q(\BLOCK[3].RAM32.Do0[27] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[4]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ),
    .Q(\BLOCK[3].RAM32.Do0[28] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[5]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ),
    .Q(\BLOCK[3].RAM32.Do0[29] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[6]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ),
    .Q(\BLOCK[3].RAM32.Do0[30] ));
 sky130_fd_sc_hd__dfxtp_1 \BLOCK[3].RAM32.Do0_REG.OUTREG_BYTE[3].Do_FF[7]  (.CLK(\BLOCK[3].RAM32.Do0_REG.CLKBUF[3] ),
    .D(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ),
    .Q(\BLOCK[3].RAM32.Do0[31] ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.Do0_REG.Root_CLKBUF  (.A(\BLOCK[3].RAM32.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.Do0_REG.CLK_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.EN0BUF.__cell__  (.A(\BLOCK[3].RAM32.EN0 ),
    .X(\BLOCK[3].RAM32.DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.FBUFENBUF0[0].__cell__  (.A(\BLOCK[3].RAM32.EN0 ),
    .X(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.FBUFENBUF0[1].__cell__  (.A(\BLOCK[3].RAM32.EN0 ),
    .X(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.FBUFENBUF0[2].__cell__  (.A(\BLOCK[3].RAM32.EN0 ),
    .X(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.FBUFENBUF0[3].__cell__  (.A(\BLOCK[3].RAM32.EN0 ),
    .X(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].TE_B ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[0].RAM8.CLKBUF.__cell__  (.A(\BLOCK[3].RAM32.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.ABUF[0]  (.A(\BLOCK[3].RAM32.A0BUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.ABUF[1]  (.A(\BLOCK[3].RAM32.A0BUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.ABUF[2]  (.A(\BLOCK[3].RAM32.A0BUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.AND0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D_N(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.AND1  (.A_N(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.AND2  (.A_N(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .D(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.AND3  (.A_N(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.AND4  (.A_N(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B_N(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.AND5  (.A_N(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.AND6  (.A_N(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.AND7  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.ENBUF  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.EN ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[0].__cell__  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[0].A ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[1].__cell__  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[1].A ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[2].__cell__  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[2].A ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[3].__cell__  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[3].A ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[1].RAM8.CLKBUF.__cell__  (.A(\BLOCK[3].RAM32.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.ABUF[0]  (.A(\BLOCK[3].RAM32.A0BUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.ABUF[1]  (.A(\BLOCK[3].RAM32.A0BUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.ABUF[2]  (.A(\BLOCK[3].RAM32.A0BUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.AND0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D_N(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.AND1  (.A_N(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.AND2  (.A_N(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .D(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.AND3  (.A_N(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.AND4  (.A_N(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B_N(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.AND5  (.A_N(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.AND6  (.A_N(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.AND7  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.ENBUF  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.EN ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[0].__cell__  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[0].A ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[1].__cell__  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[1].A ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[2].__cell__  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[2].A ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[3].__cell__  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[3].A ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[1].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[1].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[2].RAM8.CLKBUF.__cell__  (.A(\BLOCK[3].RAM32.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.ABUF[0]  (.A(\BLOCK[3].RAM32.A0BUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.ABUF[1]  (.A(\BLOCK[3].RAM32.A0BUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.ABUF[2]  (.A(\BLOCK[3].RAM32.A0BUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.AND0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D_N(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.AND1  (.A_N(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.AND2  (.A_N(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .D(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.AND3  (.A_N(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.AND4  (.A_N(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .B_N(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.AND5  (.A_N(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.AND6  (.A_N(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.AND7  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.ENBUF  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.EN ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[0].__cell__  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[0].A ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[1].__cell__  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[1].A ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[2].__cell__  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[2].A ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[3].__cell__  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[3].A ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[2].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[2].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[3].RAM8.CLKBUF.__cell__  (.A(\BLOCK[3].RAM32.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.CLKBUF.X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.ABUF[0]  (.A(\BLOCK[3].RAM32.A0BUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.ABUF[1]  (.A(\BLOCK[3].RAM32.A0BUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.ABUF[2]  (.A(\BLOCK[3].RAM32.A0BUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ));
 sky130_fd_sc_hd__nor4b_2 \BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.AND0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D_N(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.AND1  (.A_N(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.AND2  (.A_N(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .B_N(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .D(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.AND3  (.A_N(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .D(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.SEL0 ));
 sky130_fd_sc_hd__and4bb_2 \BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.AND4  (.A_N(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .B_N(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.AND5  (.A_N(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .C(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.SEL0 ));
 sky130_fd_sc_hd__and4b_2 \BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.AND6  (.A_N(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.SEL0 ));
 sky130_fd_sc_hd__and4_2 \BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.AND7  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[0] ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[1] ),
    .C(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.A_buf[2] ),
    .D(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.EN_buf ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.SEL0 ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.ENBUF  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.EN ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.DEC0.EN_buf ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[0].__cell__  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[0].A ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[0].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[1].__cell__  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[1].A ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[1].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[2].__cell__  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[2].A ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[2].X ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[3].__cell__  (.A(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[3].A ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[3].X ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[0].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[1].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[2].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[3].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[4].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[5].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[6].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[0].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[1].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[1].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[2].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[2].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[3].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[3].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[4].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[4].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[5].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[5].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[6].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[6].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[7].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[7].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[0].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[8].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[8].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[9].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[9].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[10].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[11].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[11].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[12].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[12].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[13].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[13].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[14].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[14].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[15].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[15].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[1].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[1].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[16].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[17].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[17].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[18].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[18].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[19].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[19].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[20].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[20].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[21].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[21].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[22].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[22].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[23].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[23].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[2].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[2].B.CLK_B ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[0].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[0].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[24].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[0] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[1].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[25].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[1].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[25].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[1] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[2].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[26].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[2].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[26].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[2] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[3].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[27].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[3].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[27].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[3] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[4].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[28].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[4].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[28].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[4] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[5].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[29].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[5].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[29].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[5] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[6].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[30].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[6].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[30].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[6] ));
 sky130_fd_sc_hd__ebufn_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[7].OBUF0  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ),
    .TE_B(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ),
    .Z(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[31].Z ));
 sky130_fd_sc_hd__dlxtp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.BIT[7].genblk1.STORAGE  (.D(\BLOCK[3].RAM32.DIBUF[31].X ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ),
    .Q(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.Q_WIRE[7] ));
 sky130_fd_sc_hd__and2_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CGAND  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .B(\BLOCK[3].RAM32.SLICE[3].RAM8.WEBUF[3].X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ));
 sky130_fd_sc_hd__diode_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.DIODE_CLK  (.DIODE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0INV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.SEL0_B ));
 sky130_fd_sc_hd__dlclkp_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.genblk1.CG  (.CLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CLK_B ),
    .GATE(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.WE0_WIRE ),
    .GCLK(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.GCLK ));
 sky130_fd_sc_hd__inv_1 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.genblk1.CLKINV  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ),
    .Y(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[3].B.CLK_B ));
 sky130_fd_sc_hd__clkbuf_4 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.CLKBUF  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.CLKBUF.X ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.CLK ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.SEL0BUF  (.A(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.SEL0 ),
    .X(\BLOCK[3].RAM32.SLICE[3].RAM8.WORD[7].W.BYTE[0].B.SEL0 ));
 sky130_fd_sc_hd__conb_1 \BLOCK[3].RAM32.TIE0[0].__cell__  (.LO(\BLOCK[3].RAM32.BYTE[0].FLOATBUF0[0].A ));
 sky130_fd_sc_hd__conb_1 \BLOCK[3].RAM32.TIE0[1].__cell__  (.LO(\BLOCK[3].RAM32.BYTE[1].FLOATBUF0[10].A ));
 sky130_fd_sc_hd__conb_1 \BLOCK[3].RAM32.TIE0[2].__cell__  (.LO(\BLOCK[3].RAM32.BYTE[2].FLOATBUF0[16].A ));
 sky130_fd_sc_hd__conb_1 \BLOCK[3].RAM32.TIE0[3].__cell__  (.LO(\BLOCK[3].RAM32.BYTE[3].FLOATBUF0[24].A ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.WEBUF[0].__cell__  (.A(\BLOCK[0].RAM32.WEBUF[0].A ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.WEBUF[1].__cell__  (.A(\BLOCK[0].RAM32.WEBUF[1].A ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[1].A ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.WEBUF[2].__cell__  (.A(\BLOCK[0].RAM32.WEBUF[2].A ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[2].A ));
 sky130_fd_sc_hd__clkbuf_2 \BLOCK[3].RAM32.WEBUF[3].__cell__  (.A(\BLOCK[0].RAM32.WEBUF[3].A ),
    .X(\BLOCK[3].RAM32.SLICE[0].RAM8.WEBUF[3].A ));
 sky130_fd_sc_hd__clkbuf_4 \CLKBUF.__cell__  (.A(CLK),
    .X(\BLOCK[0].RAM32.CLK ));
 sky130_fd_sc_hd__nor3b_2 \DEC0.AND0  (.A(\A0BUF[5].X ),
    .B(\A0BUF[6].X ),
    .C_N(\DEC0.EN ),
    .Y(\BLOCK[0].RAM32.EN0 ));
 sky130_fd_sc_hd__and3b_2 \DEC0.AND1  (.A_N(\A0BUF[6].X ),
    .B(\A0BUF[5].X ),
    .C(\DEC0.EN ),
    .X(\BLOCK[1].RAM32.EN0 ));
 sky130_fd_sc_hd__and3b_2 \DEC0.AND2  (.A_N(\A0BUF[5].X ),
    .B(\A0BUF[6].X ),
    .C(\DEC0.EN ),
    .X(\BLOCK[2].RAM32.EN0 ));
 sky130_fd_sc_hd__and3_2 \DEC0.AND3  (.A(\A0BUF[6].X ),
    .B(\A0BUF[5].X ),
    .C(\DEC0.EN ),
    .X(\BLOCK[3].RAM32.EN0 ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[0].__cell__  (.A(Di0[0]),
    .X(\BLOCK[0].RAM32.DIBUF[0].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[10].__cell__  (.A(Di0[10]),
    .X(\BLOCK[0].RAM32.DIBUF[10].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[11].__cell__  (.A(Di0[11]),
    .X(\BLOCK[0].RAM32.DIBUF[11].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[12].__cell__  (.A(Di0[12]),
    .X(\BLOCK[0].RAM32.DIBUF[12].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[13].__cell__  (.A(Di0[13]),
    .X(\BLOCK[0].RAM32.DIBUF[13].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[14].__cell__  (.A(Di0[14]),
    .X(\BLOCK[0].RAM32.DIBUF[14].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[15].__cell__  (.A(Di0[15]),
    .X(\BLOCK[0].RAM32.DIBUF[15].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[16].__cell__  (.A(Di0[16]),
    .X(\BLOCK[0].RAM32.DIBUF[16].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[17].__cell__  (.A(Di0[17]),
    .X(\BLOCK[0].RAM32.DIBUF[17].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[18].__cell__  (.A(Di0[18]),
    .X(\BLOCK[0].RAM32.DIBUF[18].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[19].__cell__  (.A(Di0[19]),
    .X(\BLOCK[0].RAM32.DIBUF[19].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[1].__cell__  (.A(Di0[1]),
    .X(\BLOCK[0].RAM32.DIBUF[1].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[20].__cell__  (.A(Di0[20]),
    .X(\BLOCK[0].RAM32.DIBUF[20].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[21].__cell__  (.A(Di0[21]),
    .X(\BLOCK[0].RAM32.DIBUF[21].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[22].__cell__  (.A(Di0[22]),
    .X(\BLOCK[0].RAM32.DIBUF[22].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[23].__cell__  (.A(Di0[23]),
    .X(\BLOCK[0].RAM32.DIBUF[23].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[24].__cell__  (.A(Di0[24]),
    .X(\BLOCK[0].RAM32.DIBUF[24].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[25].__cell__  (.A(Di0[25]),
    .X(\BLOCK[0].RAM32.DIBUF[25].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[26].__cell__  (.A(Di0[26]),
    .X(\BLOCK[0].RAM32.DIBUF[26].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[27].__cell__  (.A(Di0[27]),
    .X(\BLOCK[0].RAM32.DIBUF[27].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[28].__cell__  (.A(Di0[28]),
    .X(\BLOCK[0].RAM32.DIBUF[28].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[29].__cell__  (.A(Di0[29]),
    .X(\BLOCK[0].RAM32.DIBUF[29].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[2].__cell__  (.A(Di0[2]),
    .X(\BLOCK[0].RAM32.DIBUF[2].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[30].__cell__  (.A(Di0[30]),
    .X(\BLOCK[0].RAM32.DIBUF[30].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[31].__cell__  (.A(Di0[31]),
    .X(\BLOCK[0].RAM32.DIBUF[31].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[3].__cell__  (.A(Di0[3]),
    .X(\BLOCK[0].RAM32.DIBUF[3].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[4].__cell__  (.A(Di0[4]),
    .X(\BLOCK[0].RAM32.DIBUF[4].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[5].__cell__  (.A(Di0[5]),
    .X(\BLOCK[0].RAM32.DIBUF[5].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[6].__cell__  (.A(Di0[6]),
    .X(\BLOCK[0].RAM32.DIBUF[6].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[7].__cell__  (.A(Di0[7]),
    .X(\BLOCK[0].RAM32.DIBUF[7].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[8].__cell__  (.A(Di0[8]),
    .X(\BLOCK[0].RAM32.DIBUF[8].A ));
 sky130_fd_sc_hd__clkbuf_16 \DIBUF[9].__cell__  (.A(Di0[9]),
    .X(\BLOCK[0].RAM32.DIBUF[9].A ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[0]  (.DIODE(\BLOCK[0].RAM32.Do0[0] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[1]  (.DIODE(\BLOCK[0].RAM32.Do0[1] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[2]  (.DIODE(\BLOCK[0].RAM32.Do0[2] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[3]  (.DIODE(\BLOCK[0].RAM32.Do0[3] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[4]  (.DIODE(\BLOCK[0].RAM32.Do0[4] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[5]  (.DIODE(\BLOCK[0].RAM32.Do0[5] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[6]  (.DIODE(\BLOCK[0].RAM32.Do0[6] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A0MUX[7]  (.DIODE(\BLOCK[0].RAM32.Do0[7] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[0]  (.DIODE(\BLOCK[1].RAM32.Do0[0] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[1]  (.DIODE(\BLOCK[1].RAM32.Do0[1] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[2]  (.DIODE(\BLOCK[1].RAM32.Do0[2] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[3]  (.DIODE(\BLOCK[1].RAM32.Do0[3] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[4]  (.DIODE(\BLOCK[1].RAM32.Do0[4] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[5]  (.DIODE(\BLOCK[1].RAM32.Do0[5] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[6]  (.DIODE(\BLOCK[1].RAM32.Do0[6] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A1MUX[7]  (.DIODE(\BLOCK[1].RAM32.Do0[7] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A2MUX[0]  (.DIODE(\BLOCK[2].RAM32.Do0[0] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A2MUX[1]  (.DIODE(\BLOCK[2].RAM32.Do0[1] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A2MUX[2]  (.DIODE(\BLOCK[2].RAM32.Do0[2] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A2MUX[3]  (.DIODE(\BLOCK[2].RAM32.Do0[3] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A2MUX[4]  (.DIODE(\BLOCK[2].RAM32.Do0[4] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A2MUX[5]  (.DIODE(\BLOCK[2].RAM32.Do0[5] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A2MUX[6]  (.DIODE(\BLOCK[2].RAM32.Do0[6] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A2MUX[7]  (.DIODE(\BLOCK[2].RAM32.Do0[7] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A3MUX[0]  (.DIODE(\BLOCK[3].RAM32.Do0[0] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A3MUX[1]  (.DIODE(\BLOCK[3].RAM32.Do0[1] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A3MUX[2]  (.DIODE(\BLOCK[3].RAM32.Do0[2] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A3MUX[3]  (.DIODE(\BLOCK[3].RAM32.Do0[3] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A3MUX[4]  (.DIODE(\BLOCK[3].RAM32.Do0[4] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A3MUX[5]  (.DIODE(\BLOCK[3].RAM32.Do0[5] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A3MUX[6]  (.DIODE(\BLOCK[3].RAM32.Do0[6] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[0].DIODE_A3MUX[7]  (.DIODE(\BLOCK[3].RAM32.Do0[7] ));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[0].MUX[0]  (.A0(\BLOCK[0].RAM32.Do0[0] ),
    .A1(\BLOCK[1].RAM32.Do0[0] ),
    .A2(\BLOCK[2].RAM32.Do0[0] ),
    .A3(\BLOCK[3].RAM32.Do0[0] ),
    .S0(\Do0MUX.SEL0[0] ),
    .S1(\Do0MUX.SEL1[0] ),
    .X(Do0[0]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[0].MUX[1]  (.A0(\BLOCK[0].RAM32.Do0[1] ),
    .A1(\BLOCK[1].RAM32.Do0[1] ),
    .A2(\BLOCK[2].RAM32.Do0[1] ),
    .A3(\BLOCK[3].RAM32.Do0[1] ),
    .S0(\Do0MUX.SEL0[0] ),
    .S1(\Do0MUX.SEL1[0] ),
    .X(Do0[1]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[0].MUX[2]  (.A0(\BLOCK[0].RAM32.Do0[2] ),
    .A1(\BLOCK[1].RAM32.Do0[2] ),
    .A2(\BLOCK[2].RAM32.Do0[2] ),
    .A3(\BLOCK[3].RAM32.Do0[2] ),
    .S0(\Do0MUX.SEL0[0] ),
    .S1(\Do0MUX.SEL1[0] ),
    .X(Do0[2]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[0].MUX[3]  (.A0(\BLOCK[0].RAM32.Do0[3] ),
    .A1(\BLOCK[1].RAM32.Do0[3] ),
    .A2(\BLOCK[2].RAM32.Do0[3] ),
    .A3(\BLOCK[3].RAM32.Do0[3] ),
    .S0(\Do0MUX.SEL0[0] ),
    .S1(\Do0MUX.SEL1[0] ),
    .X(Do0[3]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[0].MUX[4]  (.A0(\BLOCK[0].RAM32.Do0[4] ),
    .A1(\BLOCK[1].RAM32.Do0[4] ),
    .A2(\BLOCK[2].RAM32.Do0[4] ),
    .A3(\BLOCK[3].RAM32.Do0[4] ),
    .S0(\Do0MUX.SEL0[0] ),
    .S1(\Do0MUX.SEL1[0] ),
    .X(Do0[4]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[0].MUX[5]  (.A0(\BLOCK[0].RAM32.Do0[5] ),
    .A1(\BLOCK[1].RAM32.Do0[5] ),
    .A2(\BLOCK[2].RAM32.Do0[5] ),
    .A3(\BLOCK[3].RAM32.Do0[5] ),
    .S0(\Do0MUX.SEL0[0] ),
    .S1(\Do0MUX.SEL1[0] ),
    .X(Do0[5]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[0].MUX[6]  (.A0(\BLOCK[0].RAM32.Do0[6] ),
    .A1(\BLOCK[1].RAM32.Do0[6] ),
    .A2(\BLOCK[2].RAM32.Do0[6] ),
    .A3(\BLOCK[3].RAM32.Do0[6] ),
    .S0(\Do0MUX.SEL0[0] ),
    .S1(\Do0MUX.SEL1[0] ),
    .X(Do0[6]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[0].MUX[7]  (.A0(\BLOCK[0].RAM32.Do0[7] ),
    .A1(\BLOCK[1].RAM32.Do0[7] ),
    .A2(\BLOCK[2].RAM32.Do0[7] ),
    .A3(\BLOCK[3].RAM32.Do0[7] ),
    .S0(\Do0MUX.SEL0[0] ),
    .S1(\Do0MUX.SEL1[0] ),
    .X(Do0[7]));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A0MUX[10]  (.DIODE(\BLOCK[0].RAM32.Do0[10] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A0MUX[11]  (.DIODE(\BLOCK[0].RAM32.Do0[11] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A0MUX[12]  (.DIODE(\BLOCK[0].RAM32.Do0[12] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A0MUX[13]  (.DIODE(\BLOCK[0].RAM32.Do0[13] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A0MUX[14]  (.DIODE(\BLOCK[0].RAM32.Do0[14] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A0MUX[15]  (.DIODE(\BLOCK[0].RAM32.Do0[15] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A0MUX[8]  (.DIODE(\BLOCK[0].RAM32.Do0[8] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A0MUX[9]  (.DIODE(\BLOCK[0].RAM32.Do0[9] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A1MUX[10]  (.DIODE(\BLOCK[1].RAM32.Do0[10] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A1MUX[11]  (.DIODE(\BLOCK[1].RAM32.Do0[11] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A1MUX[12]  (.DIODE(\BLOCK[1].RAM32.Do0[12] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A1MUX[13]  (.DIODE(\BLOCK[1].RAM32.Do0[13] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A1MUX[14]  (.DIODE(\BLOCK[1].RAM32.Do0[14] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A1MUX[15]  (.DIODE(\BLOCK[1].RAM32.Do0[15] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A1MUX[8]  (.DIODE(\BLOCK[1].RAM32.Do0[8] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A1MUX[9]  (.DIODE(\BLOCK[1].RAM32.Do0[9] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A2MUX[10]  (.DIODE(\BLOCK[2].RAM32.Do0[10] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A2MUX[11]  (.DIODE(\BLOCK[2].RAM32.Do0[11] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A2MUX[12]  (.DIODE(\BLOCK[2].RAM32.Do0[12] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A2MUX[13]  (.DIODE(\BLOCK[2].RAM32.Do0[13] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A2MUX[14]  (.DIODE(\BLOCK[2].RAM32.Do0[14] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A2MUX[15]  (.DIODE(\BLOCK[2].RAM32.Do0[15] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A2MUX[8]  (.DIODE(\BLOCK[2].RAM32.Do0[8] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A2MUX[9]  (.DIODE(\BLOCK[2].RAM32.Do0[9] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A3MUX[10]  (.DIODE(\BLOCK[3].RAM32.Do0[10] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A3MUX[11]  (.DIODE(\BLOCK[3].RAM32.Do0[11] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A3MUX[12]  (.DIODE(\BLOCK[3].RAM32.Do0[12] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A3MUX[13]  (.DIODE(\BLOCK[3].RAM32.Do0[13] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A3MUX[14]  (.DIODE(\BLOCK[3].RAM32.Do0[14] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A3MUX[15]  (.DIODE(\BLOCK[3].RAM32.Do0[15] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A3MUX[8]  (.DIODE(\BLOCK[3].RAM32.Do0[8] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[1].DIODE_A3MUX[9]  (.DIODE(\BLOCK[3].RAM32.Do0[9] ));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[1].MUX[0]  (.A0(\BLOCK[0].RAM32.Do0[8] ),
    .A1(\BLOCK[1].RAM32.Do0[8] ),
    .A2(\BLOCK[2].RAM32.Do0[8] ),
    .A3(\BLOCK[3].RAM32.Do0[8] ),
    .S0(\Do0MUX.SEL0[1] ),
    .S1(\Do0MUX.SEL1[1] ),
    .X(Do0[8]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[1].MUX[1]  (.A0(\BLOCK[0].RAM32.Do0[9] ),
    .A1(\BLOCK[1].RAM32.Do0[9] ),
    .A2(\BLOCK[2].RAM32.Do0[9] ),
    .A3(\BLOCK[3].RAM32.Do0[9] ),
    .S0(\Do0MUX.SEL0[1] ),
    .S1(\Do0MUX.SEL1[1] ),
    .X(Do0[9]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[1].MUX[2]  (.A0(\BLOCK[0].RAM32.Do0[10] ),
    .A1(\BLOCK[1].RAM32.Do0[10] ),
    .A2(\BLOCK[2].RAM32.Do0[10] ),
    .A3(\BLOCK[3].RAM32.Do0[10] ),
    .S0(\Do0MUX.SEL0[1] ),
    .S1(\Do0MUX.SEL1[1] ),
    .X(Do0[10]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[1].MUX[3]  (.A0(\BLOCK[0].RAM32.Do0[11] ),
    .A1(\BLOCK[1].RAM32.Do0[11] ),
    .A2(\BLOCK[2].RAM32.Do0[11] ),
    .A3(\BLOCK[3].RAM32.Do0[11] ),
    .S0(\Do0MUX.SEL0[1] ),
    .S1(\Do0MUX.SEL1[1] ),
    .X(Do0[11]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[1].MUX[4]  (.A0(\BLOCK[0].RAM32.Do0[12] ),
    .A1(\BLOCK[1].RAM32.Do0[12] ),
    .A2(\BLOCK[2].RAM32.Do0[12] ),
    .A3(\BLOCK[3].RAM32.Do0[12] ),
    .S0(\Do0MUX.SEL0[1] ),
    .S1(\Do0MUX.SEL1[1] ),
    .X(Do0[12]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[1].MUX[5]  (.A0(\BLOCK[0].RAM32.Do0[13] ),
    .A1(\BLOCK[1].RAM32.Do0[13] ),
    .A2(\BLOCK[2].RAM32.Do0[13] ),
    .A3(\BLOCK[3].RAM32.Do0[13] ),
    .S0(\Do0MUX.SEL0[1] ),
    .S1(\Do0MUX.SEL1[1] ),
    .X(Do0[13]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[1].MUX[6]  (.A0(\BLOCK[0].RAM32.Do0[14] ),
    .A1(\BLOCK[1].RAM32.Do0[14] ),
    .A2(\BLOCK[2].RAM32.Do0[14] ),
    .A3(\BLOCK[3].RAM32.Do0[14] ),
    .S0(\Do0MUX.SEL0[1] ),
    .S1(\Do0MUX.SEL1[1] ),
    .X(Do0[14]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[1].MUX[7]  (.A0(\BLOCK[0].RAM32.Do0[15] ),
    .A1(\BLOCK[1].RAM32.Do0[15] ),
    .A2(\BLOCK[2].RAM32.Do0[15] ),
    .A3(\BLOCK[3].RAM32.Do0[15] ),
    .S0(\Do0MUX.SEL0[1] ),
    .S1(\Do0MUX.SEL1[1] ),
    .X(Do0[15]));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A0MUX[16]  (.DIODE(\BLOCK[0].RAM32.Do0[16] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A0MUX[17]  (.DIODE(\BLOCK[0].RAM32.Do0[17] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A0MUX[18]  (.DIODE(\BLOCK[0].RAM32.Do0[18] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A0MUX[19]  (.DIODE(\BLOCK[0].RAM32.Do0[19] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A0MUX[20]  (.DIODE(\BLOCK[0].RAM32.Do0[20] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A0MUX[21]  (.DIODE(\BLOCK[0].RAM32.Do0[21] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A0MUX[22]  (.DIODE(\BLOCK[0].RAM32.Do0[22] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A0MUX[23]  (.DIODE(\BLOCK[0].RAM32.Do0[23] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A1MUX[16]  (.DIODE(\BLOCK[1].RAM32.Do0[16] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A1MUX[17]  (.DIODE(\BLOCK[1].RAM32.Do0[17] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A1MUX[18]  (.DIODE(\BLOCK[1].RAM32.Do0[18] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A1MUX[19]  (.DIODE(\BLOCK[1].RAM32.Do0[19] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A1MUX[20]  (.DIODE(\BLOCK[1].RAM32.Do0[20] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A1MUX[21]  (.DIODE(\BLOCK[1].RAM32.Do0[21] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A1MUX[22]  (.DIODE(\BLOCK[1].RAM32.Do0[22] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A1MUX[23]  (.DIODE(\BLOCK[1].RAM32.Do0[23] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A2MUX[16]  (.DIODE(\BLOCK[2].RAM32.Do0[16] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A2MUX[17]  (.DIODE(\BLOCK[2].RAM32.Do0[17] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A2MUX[18]  (.DIODE(\BLOCK[2].RAM32.Do0[18] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A2MUX[19]  (.DIODE(\BLOCK[2].RAM32.Do0[19] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A2MUX[20]  (.DIODE(\BLOCK[2].RAM32.Do0[20] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A2MUX[21]  (.DIODE(\BLOCK[2].RAM32.Do0[21] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A2MUX[22]  (.DIODE(\BLOCK[2].RAM32.Do0[22] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A2MUX[23]  (.DIODE(\BLOCK[2].RAM32.Do0[23] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A3MUX[16]  (.DIODE(\BLOCK[3].RAM32.Do0[16] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A3MUX[17]  (.DIODE(\BLOCK[3].RAM32.Do0[17] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A3MUX[18]  (.DIODE(\BLOCK[3].RAM32.Do0[18] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A3MUX[19]  (.DIODE(\BLOCK[3].RAM32.Do0[19] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A3MUX[20]  (.DIODE(\BLOCK[3].RAM32.Do0[20] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A3MUX[21]  (.DIODE(\BLOCK[3].RAM32.Do0[21] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A3MUX[22]  (.DIODE(\BLOCK[3].RAM32.Do0[22] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[2].DIODE_A3MUX[23]  (.DIODE(\BLOCK[3].RAM32.Do0[23] ));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[2].MUX[0]  (.A0(\BLOCK[0].RAM32.Do0[16] ),
    .A1(\BLOCK[1].RAM32.Do0[16] ),
    .A2(\BLOCK[2].RAM32.Do0[16] ),
    .A3(\BLOCK[3].RAM32.Do0[16] ),
    .S0(\Do0MUX.SEL0[2] ),
    .S1(\Do0MUX.SEL1[2] ),
    .X(Do0[16]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[2].MUX[1]  (.A0(\BLOCK[0].RAM32.Do0[17] ),
    .A1(\BLOCK[1].RAM32.Do0[17] ),
    .A2(\BLOCK[2].RAM32.Do0[17] ),
    .A3(\BLOCK[3].RAM32.Do0[17] ),
    .S0(\Do0MUX.SEL0[2] ),
    .S1(\Do0MUX.SEL1[2] ),
    .X(Do0[17]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[2].MUX[2]  (.A0(\BLOCK[0].RAM32.Do0[18] ),
    .A1(\BLOCK[1].RAM32.Do0[18] ),
    .A2(\BLOCK[2].RAM32.Do0[18] ),
    .A3(\BLOCK[3].RAM32.Do0[18] ),
    .S0(\Do0MUX.SEL0[2] ),
    .S1(\Do0MUX.SEL1[2] ),
    .X(Do0[18]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[2].MUX[3]  (.A0(\BLOCK[0].RAM32.Do0[19] ),
    .A1(\BLOCK[1].RAM32.Do0[19] ),
    .A2(\BLOCK[2].RAM32.Do0[19] ),
    .A3(\BLOCK[3].RAM32.Do0[19] ),
    .S0(\Do0MUX.SEL0[2] ),
    .S1(\Do0MUX.SEL1[2] ),
    .X(Do0[19]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[2].MUX[4]  (.A0(\BLOCK[0].RAM32.Do0[20] ),
    .A1(\BLOCK[1].RAM32.Do0[20] ),
    .A2(\BLOCK[2].RAM32.Do0[20] ),
    .A3(\BLOCK[3].RAM32.Do0[20] ),
    .S0(\Do0MUX.SEL0[2] ),
    .S1(\Do0MUX.SEL1[2] ),
    .X(Do0[20]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[2].MUX[5]  (.A0(\BLOCK[0].RAM32.Do0[21] ),
    .A1(\BLOCK[1].RAM32.Do0[21] ),
    .A2(\BLOCK[2].RAM32.Do0[21] ),
    .A3(\BLOCK[3].RAM32.Do0[21] ),
    .S0(\Do0MUX.SEL0[2] ),
    .S1(\Do0MUX.SEL1[2] ),
    .X(Do0[21]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[2].MUX[6]  (.A0(\BLOCK[0].RAM32.Do0[22] ),
    .A1(\BLOCK[1].RAM32.Do0[22] ),
    .A2(\BLOCK[2].RAM32.Do0[22] ),
    .A3(\BLOCK[3].RAM32.Do0[22] ),
    .S0(\Do0MUX.SEL0[2] ),
    .S1(\Do0MUX.SEL1[2] ),
    .X(Do0[22]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[2].MUX[7]  (.A0(\BLOCK[0].RAM32.Do0[23] ),
    .A1(\BLOCK[1].RAM32.Do0[23] ),
    .A2(\BLOCK[2].RAM32.Do0[23] ),
    .A3(\BLOCK[3].RAM32.Do0[23] ),
    .S0(\Do0MUX.SEL0[2] ),
    .S1(\Do0MUX.SEL1[2] ),
    .X(Do0[23]));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A0MUX[24]  (.DIODE(\BLOCK[0].RAM32.Do0[24] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A0MUX[25]  (.DIODE(\BLOCK[0].RAM32.Do0[25] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A0MUX[26]  (.DIODE(\BLOCK[0].RAM32.Do0[26] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A0MUX[27]  (.DIODE(\BLOCK[0].RAM32.Do0[27] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A0MUX[28]  (.DIODE(\BLOCK[0].RAM32.Do0[28] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A0MUX[29]  (.DIODE(\BLOCK[0].RAM32.Do0[29] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A0MUX[30]  (.DIODE(\BLOCK[0].RAM32.Do0[30] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A0MUX[31]  (.DIODE(\BLOCK[0].RAM32.Do0[31] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A1MUX[24]  (.DIODE(\BLOCK[1].RAM32.Do0[24] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A1MUX[25]  (.DIODE(\BLOCK[1].RAM32.Do0[25] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A1MUX[26]  (.DIODE(\BLOCK[1].RAM32.Do0[26] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A1MUX[27]  (.DIODE(\BLOCK[1].RAM32.Do0[27] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A1MUX[28]  (.DIODE(\BLOCK[1].RAM32.Do0[28] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A1MUX[29]  (.DIODE(\BLOCK[1].RAM32.Do0[29] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A1MUX[30]  (.DIODE(\BLOCK[1].RAM32.Do0[30] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A1MUX[31]  (.DIODE(\BLOCK[1].RAM32.Do0[31] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A2MUX[24]  (.DIODE(\BLOCK[2].RAM32.Do0[24] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A2MUX[25]  (.DIODE(\BLOCK[2].RAM32.Do0[25] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A2MUX[26]  (.DIODE(\BLOCK[2].RAM32.Do0[26] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A2MUX[27]  (.DIODE(\BLOCK[2].RAM32.Do0[27] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A2MUX[28]  (.DIODE(\BLOCK[2].RAM32.Do0[28] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A2MUX[29]  (.DIODE(\BLOCK[2].RAM32.Do0[29] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A2MUX[30]  (.DIODE(\BLOCK[2].RAM32.Do0[30] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A2MUX[31]  (.DIODE(\BLOCK[2].RAM32.Do0[31] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A3MUX[24]  (.DIODE(\BLOCK[3].RAM32.Do0[24] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A3MUX[25]  (.DIODE(\BLOCK[3].RAM32.Do0[25] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A3MUX[26]  (.DIODE(\BLOCK[3].RAM32.Do0[26] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A3MUX[27]  (.DIODE(\BLOCK[3].RAM32.Do0[27] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A3MUX[28]  (.DIODE(\BLOCK[3].RAM32.Do0[28] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A3MUX[29]  (.DIODE(\BLOCK[3].RAM32.Do0[29] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A3MUX[30]  (.DIODE(\BLOCK[3].RAM32.Do0[30] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.M[3].DIODE_A3MUX[31]  (.DIODE(\BLOCK[3].RAM32.Do0[31] ));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[3].MUX[0]  (.A0(\BLOCK[0].RAM32.Do0[24] ),
    .A1(\BLOCK[1].RAM32.Do0[24] ),
    .A2(\BLOCK[2].RAM32.Do0[24] ),
    .A3(\BLOCK[3].RAM32.Do0[24] ),
    .S0(\Do0MUX.SEL0[3] ),
    .S1(\Do0MUX.SEL1[3] ),
    .X(Do0[24]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[3].MUX[1]  (.A0(\BLOCK[0].RAM32.Do0[25] ),
    .A1(\BLOCK[1].RAM32.Do0[25] ),
    .A2(\BLOCK[2].RAM32.Do0[25] ),
    .A3(\BLOCK[3].RAM32.Do0[25] ),
    .S0(\Do0MUX.SEL0[3] ),
    .S1(\Do0MUX.SEL1[3] ),
    .X(Do0[25]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[3].MUX[2]  (.A0(\BLOCK[0].RAM32.Do0[26] ),
    .A1(\BLOCK[1].RAM32.Do0[26] ),
    .A2(\BLOCK[2].RAM32.Do0[26] ),
    .A3(\BLOCK[3].RAM32.Do0[26] ),
    .S0(\Do0MUX.SEL0[3] ),
    .S1(\Do0MUX.SEL1[3] ),
    .X(Do0[26]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[3].MUX[3]  (.A0(\BLOCK[0].RAM32.Do0[27] ),
    .A1(\BLOCK[1].RAM32.Do0[27] ),
    .A2(\BLOCK[2].RAM32.Do0[27] ),
    .A3(\BLOCK[3].RAM32.Do0[27] ),
    .S0(\Do0MUX.SEL0[3] ),
    .S1(\Do0MUX.SEL1[3] ),
    .X(Do0[27]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[3].MUX[4]  (.A0(\BLOCK[0].RAM32.Do0[28] ),
    .A1(\BLOCK[1].RAM32.Do0[28] ),
    .A2(\BLOCK[2].RAM32.Do0[28] ),
    .A3(\BLOCK[3].RAM32.Do0[28] ),
    .S0(\Do0MUX.SEL0[3] ),
    .S1(\Do0MUX.SEL1[3] ),
    .X(Do0[28]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[3].MUX[5]  (.A0(\BLOCK[0].RAM32.Do0[29] ),
    .A1(\BLOCK[1].RAM32.Do0[29] ),
    .A2(\BLOCK[2].RAM32.Do0[29] ),
    .A3(\BLOCK[3].RAM32.Do0[29] ),
    .S0(\Do0MUX.SEL0[3] ),
    .S1(\Do0MUX.SEL1[3] ),
    .X(Do0[29]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[3].MUX[6]  (.A0(\BLOCK[0].RAM32.Do0[30] ),
    .A1(\BLOCK[1].RAM32.Do0[30] ),
    .A2(\BLOCK[2].RAM32.Do0[30] ),
    .A3(\BLOCK[3].RAM32.Do0[30] ),
    .S0(\Do0MUX.SEL0[3] ),
    .S1(\Do0MUX.SEL1[3] ),
    .X(Do0[30]));
 sky130_fd_sc_hd__mux4_1 \Do0MUX.M[3].MUX[7]  (.A0(\BLOCK[0].RAM32.Do0[31] ),
    .A1(\BLOCK[1].RAM32.Do0[31] ),
    .A2(\BLOCK[2].RAM32.Do0[31] ),
    .A3(\BLOCK[3].RAM32.Do0[31] ),
    .S0(\Do0MUX.SEL0[3] ),
    .S1(\Do0MUX.SEL1[3] ),
    .X(Do0[31]));
 sky130_fd_sc_hd__clkbuf_2 \Do0MUX.SEL0BUF[0]  (.A(\A0BUF[5].X ),
    .X(\Do0MUX.SEL0[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Do0MUX.SEL0BUF[1]  (.A(\A0BUF[5].X ),
    .X(\Do0MUX.SEL0[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Do0MUX.SEL0BUF[2]  (.A(\A0BUF[5].X ),
    .X(\Do0MUX.SEL0[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Do0MUX.SEL0BUF[3]  (.A(\A0BUF[5].X ),
    .X(\Do0MUX.SEL0[3] ));
 sky130_fd_sc_hd__clkbuf_2 \Do0MUX.SEL1BUF[0]  (.A(\A0BUF[6].X ),
    .X(\Do0MUX.SEL1[0] ));
 sky130_fd_sc_hd__clkbuf_2 \Do0MUX.SEL1BUF[1]  (.A(\A0BUF[6].X ),
    .X(\Do0MUX.SEL1[1] ));
 sky130_fd_sc_hd__clkbuf_2 \Do0MUX.SEL1BUF[2]  (.A(\A0BUF[6].X ),
    .X(\Do0MUX.SEL1[2] ));
 sky130_fd_sc_hd__clkbuf_2 \Do0MUX.SEL1BUF[3]  (.A(\A0BUF[6].X ),
    .X(\Do0MUX.SEL1[3] ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.SEL_DIODE[0]  (.DIODE(\A0BUF[5].X ));
 sky130_fd_sc_hd__diode_2 \Do0MUX.SEL_DIODE[1]  (.DIODE(\A0BUF[6].X ));
 sky130_fd_sc_hd__clkbuf_2 \EN0BUF.__cell__  (.A(EN0),
    .X(\DEC0.EN ));
 sky130_fd_sc_hd__clkbuf_2 \WEBUF[0].__cell__  (.A(WE0[0]),
    .X(\BLOCK[0].RAM32.WEBUF[0].A ));
 sky130_fd_sc_hd__clkbuf_2 \WEBUF[1].__cell__  (.A(WE0[1]),
    .X(\BLOCK[0].RAM32.WEBUF[1].A ));
 sky130_fd_sc_hd__clkbuf_2 \WEBUF[2].__cell__  (.A(WE0[2]),
    .X(\BLOCK[0].RAM32.WEBUF[2].A ));
 sky130_fd_sc_hd__clkbuf_2 \WEBUF[3].__cell__  (.A(WE0[3]),
    .X(\BLOCK[0].RAM32.WEBUF[3].A ));
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_0_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_1_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_2_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_4_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_6_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_7_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_8_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_9_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_2_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_4_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_6_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_7_0 ();
 sky130_fd_sc_hd__decap_3 fill_7_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_1 ();
 sky130_fd_sc_hd__decap_3 fill_8_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_9_0 ();
 sky130_fd_sc_hd__decap_3 fill_9_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_12_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_14_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_15_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_16_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_17_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_10_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_12_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_15_0 ();
 sky130_fd_sc_hd__decap_3 fill_15_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_1 ();
 sky130_fd_sc_hd__decap_3 fill_16_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_0 ();
 sky130_fd_sc_hd__decap_3 fill_17_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_18_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_19_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_20_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_21_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_22_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_23_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_24_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_25_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_20_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_22_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_23_0 ();
 sky130_fd_sc_hd__decap_3 fill_23_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_1 ();
 sky130_fd_sc_hd__decap_3 fill_24_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_25_0 ();
 sky130_fd_sc_hd__decap_3 fill_25_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_26_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_27_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_28_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_29_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_30_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_31_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_32_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_33_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_26_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_28_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_30_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_31_0 ();
 sky130_fd_sc_hd__decap_3 fill_31_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_1 ();
 sky130_fd_sc_hd__decap_3 fill_32_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_0 ();
 sky130_fd_sc_hd__decap_3 fill_33_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_34_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_35_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_36_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_38_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_39_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_40_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_41_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_42_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_43_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_44_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_40_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_42_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_44_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_42_1 ();
 sky130_fd_sc_hd__decap_3 fill_42_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_43_0 ();
 sky130_fd_sc_hd__decap_3 fill_43_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_44_1 ();
 sky130_fd_sc_hd__decap_3 fill_44_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_46_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_47_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_48_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_49_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_50_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_51_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_52_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_46_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_48_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_50_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_52_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_50_1 ();
 sky130_fd_sc_hd__decap_3 fill_50_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_51_0 ();
 sky130_fd_sc_hd__decap_3 fill_51_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_52_1 ();
 sky130_fd_sc_hd__decap_3 fill_52_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_54_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_55_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_56_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_57_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_58_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_59_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_60_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_54_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_56_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_58_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_60_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_58_1 ();
 sky130_fd_sc_hd__decap_3 fill_58_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_59_0 ();
 sky130_fd_sc_hd__decap_3 fill_59_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_60_1 ();
 sky130_fd_sc_hd__decap_3 fill_60_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_61_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_62_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_63_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_64_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_65_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_66_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_67_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_68_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_62_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_64_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_66_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_68_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_66_1 ();
 sky130_fd_sc_hd__decap_3 fill_66_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_67_0 ();
 sky130_fd_sc_hd__decap_3 fill_67_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_68_1 ();
 sky130_fd_sc_hd__decap_3 fill_68_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_69_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_69_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_69_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_69_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_69_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_69_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_69_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_69_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_69_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_69_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_69_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_70_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_37_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_45_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_53_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_71_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_72_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_73_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_74_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_75_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_76_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_77_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_78_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_79_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_72_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_74_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_76_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_78_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_77_0 ();
 sky130_fd_sc_hd__decap_3 fill_77_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_78_1 ();
 sky130_fd_sc_hd__decap_3 fill_78_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_79_0 ();
 sky130_fd_sc_hd__decap_3 fill_79_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_80_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_81_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_82_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_83_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_84_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_85_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_86_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_87_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_80_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_82_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_84_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_86_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_85_0 ();
 sky130_fd_sc_hd__decap_3 fill_85_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_86_1 ();
 sky130_fd_sc_hd__decap_3 fill_86_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_87_0 ();
 sky130_fd_sc_hd__decap_3 fill_87_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_88_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_89_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_90_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_91_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_92_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_93_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_94_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_95_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_88_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_90_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_92_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_94_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_93_0 ();
 sky130_fd_sc_hd__decap_3 fill_93_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_94_1 ();
 sky130_fd_sc_hd__decap_3 fill_94_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_95_0 ();
 sky130_fd_sc_hd__decap_3 fill_95_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_96_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_97_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_98_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_99_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_100_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_101_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_102_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_103_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_96_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_98_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_100_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_102_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_101_0 ();
 sky130_fd_sc_hd__decap_3 fill_101_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_102_1 ();
 sky130_fd_sc_hd__decap_3 fill_102_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_103_0 ();
 sky130_fd_sc_hd__decap_3 fill_103_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_104_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_104_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_104_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_104_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_104_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_104_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_104_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_104_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_104_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_104_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_105_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_106_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_108_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_109_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_110_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_111_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_112_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_113_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_114_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_108_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_110_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_112_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_114_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_112_1 ();
 sky130_fd_sc_hd__decap_3 fill_112_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_113_0 ();
 sky130_fd_sc_hd__decap_3 fill_113_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_114_1 ();
 sky130_fd_sc_hd__decap_3 fill_114_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_116_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_117_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_118_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_119_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_120_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_121_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_122_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_116_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_118_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_120_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_122_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_120_1 ();
 sky130_fd_sc_hd__decap_3 fill_120_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_121_0 ();
 sky130_fd_sc_hd__decap_3 fill_121_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_122_1 ();
 sky130_fd_sc_hd__decap_3 fill_122_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_124_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_125_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_126_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_127_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_128_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_129_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_130_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_124_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_126_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_128_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_130_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_128_1 ();
 sky130_fd_sc_hd__decap_3 fill_128_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_129_0 ();
 sky130_fd_sc_hd__decap_3 fill_129_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_130_1 ();
 sky130_fd_sc_hd__decap_3 fill_130_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_131_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_132_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_133_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_134_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_135_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_136_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_137_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_138_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_132_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_134_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_136_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_138_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_136_1 ();
 sky130_fd_sc_hd__decap_3 fill_136_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_137_0 ();
 sky130_fd_sc_hd__decap_3 fill_137_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_138_1 ();
 sky130_fd_sc_hd__decap_3 fill_138_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_139_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_139_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_139_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_139_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_139_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_139_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_139_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_139_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_139_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_139_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_139_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_140_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_107_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_115_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_123_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_7 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_10 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_12 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_13 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_15 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_16 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_18 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_19 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_24 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_25 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_141_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_142_0 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_142_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_142_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_142_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_142_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_142_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_142_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_3_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_5_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_10_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_11_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 tap_13_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_0 ();
 sky130_fd_sc_hd__decap_12 fill_0_1 ();
 sky130_fd_sc_hd__decap_12 fill_0_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_3 ();
 sky130_fd_sc_hd__decap_12 fill_0_4 ();
 sky130_fd_sc_hd__decap_12 fill_0_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_6 ();
 sky130_fd_sc_hd__decap_12 fill_0_7 ();
 sky130_fd_sc_hd__decap_12 fill_0_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_9 ();
 sky130_fd_sc_hd__decap_12 fill_0_10 ();
 sky130_fd_sc_hd__decap_12 fill_0_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_12 ();
 sky130_fd_sc_hd__decap_12 fill_0_13 ();
 sky130_fd_sc_hd__decap_12 fill_0_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_15 ();
 sky130_fd_sc_hd__decap_12 fill_0_16 ();
 sky130_fd_sc_hd__decap_12 fill_0_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_18 ();
 sky130_fd_sc_hd__decap_12 fill_0_19 ();
 sky130_fd_sc_hd__decap_12 fill_0_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_0_21 ();
 sky130_fd_sc_hd__decap_8 fill_0_22 ();
 sky130_fd_sc_hd__decap_3 fill_0_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_0 ();
 sky130_fd_sc_hd__decap_12 fill_1_1 ();
 sky130_fd_sc_hd__decap_12 fill_1_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_3 ();
 sky130_fd_sc_hd__decap_12 fill_1_4 ();
 sky130_fd_sc_hd__decap_12 fill_1_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_6 ();
 sky130_fd_sc_hd__decap_12 fill_1_7 ();
 sky130_fd_sc_hd__decap_12 fill_1_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_9 ();
 sky130_fd_sc_hd__decap_12 fill_1_10 ();
 sky130_fd_sc_hd__decap_12 fill_1_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_12 ();
 sky130_fd_sc_hd__decap_12 fill_1_13 ();
 sky130_fd_sc_hd__decap_12 fill_1_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_15 ();
 sky130_fd_sc_hd__decap_12 fill_1_16 ();
 sky130_fd_sc_hd__decap_12 fill_1_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_18 ();
 sky130_fd_sc_hd__decap_12 fill_1_19 ();
 sky130_fd_sc_hd__decap_12 fill_1_20 ();
 sky130_fd_sc_hd__decap_6 fill_1_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_1_22 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_2_1 ();
 sky130_fd_sc_hd__decap_6 fill_2_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_3_0 ();
 sky130_fd_sc_hd__decap_6 fill_3_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_3_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_4_1 ();
 sky130_fd_sc_hd__decap_8 fill_4_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_5_0 ();
 sky130_fd_sc_hd__decap_8 fill_5_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_6_1 ();
 sky130_fd_sc_hd__decap_12 fill_6_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_7_2 ();
 sky130_fd_sc_hd__decap_6 fill_7_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_7_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_8_3 ();
 sky130_fd_sc_hd__decap_3 fill_8_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_9_2 ();
 sky130_fd_sc_hd__decap_6 fill_9_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_11_0 ();
 sky130_fd_sc_hd__decap_4 fill_11_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_11_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_12_1 ();
 sky130_fd_sc_hd__decap_6 fill_12_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_13_0 ();
 sky130_fd_sc_hd__decap_8 fill_13_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_14_1 ();
 sky130_fd_sc_hd__decap_12 fill_14_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_15_2 ();
 sky130_fd_sc_hd__decap_8 fill_15_3 ();
 sky130_fd_sc_hd__decap_3 fill_15_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_3 ();
 sky130_fd_sc_hd__decap_12 fill_16_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_16_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_17_2 ();
 sky130_fd_sc_hd__decap_12 fill_17_3 ();
 sky130_fd_sc_hd__decap_6 fill_17_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_18_1 ();
 sky130_fd_sc_hd__decap_8 fill_18_2 ();
 sky130_fd_sc_hd__fill_2 fill_18_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_19_0 ();
 sky130_fd_sc_hd__decap_12 fill_19_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_20_1 ();
 sky130_fd_sc_hd__decap_12 fill_20_2 ();
 sky130_fd_sc_hd__decap_4 fill_20_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_21_0 ();
 sky130_fd_sc_hd__decap_12 fill_21_1 ();
 sky130_fd_sc_hd__decap_4 fill_21_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_21_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_22_1 ();
 sky130_fd_sc_hd__decap_12 fill_22_2 ();
 sky130_fd_sc_hd__decap_8 fill_22_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_23_2 ();
 sky130_fd_sc_hd__decap_12 fill_23_3 ();
 sky130_fd_sc_hd__decap_8 fill_23_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_23_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_3 ();
 sky130_fd_sc_hd__decap_12 fill_24_4 ();
 sky130_fd_sc_hd__decap_8 fill_24_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_24_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_25_2 ();
 sky130_fd_sc_hd__decap_12 fill_25_3 ();
 sky130_fd_sc_hd__decap_8 fill_25_4 ();
 sky130_fd_sc_hd__fill_2 fill_25_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_26_1 ();
 sky130_fd_sc_hd__decap_12 fill_26_2 ();
 sky130_fd_sc_hd__fill_2 fill_26_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_27_0 ();
 sky130_fd_sc_hd__decap_12 fill_27_1 ();
 sky130_fd_sc_hd__decap_4 fill_27_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_28_1 ();
 sky130_fd_sc_hd__decap_12 fill_28_2 ();
 sky130_fd_sc_hd__decap_4 fill_28_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_29_0 ();
 sky130_fd_sc_hd__decap_12 fill_29_1 ();
 sky130_fd_sc_hd__decap_4 fill_29_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_29_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_30_1 ();
 sky130_fd_sc_hd__decap_12 fill_30_2 ();
 sky130_fd_sc_hd__decap_8 fill_30_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_31_2 ();
 sky130_fd_sc_hd__decap_12 fill_31_3 ();
 sky130_fd_sc_hd__decap_8 fill_31_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_31_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_3 ();
 sky130_fd_sc_hd__decap_12 fill_32_4 ();
 sky130_fd_sc_hd__decap_8 fill_32_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_32_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_33_2 ();
 sky130_fd_sc_hd__decap_12 fill_33_3 ();
 sky130_fd_sc_hd__decap_8 fill_33_4 ();
 sky130_fd_sc_hd__fill_2 fill_33_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_0 ();
 sky130_fd_sc_hd__decap_12 fill_34_1 ();
 sky130_fd_sc_hd__decap_12 fill_34_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_3 ();
 sky130_fd_sc_hd__decap_12 fill_34_4 ();
 sky130_fd_sc_hd__decap_12 fill_34_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_6 ();
 sky130_fd_sc_hd__decap_12 fill_34_7 ();
 sky130_fd_sc_hd__decap_12 fill_34_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_9 ();
 sky130_fd_sc_hd__decap_12 fill_34_10 ();
 sky130_fd_sc_hd__decap_12 fill_34_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_12 ();
 sky130_fd_sc_hd__decap_12 fill_34_13 ();
 sky130_fd_sc_hd__decap_12 fill_34_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_15 ();
 sky130_fd_sc_hd__decap_12 fill_34_16 ();
 sky130_fd_sc_hd__decap_12 fill_34_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_18 ();
 sky130_fd_sc_hd__decap_12 fill_34_19 ();
 sky130_fd_sc_hd__decap_12 fill_34_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_21 ();
 sky130_fd_sc_hd__decap_12 fill_34_22 ();
 sky130_fd_sc_hd__decap_12 fill_34_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_24 ();
 sky130_fd_sc_hd__decap_12 fill_34_25 ();
 sky130_fd_sc_hd__decap_12 fill_34_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_27 ();
 sky130_fd_sc_hd__decap_12 fill_34_28 ();
 sky130_fd_sc_hd__decap_12 fill_34_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_30 ();
 sky130_fd_sc_hd__decap_12 fill_34_31 ();
 sky130_fd_sc_hd__decap_12 fill_34_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_33 ();
 sky130_fd_sc_hd__decap_12 fill_34_34 ();
 sky130_fd_sc_hd__decap_12 fill_34_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_36 ();
 sky130_fd_sc_hd__decap_12 fill_34_37 ();
 sky130_fd_sc_hd__decap_12 fill_34_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_39 ();
 sky130_fd_sc_hd__decap_12 fill_34_40 ();
 sky130_fd_sc_hd__decap_12 fill_34_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_42 ();
 sky130_fd_sc_hd__decap_12 fill_34_43 ();
 sky130_fd_sc_hd__decap_12 fill_34_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_45 ();
 sky130_fd_sc_hd__decap_12 fill_34_46 ();
 sky130_fd_sc_hd__decap_12 fill_34_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_48 ();
 sky130_fd_sc_hd__decap_12 fill_34_49 ();
 sky130_fd_sc_hd__decap_12 fill_34_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_51 ();
 sky130_fd_sc_hd__decap_12 fill_34_52 ();
 sky130_fd_sc_hd__decap_12 fill_34_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_54 ();
 sky130_fd_sc_hd__decap_12 fill_34_55 ();
 sky130_fd_sc_hd__decap_12 fill_34_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_57 ();
 sky130_fd_sc_hd__decap_12 fill_34_58 ();
 sky130_fd_sc_hd__decap_12 fill_34_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_60 ();
 sky130_fd_sc_hd__decap_12 fill_34_61 ();
 sky130_fd_sc_hd__decap_12 fill_34_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_34_63 ();
 sky130_fd_sc_hd__decap_12 fill_34_64 ();
 sky130_fd_sc_hd__decap_12 fill_34_65 ();
 sky130_fd_sc_hd__fill_2 fill_34_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_0 ();
 sky130_fd_sc_hd__decap_12 fill_35_1 ();
 sky130_fd_sc_hd__decap_12 fill_35_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_3 ();
 sky130_fd_sc_hd__decap_12 fill_35_4 ();
 sky130_fd_sc_hd__decap_12 fill_35_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_6 ();
 sky130_fd_sc_hd__decap_12 fill_35_7 ();
 sky130_fd_sc_hd__decap_12 fill_35_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_9 ();
 sky130_fd_sc_hd__decap_12 fill_35_10 ();
 sky130_fd_sc_hd__decap_12 fill_35_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_12 ();
 sky130_fd_sc_hd__decap_12 fill_35_13 ();
 sky130_fd_sc_hd__decap_12 fill_35_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_15 ();
 sky130_fd_sc_hd__decap_12 fill_35_16 ();
 sky130_fd_sc_hd__decap_12 fill_35_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_18 ();
 sky130_fd_sc_hd__decap_12 fill_35_19 ();
 sky130_fd_sc_hd__decap_12 fill_35_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_21 ();
 sky130_fd_sc_hd__decap_12 fill_35_22 ();
 sky130_fd_sc_hd__decap_12 fill_35_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_35_24 ();
 sky130_fd_sc_hd__decap_12 fill_35_25 ();
 sky130_fd_sc_hd__decap_8 fill_35_26 ();
 sky130_fd_sc_hd__decap_3 fill_35_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_36_0 ();
 sky130_fd_sc_hd__decap_12 fill_36_1 ();
 sky130_fd_sc_hd__decap_12 fill_36_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_36_3 ();
 sky130_fd_sc_hd__decap_12 fill_36_4 ();
 sky130_fd_sc_hd__decap_12 fill_36_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_36_6 ();
 sky130_fd_sc_hd__decap_12 fill_36_7 ();
 sky130_fd_sc_hd__decap_12 fill_36_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_36_9 ();
 sky130_fd_sc_hd__decap_12 fill_36_10 ();
 sky130_fd_sc_hd__decap_12 fill_36_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_36_12 ();
 sky130_fd_sc_hd__decap_12 fill_36_13 ();
 sky130_fd_sc_hd__decap_12 fill_36_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_36_15 ();
 sky130_fd_sc_hd__decap_12 fill_36_16 ();
 sky130_fd_sc_hd__decap_12 fill_36_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_36_18 ();
 sky130_fd_sc_hd__decap_12 fill_36_19 ();
 sky130_fd_sc_hd__decap_12 fill_36_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_36_21 ();
 sky130_fd_sc_hd__decap_8 fill_36_22 ();
 sky130_fd_sc_hd__decap_3 fill_36_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_0 ();
 sky130_fd_sc_hd__decap_8 fill_37_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_37_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_38_1 ();
 sky130_fd_sc_hd__decap_12 fill_38_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_39_0 ();
 sky130_fd_sc_hd__decap_12 fill_39_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_40_1 ();
 sky130_fd_sc_hd__decap_12 fill_40_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_40_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_41_0 ();
 sky130_fd_sc_hd__decap_12 fill_41_1 ();
 sky130_fd_sc_hd__decap_4 fill_41_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_42_3 ();
 sky130_fd_sc_hd__decap_8 fill_42_4 ();
 sky130_fd_sc_hd__decap_3 fill_42_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_43_2 ();
 sky130_fd_sc_hd__decap_12 fill_43_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_43_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_44_3 ();
 sky130_fd_sc_hd__decap_12 fill_44_4 ();
 sky130_fd_sc_hd__fill_2 fill_44_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_45_0 ();
 sky130_fd_sc_hd__decap_6 fill_45_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_45_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_46_1 ();
 sky130_fd_sc_hd__decap_12 fill_46_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_47_0 ();
 sky130_fd_sc_hd__decap_12 fill_47_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_48_1 ();
 sky130_fd_sc_hd__decap_12 fill_48_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_48_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_49_0 ();
 sky130_fd_sc_hd__decap_12 fill_49_1 ();
 sky130_fd_sc_hd__decap_4 fill_49_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_50_3 ();
 sky130_fd_sc_hd__decap_12 fill_50_4 ();
 sky130_fd_sc_hd__decap_3 fill_50_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_51_2 ();
 sky130_fd_sc_hd__decap_12 fill_51_3 ();
 sky130_fd_sc_hd__decap_4 fill_51_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_51_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_52_3 ();
 sky130_fd_sc_hd__decap_12 fill_52_4 ();
 sky130_fd_sc_hd__decap_6 fill_52_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_53_0 ();
 sky130_fd_sc_hd__decap_8 fill_53_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_53_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_54_1 ();
 sky130_fd_sc_hd__decap_12 fill_54_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_55_0 ();
 sky130_fd_sc_hd__decap_12 fill_55_1 ();
 sky130_fd_sc_hd__decap_4 fill_55_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_56_1 ();
 sky130_fd_sc_hd__decap_12 fill_56_2 ();
 sky130_fd_sc_hd__decap_4 fill_56_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_56_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_57_0 ();
 sky130_fd_sc_hd__decap_12 fill_57_1 ();
 sky130_fd_sc_hd__decap_8 fill_57_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_58_3 ();
 sky130_fd_sc_hd__decap_12 fill_58_4 ();
 sky130_fd_sc_hd__decap_8 fill_58_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_58_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_59_2 ();
 sky130_fd_sc_hd__decap_12 fill_59_3 ();
 sky130_fd_sc_hd__decap_8 fill_59_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_59_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_60_3 ();
 sky130_fd_sc_hd__decap_12 fill_60_4 ();
 sky130_fd_sc_hd__decap_8 fill_60_5 ();
 sky130_fd_sc_hd__fill_2 fill_60_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_61_0 ();
 sky130_fd_sc_hd__decap_12 fill_61_1 ();
 sky130_fd_sc_hd__fill_2 fill_61_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_62_1 ();
 sky130_fd_sc_hd__decap_12 fill_62_2 ();
 sky130_fd_sc_hd__decap_4 fill_62_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_63_0 ();
 sky130_fd_sc_hd__decap_12 fill_63_1 ();
 sky130_fd_sc_hd__decap_4 fill_63_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_64_1 ();
 sky130_fd_sc_hd__decap_12 fill_64_2 ();
 sky130_fd_sc_hd__decap_4 fill_64_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_64_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_65_0 ();
 sky130_fd_sc_hd__decap_12 fill_65_1 ();
 sky130_fd_sc_hd__decap_8 fill_65_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_66_3 ();
 sky130_fd_sc_hd__decap_12 fill_66_4 ();
 sky130_fd_sc_hd__decap_8 fill_66_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_66_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_67_2 ();
 sky130_fd_sc_hd__decap_12 fill_67_3 ();
 sky130_fd_sc_hd__decap_8 fill_67_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_67_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_68_3 ();
 sky130_fd_sc_hd__decap_12 fill_68_4 ();
 sky130_fd_sc_hd__decap_8 fill_68_5 ();
 sky130_fd_sc_hd__fill_2 fill_68_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_0 ();
 sky130_fd_sc_hd__decap_12 fill_69_1 ();
 sky130_fd_sc_hd__decap_12 fill_69_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_3 ();
 sky130_fd_sc_hd__decap_12 fill_69_4 ();
 sky130_fd_sc_hd__decap_12 fill_69_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_6 ();
 sky130_fd_sc_hd__decap_12 fill_69_7 ();
 sky130_fd_sc_hd__decap_12 fill_69_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_9 ();
 sky130_fd_sc_hd__decap_12 fill_69_10 ();
 sky130_fd_sc_hd__decap_12 fill_69_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_12 ();
 sky130_fd_sc_hd__decap_12 fill_69_13 ();
 sky130_fd_sc_hd__decap_12 fill_69_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_15 ();
 sky130_fd_sc_hd__decap_12 fill_69_16 ();
 sky130_fd_sc_hd__decap_12 fill_69_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_18 ();
 sky130_fd_sc_hd__decap_12 fill_69_19 ();
 sky130_fd_sc_hd__decap_12 fill_69_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_21 ();
 sky130_fd_sc_hd__decap_12 fill_69_22 ();
 sky130_fd_sc_hd__decap_12 fill_69_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_24 ();
 sky130_fd_sc_hd__decap_12 fill_69_25 ();
 sky130_fd_sc_hd__decap_12 fill_69_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_27 ();
 sky130_fd_sc_hd__decap_12 fill_69_28 ();
 sky130_fd_sc_hd__decap_12 fill_69_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_30 ();
 sky130_fd_sc_hd__decap_12 fill_69_31 ();
 sky130_fd_sc_hd__decap_12 fill_69_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_33 ();
 sky130_fd_sc_hd__decap_12 fill_69_34 ();
 sky130_fd_sc_hd__decap_12 fill_69_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_36 ();
 sky130_fd_sc_hd__decap_12 fill_69_37 ();
 sky130_fd_sc_hd__decap_12 fill_69_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_39 ();
 sky130_fd_sc_hd__decap_12 fill_69_40 ();
 sky130_fd_sc_hd__decap_12 fill_69_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_42 ();
 sky130_fd_sc_hd__decap_12 fill_69_43 ();
 sky130_fd_sc_hd__decap_12 fill_69_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_45 ();
 sky130_fd_sc_hd__decap_12 fill_69_46 ();
 sky130_fd_sc_hd__decap_12 fill_69_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_48 ();
 sky130_fd_sc_hd__decap_12 fill_69_49 ();
 sky130_fd_sc_hd__decap_12 fill_69_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_51 ();
 sky130_fd_sc_hd__decap_12 fill_69_52 ();
 sky130_fd_sc_hd__decap_12 fill_69_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_54 ();
 sky130_fd_sc_hd__decap_12 fill_69_55 ();
 sky130_fd_sc_hd__decap_12 fill_69_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_57 ();
 sky130_fd_sc_hd__decap_12 fill_69_58 ();
 sky130_fd_sc_hd__decap_12 fill_69_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_60 ();
 sky130_fd_sc_hd__decap_12 fill_69_61 ();
 sky130_fd_sc_hd__decap_12 fill_69_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_63 ();
 sky130_fd_sc_hd__decap_12 fill_69_64 ();
 sky130_fd_sc_hd__decap_12 fill_69_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_69_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_70_0 ();
 sky130_fd_sc_hd__decap_12 fill_70_1 ();
 sky130_fd_sc_hd__decap_12 fill_70_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_70_3 ();
 sky130_fd_sc_hd__decap_12 fill_70_4 ();
 sky130_fd_sc_hd__decap_12 fill_70_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_70_6 ();
 sky130_fd_sc_hd__decap_12 fill_70_7 ();
 sky130_fd_sc_hd__decap_12 fill_70_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_70_9 ();
 sky130_fd_sc_hd__decap_12 fill_70_10 ();
 sky130_fd_sc_hd__decap_12 fill_70_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_70_12 ();
 sky130_fd_sc_hd__decap_12 fill_70_13 ();
 sky130_fd_sc_hd__decap_12 fill_70_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_70_15 ();
 sky130_fd_sc_hd__decap_12 fill_70_16 ();
 sky130_fd_sc_hd__decap_12 fill_70_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_70_18 ();
 sky130_fd_sc_hd__decap_12 fill_70_19 ();
 sky130_fd_sc_hd__decap_12 fill_70_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_70_21 ();
 sky130_fd_sc_hd__decap_12 fill_70_22 ();
 sky130_fd_sc_hd__decap_12 fill_70_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_70_24 ();
 sky130_fd_sc_hd__decap_12 fill_70_25 ();
 sky130_fd_sc_hd__decap_12 fill_70_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_71_0 ();
 sky130_fd_sc_hd__decap_12 fill_71_1 ();
 sky130_fd_sc_hd__decap_12 fill_71_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_71_3 ();
 sky130_fd_sc_hd__decap_12 fill_71_4 ();
 sky130_fd_sc_hd__decap_12 fill_71_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_71_6 ();
 sky130_fd_sc_hd__decap_12 fill_71_7 ();
 sky130_fd_sc_hd__decap_12 fill_71_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_71_9 ();
 sky130_fd_sc_hd__decap_12 fill_71_10 ();
 sky130_fd_sc_hd__decap_12 fill_71_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_71_12 ();
 sky130_fd_sc_hd__decap_12 fill_71_13 ();
 sky130_fd_sc_hd__decap_12 fill_71_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_71_15 ();
 sky130_fd_sc_hd__decap_12 fill_71_16 ();
 sky130_fd_sc_hd__decap_12 fill_71_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_71_18 ();
 sky130_fd_sc_hd__decap_12 fill_71_19 ();
 sky130_fd_sc_hd__decap_12 fill_71_20 ();
 sky130_fd_sc_hd__decap_8 fill_71_21 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_71_22 ();
 sky130_fd_sc_hd__fill_2 fill_71_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_72_1 ();
 sky130_fd_sc_hd__decap_8 fill_72_2 ();
 sky130_fd_sc_hd__fill_2 fill_72_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_73_0 ();
 sky130_fd_sc_hd__decap_12 fill_73_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_74_1 ();
 sky130_fd_sc_hd__decap_12 fill_74_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_75_0 ();
 sky130_fd_sc_hd__decap_12 fill_75_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_75_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_76_1 ();
 sky130_fd_sc_hd__decap_12 fill_76_2 ();
 sky130_fd_sc_hd__decap_4 fill_76_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_77_2 ();
 sky130_fd_sc_hd__decap_8 fill_77_3 ();
 sky130_fd_sc_hd__decap_3 fill_77_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_78_3 ();
 sky130_fd_sc_hd__decap_12 fill_78_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_78_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_79_2 ();
 sky130_fd_sc_hd__decap_12 fill_79_3 ();
 sky130_fd_sc_hd__fill_2 fill_79_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_80_1 ();
 sky130_fd_sc_hd__decap_8 fill_80_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_81_0 ();
 sky130_fd_sc_hd__decap_12 fill_81_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_82_1 ();
 sky130_fd_sc_hd__decap_12 fill_82_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_83_0 ();
 sky130_fd_sc_hd__decap_12 fill_83_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_83_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_84_1 ();
 sky130_fd_sc_hd__decap_12 fill_84_2 ();
 sky130_fd_sc_hd__decap_4 fill_84_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_85_2 ();
 sky130_fd_sc_hd__decap_12 fill_85_3 ();
 sky130_fd_sc_hd__decap_3 fill_85_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_86_3 ();
 sky130_fd_sc_hd__decap_12 fill_86_4 ();
 sky130_fd_sc_hd__decap_4 fill_86_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_86_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_87_2 ();
 sky130_fd_sc_hd__decap_12 fill_87_3 ();
 sky130_fd_sc_hd__decap_6 fill_87_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_88_1 ();
 sky130_fd_sc_hd__decap_8 fill_88_2 ();
 sky130_fd_sc_hd__fill_2 fill_88_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_89_0 ();
 sky130_fd_sc_hd__decap_12 fill_89_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_90_1 ();
 sky130_fd_sc_hd__decap_12 fill_90_2 ();
 sky130_fd_sc_hd__decap_4 fill_90_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_91_0 ();
 sky130_fd_sc_hd__decap_12 fill_91_1 ();
 sky130_fd_sc_hd__decap_4 fill_91_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_91_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_92_1 ();
 sky130_fd_sc_hd__decap_12 fill_92_2 ();
 sky130_fd_sc_hd__decap_8 fill_92_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_93_2 ();
 sky130_fd_sc_hd__decap_12 fill_93_3 ();
 sky130_fd_sc_hd__decap_8 fill_93_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_93_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_94_3 ();
 sky130_fd_sc_hd__decap_12 fill_94_4 ();
 sky130_fd_sc_hd__decap_8 fill_94_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_94_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_95_2 ();
 sky130_fd_sc_hd__decap_12 fill_95_3 ();
 sky130_fd_sc_hd__decap_8 fill_95_4 ();
 sky130_fd_sc_hd__fill_2 fill_95_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_96_1 ();
 sky130_fd_sc_hd__decap_12 fill_96_2 ();
 sky130_fd_sc_hd__fill_2 fill_96_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_97_0 ();
 sky130_fd_sc_hd__decap_12 fill_97_1 ();
 sky130_fd_sc_hd__decap_4 fill_97_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_98_1 ();
 sky130_fd_sc_hd__decap_12 fill_98_2 ();
 sky130_fd_sc_hd__decap_4 fill_98_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_99_0 ();
 sky130_fd_sc_hd__decap_12 fill_99_1 ();
 sky130_fd_sc_hd__decap_4 fill_99_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_99_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_100_1 ();
 sky130_fd_sc_hd__decap_12 fill_100_2 ();
 sky130_fd_sc_hd__decap_8 fill_100_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_101_2 ();
 sky130_fd_sc_hd__decap_12 fill_101_3 ();
 sky130_fd_sc_hd__decap_8 fill_101_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_101_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_102_3 ();
 sky130_fd_sc_hd__decap_12 fill_102_4 ();
 sky130_fd_sc_hd__decap_8 fill_102_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_102_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_103_2 ();
 sky130_fd_sc_hd__decap_12 fill_103_3 ();
 sky130_fd_sc_hd__decap_8 fill_103_4 ();
 sky130_fd_sc_hd__fill_2 fill_103_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_0 ();
 sky130_fd_sc_hd__decap_12 fill_104_1 ();
 sky130_fd_sc_hd__decap_12 fill_104_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_3 ();
 sky130_fd_sc_hd__decap_12 fill_104_4 ();
 sky130_fd_sc_hd__decap_12 fill_104_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_6 ();
 sky130_fd_sc_hd__decap_12 fill_104_7 ();
 sky130_fd_sc_hd__decap_12 fill_104_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_9 ();
 sky130_fd_sc_hd__decap_12 fill_104_10 ();
 sky130_fd_sc_hd__decap_12 fill_104_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_12 ();
 sky130_fd_sc_hd__decap_12 fill_104_13 ();
 sky130_fd_sc_hd__decap_12 fill_104_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_15 ();
 sky130_fd_sc_hd__decap_12 fill_104_16 ();
 sky130_fd_sc_hd__decap_12 fill_104_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_18 ();
 sky130_fd_sc_hd__decap_12 fill_104_19 ();
 sky130_fd_sc_hd__decap_12 fill_104_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_21 ();
 sky130_fd_sc_hd__decap_12 fill_104_22 ();
 sky130_fd_sc_hd__decap_12 fill_104_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_24 ();
 sky130_fd_sc_hd__decap_12 fill_104_25 ();
 sky130_fd_sc_hd__decap_12 fill_104_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_27 ();
 sky130_fd_sc_hd__decap_12 fill_104_28 ();
 sky130_fd_sc_hd__decap_12 fill_104_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_30 ();
 sky130_fd_sc_hd__decap_12 fill_104_31 ();
 sky130_fd_sc_hd__decap_12 fill_104_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_33 ();
 sky130_fd_sc_hd__decap_12 fill_104_34 ();
 sky130_fd_sc_hd__decap_12 fill_104_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_36 ();
 sky130_fd_sc_hd__decap_12 fill_104_37 ();
 sky130_fd_sc_hd__decap_12 fill_104_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_39 ();
 sky130_fd_sc_hd__decap_12 fill_104_40 ();
 sky130_fd_sc_hd__decap_12 fill_104_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_42 ();
 sky130_fd_sc_hd__decap_12 fill_104_43 ();
 sky130_fd_sc_hd__decap_12 fill_104_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_45 ();
 sky130_fd_sc_hd__decap_12 fill_104_46 ();
 sky130_fd_sc_hd__decap_12 fill_104_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_48 ();
 sky130_fd_sc_hd__decap_12 fill_104_49 ();
 sky130_fd_sc_hd__decap_12 fill_104_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_51 ();
 sky130_fd_sc_hd__decap_12 fill_104_52 ();
 sky130_fd_sc_hd__decap_12 fill_104_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_54 ();
 sky130_fd_sc_hd__decap_12 fill_104_55 ();
 sky130_fd_sc_hd__decap_12 fill_104_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_57 ();
 sky130_fd_sc_hd__decap_12 fill_104_58 ();
 sky130_fd_sc_hd__decap_12 fill_104_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_60 ();
 sky130_fd_sc_hd__decap_12 fill_104_61 ();
 sky130_fd_sc_hd__decap_12 fill_104_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_104_63 ();
 sky130_fd_sc_hd__decap_12 fill_104_64 ();
 sky130_fd_sc_hd__decap_12 fill_104_65 ();
 sky130_fd_sc_hd__fill_2 fill_104_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_105_0 ();
 sky130_fd_sc_hd__decap_12 fill_105_1 ();
 sky130_fd_sc_hd__decap_12 fill_105_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_105_3 ();
 sky130_fd_sc_hd__decap_12 fill_105_4 ();
 sky130_fd_sc_hd__decap_12 fill_105_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_105_6 ();
 sky130_fd_sc_hd__decap_12 fill_105_7 ();
 sky130_fd_sc_hd__decap_12 fill_105_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_105_9 ();
 sky130_fd_sc_hd__decap_12 fill_105_10 ();
 sky130_fd_sc_hd__decap_12 fill_105_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_105_12 ();
 sky130_fd_sc_hd__decap_12 fill_105_13 ();
 sky130_fd_sc_hd__decap_12 fill_105_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_105_15 ();
 sky130_fd_sc_hd__decap_12 fill_105_16 ();
 sky130_fd_sc_hd__decap_12 fill_105_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_105_18 ();
 sky130_fd_sc_hd__decap_12 fill_105_19 ();
 sky130_fd_sc_hd__decap_12 fill_105_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_105_21 ();
 sky130_fd_sc_hd__decap_12 fill_105_22 ();
 sky130_fd_sc_hd__decap_12 fill_105_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_105_24 ();
 sky130_fd_sc_hd__decap_12 fill_105_25 ();
 sky130_fd_sc_hd__decap_8 fill_105_26 ();
 sky130_fd_sc_hd__decap_3 fill_105_27 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_106_0 ();
 sky130_fd_sc_hd__decap_12 fill_106_1 ();
 sky130_fd_sc_hd__decap_12 fill_106_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_106_3 ();
 sky130_fd_sc_hd__decap_12 fill_106_4 ();
 sky130_fd_sc_hd__decap_12 fill_106_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_106_6 ();
 sky130_fd_sc_hd__decap_12 fill_106_7 ();
 sky130_fd_sc_hd__decap_12 fill_106_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_106_9 ();
 sky130_fd_sc_hd__decap_12 fill_106_10 ();
 sky130_fd_sc_hd__decap_12 fill_106_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_106_12 ();
 sky130_fd_sc_hd__decap_12 fill_106_13 ();
 sky130_fd_sc_hd__decap_12 fill_106_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_106_15 ();
 sky130_fd_sc_hd__decap_12 fill_106_16 ();
 sky130_fd_sc_hd__decap_12 fill_106_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_106_18 ();
 sky130_fd_sc_hd__decap_12 fill_106_19 ();
 sky130_fd_sc_hd__decap_12 fill_106_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_106_21 ();
 sky130_fd_sc_hd__decap_8 fill_106_22 ();
 sky130_fd_sc_hd__decap_3 fill_106_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_107_0 ();
 sky130_fd_sc_hd__decap_8 fill_107_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_107_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_108_1 ();
 sky130_fd_sc_hd__decap_12 fill_108_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_109_0 ();
 sky130_fd_sc_hd__decap_12 fill_109_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_110_1 ();
 sky130_fd_sc_hd__decap_12 fill_110_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_110_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_111_0 ();
 sky130_fd_sc_hd__decap_12 fill_111_1 ();
 sky130_fd_sc_hd__decap_4 fill_111_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_112_3 ();
 sky130_fd_sc_hd__decap_8 fill_112_4 ();
 sky130_fd_sc_hd__decap_3 fill_112_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_113_2 ();
 sky130_fd_sc_hd__decap_12 fill_113_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_113_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_114_3 ();
 sky130_fd_sc_hd__decap_12 fill_114_4 ();
 sky130_fd_sc_hd__fill_2 fill_114_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_115_0 ();
 sky130_fd_sc_hd__decap_6 fill_115_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_115_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_116_1 ();
 sky130_fd_sc_hd__decap_12 fill_116_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_117_0 ();
 sky130_fd_sc_hd__decap_12 fill_117_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_118_1 ();
 sky130_fd_sc_hd__decap_12 fill_118_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_118_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_119_0 ();
 sky130_fd_sc_hd__decap_12 fill_119_1 ();
 sky130_fd_sc_hd__decap_4 fill_119_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_120_3 ();
 sky130_fd_sc_hd__decap_12 fill_120_4 ();
 sky130_fd_sc_hd__decap_3 fill_120_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_121_2 ();
 sky130_fd_sc_hd__decap_12 fill_121_3 ();
 sky130_fd_sc_hd__decap_4 fill_121_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_121_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_122_3 ();
 sky130_fd_sc_hd__decap_12 fill_122_4 ();
 sky130_fd_sc_hd__decap_6 fill_122_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_123_0 ();
 sky130_fd_sc_hd__decap_8 fill_123_1 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_123_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_124_1 ();
 sky130_fd_sc_hd__decap_12 fill_124_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_125_0 ();
 sky130_fd_sc_hd__decap_12 fill_125_1 ();
 sky130_fd_sc_hd__decap_4 fill_125_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_126_1 ();
 sky130_fd_sc_hd__decap_12 fill_126_2 ();
 sky130_fd_sc_hd__decap_4 fill_126_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_126_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_127_0 ();
 sky130_fd_sc_hd__decap_12 fill_127_1 ();
 sky130_fd_sc_hd__decap_8 fill_127_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_128_3 ();
 sky130_fd_sc_hd__decap_12 fill_128_4 ();
 sky130_fd_sc_hd__decap_8 fill_128_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_128_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_129_2 ();
 sky130_fd_sc_hd__decap_12 fill_129_3 ();
 sky130_fd_sc_hd__decap_8 fill_129_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_129_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_130_3 ();
 sky130_fd_sc_hd__decap_12 fill_130_4 ();
 sky130_fd_sc_hd__decap_8 fill_130_5 ();
 sky130_fd_sc_hd__fill_2 fill_130_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_131_0 ();
 sky130_fd_sc_hd__decap_12 fill_131_1 ();
 sky130_fd_sc_hd__fill_2 fill_131_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_132_1 ();
 sky130_fd_sc_hd__decap_12 fill_132_2 ();
 sky130_fd_sc_hd__decap_4 fill_132_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_133_0 ();
 sky130_fd_sc_hd__decap_12 fill_133_1 ();
 sky130_fd_sc_hd__decap_4 fill_133_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_134_1 ();
 sky130_fd_sc_hd__decap_12 fill_134_2 ();
 sky130_fd_sc_hd__decap_4 fill_134_3 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_134_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_135_0 ();
 sky130_fd_sc_hd__decap_12 fill_135_1 ();
 sky130_fd_sc_hd__decap_8 fill_135_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_136_3 ();
 sky130_fd_sc_hd__decap_12 fill_136_4 ();
 sky130_fd_sc_hd__decap_8 fill_136_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_136_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_137_2 ();
 sky130_fd_sc_hd__decap_12 fill_137_3 ();
 sky130_fd_sc_hd__decap_8 fill_137_4 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_137_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_138_3 ();
 sky130_fd_sc_hd__decap_12 fill_138_4 ();
 sky130_fd_sc_hd__decap_8 fill_138_5 ();
 sky130_fd_sc_hd__fill_2 fill_138_6 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_0 ();
 sky130_fd_sc_hd__decap_12 fill_139_1 ();
 sky130_fd_sc_hd__decap_12 fill_139_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_3 ();
 sky130_fd_sc_hd__decap_12 fill_139_4 ();
 sky130_fd_sc_hd__decap_12 fill_139_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_6 ();
 sky130_fd_sc_hd__decap_12 fill_139_7 ();
 sky130_fd_sc_hd__decap_12 fill_139_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_9 ();
 sky130_fd_sc_hd__decap_12 fill_139_10 ();
 sky130_fd_sc_hd__decap_12 fill_139_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_12 ();
 sky130_fd_sc_hd__decap_12 fill_139_13 ();
 sky130_fd_sc_hd__decap_12 fill_139_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_15 ();
 sky130_fd_sc_hd__decap_12 fill_139_16 ();
 sky130_fd_sc_hd__decap_12 fill_139_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_18 ();
 sky130_fd_sc_hd__decap_12 fill_139_19 ();
 sky130_fd_sc_hd__decap_12 fill_139_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_21 ();
 sky130_fd_sc_hd__decap_12 fill_139_22 ();
 sky130_fd_sc_hd__decap_12 fill_139_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_24 ();
 sky130_fd_sc_hd__decap_12 fill_139_25 ();
 sky130_fd_sc_hd__decap_12 fill_139_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_27 ();
 sky130_fd_sc_hd__decap_12 fill_139_28 ();
 sky130_fd_sc_hd__decap_12 fill_139_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_30 ();
 sky130_fd_sc_hd__decap_12 fill_139_31 ();
 sky130_fd_sc_hd__decap_12 fill_139_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_33 ();
 sky130_fd_sc_hd__decap_12 fill_139_34 ();
 sky130_fd_sc_hd__decap_12 fill_139_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_36 ();
 sky130_fd_sc_hd__decap_12 fill_139_37 ();
 sky130_fd_sc_hd__decap_12 fill_139_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_39 ();
 sky130_fd_sc_hd__decap_12 fill_139_40 ();
 sky130_fd_sc_hd__decap_12 fill_139_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_42 ();
 sky130_fd_sc_hd__decap_12 fill_139_43 ();
 sky130_fd_sc_hd__decap_12 fill_139_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_45 ();
 sky130_fd_sc_hd__decap_12 fill_139_46 ();
 sky130_fd_sc_hd__decap_12 fill_139_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_48 ();
 sky130_fd_sc_hd__decap_12 fill_139_49 ();
 sky130_fd_sc_hd__decap_12 fill_139_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_51 ();
 sky130_fd_sc_hd__decap_12 fill_139_52 ();
 sky130_fd_sc_hd__decap_12 fill_139_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_54 ();
 sky130_fd_sc_hd__decap_12 fill_139_55 ();
 sky130_fd_sc_hd__decap_12 fill_139_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_57 ();
 sky130_fd_sc_hd__decap_12 fill_139_58 ();
 sky130_fd_sc_hd__decap_12 fill_139_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_60 ();
 sky130_fd_sc_hd__decap_12 fill_139_61 ();
 sky130_fd_sc_hd__decap_12 fill_139_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_63 ();
 sky130_fd_sc_hd__decap_12 fill_139_64 ();
 sky130_fd_sc_hd__decap_12 fill_139_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_139_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_140_0 ();
 sky130_fd_sc_hd__decap_12 fill_140_1 ();
 sky130_fd_sc_hd__decap_12 fill_140_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_140_3 ();
 sky130_fd_sc_hd__decap_12 fill_140_4 ();
 sky130_fd_sc_hd__decap_12 fill_140_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_140_6 ();
 sky130_fd_sc_hd__decap_12 fill_140_7 ();
 sky130_fd_sc_hd__decap_12 fill_140_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_140_9 ();
 sky130_fd_sc_hd__decap_12 fill_140_10 ();
 sky130_fd_sc_hd__decap_12 fill_140_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_140_12 ();
 sky130_fd_sc_hd__decap_12 fill_140_13 ();
 sky130_fd_sc_hd__decap_12 fill_140_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_140_15 ();
 sky130_fd_sc_hd__decap_12 fill_140_16 ();
 sky130_fd_sc_hd__decap_12 fill_140_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_140_18 ();
 sky130_fd_sc_hd__decap_12 fill_140_19 ();
 sky130_fd_sc_hd__decap_12 fill_140_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_140_21 ();
 sky130_fd_sc_hd__decap_12 fill_140_22 ();
 sky130_fd_sc_hd__decap_12 fill_140_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_140_24 ();
 sky130_fd_sc_hd__decap_12 fill_140_25 ();
 sky130_fd_sc_hd__decap_12 fill_140_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_141_0 ();
 sky130_fd_sc_hd__decap_12 fill_141_1 ();
 sky130_fd_sc_hd__decap_12 fill_141_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_141_3 ();
 sky130_fd_sc_hd__decap_12 fill_141_4 ();
 sky130_fd_sc_hd__decap_12 fill_141_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_141_6 ();
 sky130_fd_sc_hd__decap_12 fill_141_7 ();
 sky130_fd_sc_hd__decap_12 fill_141_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_141_9 ();
 sky130_fd_sc_hd__decap_12 fill_141_10 ();
 sky130_fd_sc_hd__decap_12 fill_141_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_141_12 ();
 sky130_fd_sc_hd__decap_12 fill_141_13 ();
 sky130_fd_sc_hd__decap_8 fill_141_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_0 ();
 sky130_fd_sc_hd__decap_12 fill_142_1 ();
 sky130_fd_sc_hd__decap_12 fill_142_2 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_3 ();
 sky130_fd_sc_hd__decap_12 fill_142_4 ();
 sky130_fd_sc_hd__decap_12 fill_142_5 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_6 ();
 sky130_fd_sc_hd__decap_12 fill_142_7 ();
 sky130_fd_sc_hd__decap_12 fill_142_8 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_9 ();
 sky130_fd_sc_hd__decap_12 fill_142_10 ();
 sky130_fd_sc_hd__decap_12 fill_142_11 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_12 ();
 sky130_fd_sc_hd__decap_12 fill_142_13 ();
 sky130_fd_sc_hd__decap_12 fill_142_14 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_15 ();
 sky130_fd_sc_hd__decap_12 fill_142_16 ();
 sky130_fd_sc_hd__decap_12 fill_142_17 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_18 ();
 sky130_fd_sc_hd__decap_12 fill_142_19 ();
 sky130_fd_sc_hd__decap_12 fill_142_20 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_21 ();
 sky130_fd_sc_hd__decap_12 fill_142_22 ();
 sky130_fd_sc_hd__decap_12 fill_142_23 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_24 ();
 sky130_fd_sc_hd__decap_12 fill_142_25 ();
 sky130_fd_sc_hd__decap_12 fill_142_26 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_27 ();
 sky130_fd_sc_hd__decap_12 fill_142_28 ();
 sky130_fd_sc_hd__decap_12 fill_142_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_30 ();
 sky130_fd_sc_hd__decap_12 fill_142_31 ();
 sky130_fd_sc_hd__decap_12 fill_142_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_33 ();
 sky130_fd_sc_hd__decap_12 fill_142_34 ();
 sky130_fd_sc_hd__decap_12 fill_142_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_36 ();
 sky130_fd_sc_hd__decap_12 fill_142_37 ();
 sky130_fd_sc_hd__decap_12 fill_142_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_39 ();
 sky130_fd_sc_hd__decap_12 fill_142_40 ();
 sky130_fd_sc_hd__decap_12 fill_142_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_42 ();
 sky130_fd_sc_hd__decap_12 fill_142_43 ();
 sky130_fd_sc_hd__decap_12 fill_142_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_45 ();
 sky130_fd_sc_hd__decap_12 fill_142_46 ();
 sky130_fd_sc_hd__decap_12 fill_142_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_48 ();
 sky130_fd_sc_hd__decap_12 fill_142_49 ();
 sky130_fd_sc_hd__decap_12 fill_142_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_51 ();
 sky130_fd_sc_hd__decap_12 fill_142_52 ();
 sky130_fd_sc_hd__decap_12 fill_142_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_54 ();
 sky130_fd_sc_hd__decap_12 fill_142_55 ();
 sky130_fd_sc_hd__decap_12 fill_142_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_57 ();
 sky130_fd_sc_hd__decap_12 fill_142_58 ();
 sky130_fd_sc_hd__decap_12 fill_142_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_60 ();
 sky130_fd_sc_hd__decap_12 fill_142_61 ();
 sky130_fd_sc_hd__decap_12 fill_142_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_63 ();
 sky130_fd_sc_hd__decap_12 fill_142_64 ();
 sky130_fd_sc_hd__decap_12 fill_142_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_66 ();
 sky130_fd_sc_hd__decap_12 fill_142_67 ();
 sky130_fd_sc_hd__decap_12 fill_142_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 fill_142_69 ();
 sky130_fd_sc_hd__decap_12 fill_142_70 ();
 sky130_fd_sc_hd__decap_8 fill_142_71 ();
 sky130_fd_sc_hd__decap_3 fill_142_72 ();
endmodule

