magic
tech sky130A
magscale 1 2
timestamp 1638728696
<< metal1 >>
rect 129918 160760 129924 160812
rect 129976 160800 129982 160812
rect 134150 160800 134156 160812
rect 129976 160772 134156 160800
rect 129976 160760 129982 160772
rect 134150 160760 134156 160772
rect 134208 160760 134214 160812
rect 63402 160012 63408 160064
rect 63460 160052 63466 160064
rect 143258 160052 143264 160064
rect 63460 160024 143264 160052
rect 63460 160012 63466 160024
rect 143258 160012 143264 160024
rect 143316 160012 143322 160064
rect 143350 160012 143356 160064
rect 143408 160052 143414 160064
rect 156598 160052 156604 160064
rect 143408 160024 156604 160052
rect 143408 160012 143414 160024
rect 156598 160012 156604 160024
rect 156656 160012 156662 160064
rect 156782 160012 156788 160064
rect 156840 160052 156846 160064
rect 191742 160052 191748 160064
rect 156840 160024 191748 160052
rect 156840 160012 156846 160024
rect 191742 160012 191748 160024
rect 191800 160012 191806 160064
rect 197170 160012 197176 160064
rect 197228 160052 197234 160064
rect 207014 160052 207020 160064
rect 197228 160024 207020 160052
rect 197228 160012 197234 160024
rect 207014 160012 207020 160024
rect 207072 160012 207078 160064
rect 211430 160012 211436 160064
rect 211488 160052 211494 160064
rect 280338 160052 280344 160064
rect 211488 160024 280344 160052
rect 211488 160012 211494 160024
rect 280338 160012 280344 160024
rect 280396 160012 280402 160064
rect 281258 160012 281264 160064
rect 281316 160052 281322 160064
rect 332686 160052 332692 160064
rect 281316 160024 332692 160052
rect 281316 160012 281322 160024
rect 332686 160012 332692 160024
rect 332744 160012 332750 160064
rect 334250 160012 334256 160064
rect 334308 160052 334314 160064
rect 374086 160052 374092 160064
rect 334308 160024 374092 160052
rect 334308 160012 334314 160024
rect 374086 160012 374092 160024
rect 374144 160012 374150 160064
rect 378870 160012 378876 160064
rect 378928 160052 378934 160064
rect 398558 160052 398564 160064
rect 378928 160024 398564 160052
rect 378928 160012 378934 160024
rect 398558 160012 398564 160024
rect 398616 160012 398622 160064
rect 25590 159944 25596 159996
rect 25648 159984 25654 159996
rect 109770 159984 109776 159996
rect 25648 159956 109776 159984
rect 25648 159944 25654 159956
rect 109770 159944 109776 159956
rect 109828 159944 109834 159996
rect 117222 159944 117228 159996
rect 117280 159984 117286 159996
rect 191466 159984 191472 159996
rect 117280 159956 191472 159984
rect 117280 159944 117286 159956
rect 191466 159944 191472 159956
rect 191524 159944 191530 159996
rect 197998 159944 198004 159996
rect 198056 159984 198062 159996
rect 269114 159984 269120 159996
rect 198056 159956 269120 159984
rect 198056 159944 198062 159956
rect 269114 159944 269120 159956
rect 269172 159944 269178 159996
rect 271230 159944 271236 159996
rect 271288 159984 271294 159996
rect 271874 159984 271880 159996
rect 271288 159956 271880 159984
rect 271288 159944 271294 159956
rect 271874 159944 271880 159956
rect 271932 159944 271938 159996
rect 275370 159944 275376 159996
rect 275428 159984 275434 159996
rect 329098 159984 329104 159996
rect 275428 159956 329104 159984
rect 275428 159944 275434 159956
rect 329098 159944 329104 159956
rect 329156 159944 329162 159996
rect 329190 159944 329196 159996
rect 329248 159984 329254 159996
rect 369946 159984 369952 159996
rect 329248 159956 369952 159984
rect 329248 159944 329254 159956
rect 369946 159944 369952 159956
rect 370004 159944 370010 159996
rect 374638 159944 374644 159996
rect 374696 159984 374702 159996
rect 388162 159984 388168 159996
rect 374696 159956 388168 159984
rect 374696 159944 374702 159956
rect 388162 159944 388168 159956
rect 388220 159944 388226 159996
rect 389818 159944 389824 159996
rect 389876 159984 389882 159996
rect 413830 159984 413836 159996
rect 389876 159956 413836 159984
rect 389876 159944 389882 159956
rect 413830 159944 413836 159956
rect 413888 159944 413894 159996
rect 76926 159876 76932 159928
rect 76984 159916 76990 159928
rect 162486 159916 162492 159928
rect 76984 159888 162492 159916
rect 76984 159876 76990 159888
rect 162486 159876 162492 159888
rect 162544 159876 162550 159928
rect 166902 159876 166908 159928
rect 166960 159916 166966 159928
rect 186682 159916 186688 159928
rect 166960 159888 186688 159916
rect 166960 159876 166966 159888
rect 186682 159876 186688 159888
rect 186740 159876 186746 159928
rect 191282 159876 191288 159928
rect 191340 159916 191346 159928
rect 264882 159916 264888 159928
rect 191340 159888 264888 159916
rect 191340 159876 191346 159888
rect 264882 159876 264888 159888
rect 264940 159876 264946 159928
rect 268654 159876 268660 159928
rect 268712 159916 268718 159928
rect 324038 159916 324044 159928
rect 268712 159888 324044 159916
rect 268712 159876 268718 159888
rect 324038 159876 324044 159888
rect 324096 159876 324102 159928
rect 328362 159876 328368 159928
rect 328420 159916 328426 159928
rect 369486 159916 369492 159928
rect 328420 159888 369492 159916
rect 328420 159876 328426 159888
rect 369486 159876 369492 159888
rect 369544 159876 369550 159928
rect 372154 159876 372160 159928
rect 372212 159916 372218 159928
rect 396166 159916 396172 159928
rect 372212 159888 396172 159916
rect 372212 159876 372218 159888
rect 396166 159876 396172 159888
rect 396224 159876 396230 159928
rect 403250 159876 403256 159928
rect 403308 159916 403314 159928
rect 416590 159916 416596 159928
rect 403308 159888 416596 159916
rect 403308 159876 403314 159888
rect 416590 159876 416596 159888
rect 416648 159876 416654 159928
rect 476114 159916 476120 159928
rect 470566 159888 476120 159916
rect 470566 159860 470594 159888
rect 476114 159876 476120 159888
rect 476172 159876 476178 159928
rect 480622 159876 480628 159928
rect 480680 159916 480686 159928
rect 485958 159916 485964 159928
rect 480680 159888 485964 159916
rect 480680 159876 480686 159888
rect 485958 159876 485964 159888
rect 486016 159876 486022 159928
rect 56686 159808 56692 159860
rect 56744 159848 56750 159860
rect 132954 159848 132960 159860
rect 56744 159820 132960 159848
rect 56744 159808 56750 159820
rect 132954 159808 132960 159820
rect 133012 159808 133018 159860
rect 133138 159808 133144 159860
rect 133196 159848 133202 159860
rect 143166 159848 143172 159860
rect 133196 159820 143172 159848
rect 133196 159808 133202 159820
rect 143166 159808 143172 159820
rect 143224 159808 143230 159860
rect 143258 159808 143264 159860
rect 143316 159848 143322 159860
rect 146570 159848 146576 159860
rect 143316 159820 146576 159848
rect 143316 159808 143322 159820
rect 146570 159808 146576 159820
rect 146628 159808 146634 159860
rect 146662 159808 146668 159860
rect 146720 159848 146726 159860
rect 176654 159848 176660 159860
rect 146720 159820 176660 159848
rect 146720 159808 146726 159820
rect 176654 159808 176660 159820
rect 176712 159808 176718 159860
rect 184566 159808 184572 159860
rect 184624 159848 184630 159860
rect 259546 159848 259552 159860
rect 184624 159820 259552 159848
rect 184624 159808 184630 159820
rect 259546 159808 259552 159820
rect 259604 159808 259610 159860
rect 261938 159808 261944 159860
rect 261996 159848 262002 159860
rect 318886 159848 318892 159860
rect 261996 159820 318892 159848
rect 261996 159808 262002 159820
rect 318886 159808 318892 159820
rect 318944 159808 318950 159860
rect 320818 159808 320824 159860
rect 320876 159848 320882 159860
rect 362954 159848 362960 159860
rect 320876 159820 362960 159848
rect 320876 159808 320882 159820
rect 362954 159808 362960 159820
rect 363012 159808 363018 159860
rect 376294 159808 376300 159860
rect 376352 159848 376358 159860
rect 406194 159848 406200 159860
rect 376352 159820 406200 159848
rect 376352 159808 376358 159820
rect 406194 159808 406200 159820
rect 406252 159808 406258 159860
rect 409966 159808 409972 159860
rect 410024 159848 410030 159860
rect 417878 159848 417884 159860
rect 410024 159820 417884 159848
rect 410024 159808 410030 159820
rect 417878 159808 417884 159820
rect 417936 159808 417942 159860
rect 424318 159808 424324 159860
rect 424376 159848 424382 159860
rect 442810 159848 442816 159860
rect 424376 159820 442816 159848
rect 424376 159808 424382 159820
rect 442810 159808 442816 159820
rect 442868 159808 442874 159860
rect 446122 159808 446128 159860
rect 446180 159848 446186 159860
rect 456794 159848 456800 159860
rect 446180 159820 456800 159848
rect 446180 159808 446186 159820
rect 456794 159808 456800 159820
rect 456852 159808 456858 159860
rect 458726 159808 458732 159860
rect 458784 159848 458790 159860
rect 465074 159848 465080 159860
rect 458784 159820 465080 159848
rect 458784 159808 458790 159820
rect 465074 159808 465080 159820
rect 465132 159808 465138 159860
rect 470502 159808 470508 159860
rect 470560 159820 470594 159860
rect 470560 159808 470566 159820
rect 471422 159808 471428 159860
rect 471480 159848 471486 159860
rect 477678 159848 477684 159860
rect 471480 159820 477684 159848
rect 471480 159808 471486 159820
rect 477678 159808 477684 159820
rect 477736 159808 477742 159860
rect 70118 159740 70124 159792
rect 70176 159780 70182 159792
rect 156322 159780 156328 159792
rect 70176 159752 156328 159780
rect 70176 159740 70182 159752
rect 156322 159740 156328 159752
rect 156380 159740 156386 159792
rect 156598 159740 156604 159792
rect 156656 159780 156662 159792
rect 160094 159780 160100 159792
rect 156656 159752 160100 159780
rect 156656 159740 156662 159752
rect 160094 159740 160100 159752
rect 160152 159740 160158 159792
rect 177850 159740 177856 159792
rect 177908 159780 177914 159792
rect 253934 159780 253940 159792
rect 177908 159752 253940 159780
rect 177908 159740 177914 159752
rect 253934 159740 253940 159752
rect 253992 159740 253998 159792
rect 255222 159740 255228 159792
rect 255280 159780 255286 159792
rect 313458 159780 313464 159792
rect 255280 159752 313464 159780
rect 255280 159740 255286 159752
rect 313458 159740 313464 159752
rect 313516 159740 313522 159792
rect 314102 159740 314108 159792
rect 314160 159780 314166 159792
rect 357986 159780 357992 159792
rect 314160 159752 357992 159780
rect 314160 159740 314166 159752
rect 357986 159740 357992 159752
rect 358044 159740 358050 159792
rect 365438 159740 365444 159792
rect 365496 159780 365502 159792
rect 395522 159780 395528 159792
rect 365496 159752 395528 159780
rect 365496 159740 365502 159752
rect 395522 159740 395528 159752
rect 395580 159740 395586 159792
rect 396534 159740 396540 159792
rect 396592 159780 396598 159792
rect 413922 159780 413928 159792
rect 396592 159752 413928 159780
rect 396592 159740 396598 159752
rect 413922 159740 413928 159752
rect 413980 159740 413986 159792
rect 420914 159740 420920 159792
rect 420972 159780 420978 159792
rect 440418 159780 440424 159792
rect 420972 159752 440424 159780
rect 420972 159740 420978 159752
rect 440418 159740 440424 159752
rect 440476 159740 440482 159792
rect 450354 159740 450360 159792
rect 450412 159780 450418 159792
rect 462314 159780 462320 159792
rect 450412 159752 462320 159780
rect 450412 159740 450418 159752
rect 462314 159740 462320 159752
rect 462372 159740 462378 159792
rect 473078 159740 473084 159792
rect 473136 159780 473142 159792
rect 480070 159780 480076 159792
rect 473136 159752 480076 159780
rect 473136 159740 473142 159752
rect 480070 159740 480076 159752
rect 480128 159740 480134 159792
rect 18874 159672 18880 159724
rect 18932 159712 18938 159724
rect 109126 159712 109132 159724
rect 18932 159684 109132 159712
rect 18932 159672 18938 159684
rect 109126 159672 109132 159684
rect 109184 159672 109190 159724
rect 113082 159672 113088 159724
rect 113140 159712 113146 159724
rect 126422 159712 126428 159724
rect 113140 159684 126428 159712
rect 113140 159672 113146 159684
rect 126422 159672 126428 159684
rect 126480 159672 126486 159724
rect 126514 159672 126520 159724
rect 126572 159712 126578 159724
rect 156506 159712 156512 159724
rect 126572 159684 156512 159712
rect 126572 159672 126578 159684
rect 156506 159672 156512 159684
rect 156564 159672 156570 159724
rect 163774 159712 163780 159724
rect 156616 159684 163780 159712
rect 49970 159604 49976 159656
rect 50028 159644 50034 159656
rect 132862 159644 132868 159656
rect 50028 159616 132868 159644
rect 50028 159604 50034 159616
rect 132862 159604 132868 159616
rect 132920 159604 132926 159656
rect 136542 159644 136548 159656
rect 132972 159616 136548 159644
rect 43254 159536 43260 159588
rect 43312 159576 43318 159588
rect 132972 159576 133000 159616
rect 136542 159604 136548 159616
rect 136600 159604 136606 159656
rect 136634 159604 136640 159656
rect 136692 159644 136698 159656
rect 139394 159644 139400 159656
rect 136692 159616 139400 159644
rect 136692 159604 136698 159616
rect 139394 159604 139400 159616
rect 139452 159604 139458 159656
rect 139946 159604 139952 159656
rect 140004 159644 140010 159656
rect 156616 159644 156644 159684
rect 163774 159672 163780 159684
rect 163832 159672 163838 159724
rect 167730 159672 167736 159724
rect 167788 159712 167794 159724
rect 246942 159712 246948 159724
rect 167788 159684 246948 159712
rect 167788 159672 167794 159684
rect 246942 159672 246948 159684
rect 247000 159672 247006 159724
rect 248506 159672 248512 159724
rect 248564 159712 248570 159724
rect 248564 159684 306374 159712
rect 248564 159672 248570 159684
rect 140004 159616 156644 159644
rect 140004 159604 140010 159616
rect 161014 159604 161020 159656
rect 161072 159644 161078 159656
rect 240318 159644 240324 159656
rect 161072 159616 240324 159644
rect 161072 159604 161078 159616
rect 240318 159604 240324 159616
rect 240376 159604 240382 159656
rect 244274 159604 244280 159656
rect 244332 159644 244338 159656
rect 305362 159644 305368 159656
rect 244332 159616 305368 159644
rect 244332 159604 244338 159616
rect 305362 159604 305368 159616
rect 305420 159604 305426 159656
rect 306346 159644 306374 159684
rect 308214 159672 308220 159724
rect 308272 159712 308278 159724
rect 342622 159712 342628 159724
rect 308272 159684 342628 159712
rect 308272 159672 308278 159684
rect 342622 159672 342628 159684
rect 342680 159672 342686 159724
rect 342714 159672 342720 159724
rect 342772 159712 342778 159724
rect 343818 159712 343824 159724
rect 342772 159684 343824 159712
rect 342772 159672 342778 159684
rect 343818 159672 343824 159684
rect 343876 159672 343882 159724
rect 347774 159672 347780 159724
rect 347832 159712 347838 159724
rect 378778 159712 378784 159724
rect 347832 159684 378784 159712
rect 347832 159672 347838 159684
rect 378778 159672 378784 159684
rect 378836 159672 378842 159724
rect 379698 159672 379704 159724
rect 379756 159712 379762 159724
rect 405826 159712 405832 159724
rect 379756 159684 405832 159712
rect 379756 159672 379762 159684
rect 405826 159672 405832 159684
rect 405884 159672 405890 159724
rect 417510 159672 417516 159724
rect 417568 159712 417574 159724
rect 437658 159712 437664 159724
rect 417568 159684 437664 159712
rect 417568 159672 417574 159684
rect 437658 159672 437664 159684
rect 437716 159672 437722 159724
rect 449526 159672 449532 159724
rect 449584 159712 449590 159724
rect 460934 159712 460940 159724
rect 449584 159684 460940 159712
rect 449584 159672 449590 159684
rect 460934 159672 460940 159684
rect 460992 159672 460998 159724
rect 463786 159672 463792 159724
rect 463844 159712 463850 159724
rect 471422 159712 471428 159724
rect 463844 159684 471428 159712
rect 463844 159672 463850 159684
rect 471422 159672 471428 159684
rect 471480 159672 471486 159724
rect 478966 159672 478972 159724
rect 479024 159712 479030 159724
rect 484670 159712 484676 159724
rect 479024 159684 484676 159712
rect 479024 159672 479030 159684
rect 484670 159672 484676 159684
rect 484728 159672 484734 159724
rect 308582 159644 308588 159656
rect 306346 159616 308588 159644
rect 308582 159604 308588 159616
rect 308640 159604 308646 159656
rect 309042 159604 309048 159656
rect 309100 159644 309106 159656
rect 341610 159644 341616 159656
rect 309100 159616 341616 159644
rect 309100 159604 309106 159616
rect 341610 159604 341616 159616
rect 341668 159604 341674 159656
rect 342456 159616 342668 159644
rect 43312 159548 133000 159576
rect 43312 159536 43318 159548
rect 134150 159536 134156 159588
rect 134208 159576 134214 159588
rect 154482 159576 154488 159588
rect 134208 159548 154488 159576
rect 134208 159536 134214 159548
rect 154482 159536 154488 159548
rect 154540 159536 154546 159588
rect 157610 159536 157616 159588
rect 157668 159576 157674 159588
rect 239306 159576 239312 159588
rect 157668 159548 239312 159576
rect 157668 159536 157674 159548
rect 239306 159536 239312 159548
rect 239364 159536 239370 159588
rect 250990 159536 250996 159588
rect 251048 159576 251054 159588
rect 310606 159576 310612 159588
rect 251048 159548 310612 159576
rect 251048 159536 251054 159548
rect 310606 159536 310612 159548
rect 310664 159536 310670 159588
rect 315758 159536 315764 159588
rect 315816 159576 315822 159588
rect 342456 159576 342484 159616
rect 315816 159548 342484 159576
rect 342640 159576 342668 159616
rect 342806 159604 342812 159656
rect 342864 159644 342870 159656
rect 354214 159644 354220 159656
rect 342864 159616 354220 159644
rect 342864 159604 342870 159616
rect 354214 159604 354220 159616
rect 354272 159604 354278 159656
rect 357802 159604 357808 159656
rect 357860 159644 357866 159656
rect 369210 159644 369216 159656
rect 357860 159616 369216 159644
rect 357860 159604 357866 159616
rect 369210 159604 369216 159616
rect 369268 159604 369274 159656
rect 369578 159604 369584 159656
rect 369636 159644 369642 159656
rect 401042 159644 401048 159656
rect 369636 159616 401048 159644
rect 369636 159604 369642 159616
rect 401042 159604 401048 159616
rect 401100 159604 401106 159656
rect 407482 159604 407488 159656
rect 407540 159644 407546 159656
rect 429930 159644 429936 159656
rect 407540 159616 429936 159644
rect 407540 159604 407546 159616
rect 429930 159604 429936 159616
rect 429988 159604 429994 159656
rect 453758 159604 453764 159656
rect 453816 159644 453822 159656
rect 465258 159644 465264 159656
rect 453816 159616 465264 159644
rect 453816 159604 453822 159616
rect 465258 159604 465264 159616
rect 465316 159604 465322 159656
rect 468018 159604 468024 159656
rect 468076 159644 468082 159656
rect 476022 159644 476028 159656
rect 468076 159616 476028 159644
rect 468076 159604 468082 159616
rect 476022 159604 476028 159616
rect 476080 159604 476086 159656
rect 479794 159604 479800 159656
rect 479852 159644 479858 159656
rect 485222 159644 485228 159656
rect 479852 159616 485228 159644
rect 479852 159604 479858 159616
rect 485222 159604 485228 159616
rect 485280 159604 485286 159656
rect 358906 159576 358912 159588
rect 342640 159548 358912 159576
rect 315816 159536 315822 159548
rect 358906 159536 358912 159548
rect 358964 159536 358970 159588
rect 362862 159536 362868 159588
rect 362920 159576 362926 159588
rect 394970 159576 394976 159588
rect 362920 159548 394976 159576
rect 362920 159536 362926 159548
rect 394970 159536 394976 159548
rect 395028 159536 395034 159588
rect 399018 159536 399024 159588
rect 399076 159576 399082 159588
rect 408494 159576 408500 159588
rect 399076 159548 408500 159576
rect 399076 159536 399082 159548
rect 408494 159536 408500 159548
rect 408552 159536 408558 159588
rect 410794 159536 410800 159588
rect 410852 159576 410858 159588
rect 432506 159576 432512 159588
rect 410852 159548 432512 159576
rect 410852 159536 410858 159548
rect 432506 159536 432512 159548
rect 432564 159536 432570 159588
rect 452010 159536 452016 159588
rect 452068 159576 452074 159588
rect 463970 159576 463976 159588
rect 452068 159548 463976 159576
rect 452068 159536 452074 159548
rect 463970 159536 463976 159548
rect 464028 159536 464034 159588
rect 467190 159536 467196 159588
rect 467248 159576 467254 159588
rect 473354 159576 473360 159588
rect 467248 159548 473360 159576
rect 467248 159536 467254 159548
rect 473354 159536 473360 159548
rect 473412 159536 473418 159588
rect 32306 159468 32312 159520
rect 32364 159508 32370 159520
rect 32364 159480 126376 159508
rect 32364 159468 32370 159480
rect 36538 159400 36544 159452
rect 36596 159440 36602 159452
rect 126238 159440 126244 159452
rect 36596 159412 126244 159440
rect 36596 159400 36602 159412
rect 126238 159400 126244 159412
rect 126296 159400 126302 159452
rect 126348 159440 126376 159480
rect 126422 159468 126428 159520
rect 126480 159508 126486 159520
rect 127618 159508 127624 159520
rect 126480 159480 127624 159508
rect 126480 159468 126486 159480
rect 127618 159468 127624 159480
rect 127676 159468 127682 159520
rect 133230 159468 133236 159520
rect 133288 159508 133294 159520
rect 144086 159508 144092 159520
rect 133288 159480 144092 159508
rect 133288 159468 133294 159480
rect 144086 159468 144092 159480
rect 144144 159468 144150 159520
rect 144178 159468 144184 159520
rect 144236 159508 144242 159520
rect 225322 159508 225328 159520
rect 144236 159480 225328 159508
rect 144236 159468 144242 159480
rect 225322 159468 225328 159480
rect 225380 159468 225386 159520
rect 230842 159468 230848 159520
rect 230900 159508 230906 159520
rect 293954 159508 293960 159520
rect 230900 159480 293960 159508
rect 230900 159468 230906 159480
rect 293954 159468 293960 159480
rect 294012 159468 294018 159520
rect 294782 159468 294788 159520
rect 294840 159508 294846 159520
rect 294840 159480 341564 159508
rect 294840 159468 294846 159480
rect 126790 159440 126796 159452
rect 126348 159412 126796 159440
rect 126790 159400 126796 159412
rect 126848 159400 126854 159452
rect 147766 159440 147772 159452
rect 128326 159412 147772 159440
rect 6270 159332 6276 159384
rect 6328 159372 6334 159384
rect 122834 159372 122840 159384
rect 6328 159344 122840 159372
rect 6328 159332 6334 159344
rect 122834 159332 122840 159344
rect 122892 159332 122898 159384
rect 123110 159332 123116 159384
rect 123168 159372 123174 159384
rect 128326 159372 128354 159412
rect 147766 159400 147772 159412
rect 147824 159400 147830 159452
rect 150894 159400 150900 159452
rect 150952 159440 150958 159452
rect 233234 159440 233240 159452
rect 150952 159412 233240 159440
rect 150952 159400 150958 159412
rect 233234 159400 233240 159412
rect 233292 159400 233298 159452
rect 234982 159400 234988 159452
rect 235040 159440 235046 159452
rect 298002 159440 298008 159452
rect 235040 159412 298008 159440
rect 235040 159400 235046 159412
rect 298002 159400 298008 159412
rect 298060 159400 298066 159452
rect 301498 159400 301504 159452
rect 301556 159440 301562 159452
rect 341426 159440 341432 159452
rect 301556 159412 341432 159440
rect 301556 159400 301562 159412
rect 341426 159400 341432 159412
rect 341484 159400 341490 159452
rect 341536 159440 341564 159480
rect 341610 159468 341616 159520
rect 341668 159508 341674 159520
rect 354858 159508 354864 159520
rect 341668 159480 354864 159508
rect 341668 159468 341674 159480
rect 354858 159468 354864 159480
rect 354916 159468 354922 159520
rect 356146 159468 356152 159520
rect 356204 159508 356210 159520
rect 390554 159508 390560 159520
rect 356204 159480 390560 159508
rect 356204 159468 356210 159480
rect 390554 159468 390560 159480
rect 390612 159468 390618 159520
rect 400766 159468 400772 159520
rect 400824 159508 400830 159520
rect 424870 159508 424876 159520
rect 400824 159480 424876 159508
rect 400824 159468 400830 159480
rect 424870 159468 424876 159480
rect 424928 159468 424934 159520
rect 459646 159468 459652 159520
rect 459704 159508 459710 159520
rect 466638 159508 466644 159520
rect 459704 159480 466644 159508
rect 459704 159468 459710 159480
rect 466638 159468 466644 159480
rect 466696 159468 466702 159520
rect 468846 159468 468852 159520
rect 468904 159508 468910 159520
rect 474826 159508 474832 159520
rect 468904 159480 474832 159508
rect 468904 159468 468910 159480
rect 474826 159468 474832 159480
rect 474884 159468 474890 159520
rect 477310 159468 477316 159520
rect 477368 159508 477374 159520
rect 483290 159508 483296 159520
rect 477368 159480 483296 159508
rect 477368 159468 477374 159480
rect 483290 159468 483296 159480
rect 483348 159468 483354 159520
rect 342254 159440 342260 159452
rect 341536 159412 342260 159440
rect 342254 159400 342260 159412
rect 342312 159400 342318 159452
rect 342346 159400 342352 159452
rect 342404 159440 342410 159452
rect 349338 159440 349344 159452
rect 342404 159412 349344 159440
rect 342404 159400 342410 159412
rect 349338 159400 349344 159412
rect 349396 159400 349402 159452
rect 358630 159400 358636 159452
rect 358688 159440 358694 159452
rect 392762 159440 392768 159452
rect 358688 159412 392768 159440
rect 358688 159400 358694 159412
rect 392762 159400 392768 159412
rect 392820 159400 392826 159452
rect 404078 159400 404084 159452
rect 404136 159440 404142 159452
rect 427354 159440 427360 159452
rect 404136 159412 427360 159440
rect 404136 159400 404142 159412
rect 427354 159400 427360 159412
rect 427412 159400 427418 159452
rect 427630 159400 427636 159452
rect 427688 159440 427694 159452
rect 445386 159440 445392 159452
rect 427688 159412 445392 159440
rect 427688 159400 427694 159412
rect 445386 159400 445392 159412
rect 445444 159400 445450 159452
rect 451182 159400 451188 159452
rect 451240 159440 451246 159452
rect 462866 159440 462872 159452
rect 451240 159412 462872 159440
rect 451240 159400 451246 159412
rect 462866 159400 462872 159412
rect 462924 159400 462930 159452
rect 518802 159400 518808 159452
rect 518860 159440 518866 159452
rect 522666 159440 522672 159452
rect 518860 159412 522672 159440
rect 518860 159400 518866 159412
rect 522666 159400 522672 159412
rect 522724 159400 522730 159452
rect 123168 159344 128354 159372
rect 123168 159332 123174 159344
rect 132678 159332 132684 159384
rect 132736 159372 132742 159384
rect 137094 159372 137100 159384
rect 132736 159344 137100 159372
rect 132736 159332 132742 159344
rect 137094 159332 137100 159344
rect 137152 159332 137158 159384
rect 137462 159332 137468 159384
rect 137520 159372 137526 159384
rect 223574 159372 223580 159384
rect 137520 159344 223580 159372
rect 137520 159332 137526 159344
rect 223574 159332 223580 159344
rect 223632 159332 223638 159384
rect 231670 159332 231676 159384
rect 231728 159372 231734 159384
rect 295518 159372 295524 159384
rect 231728 159344 295524 159372
rect 231728 159332 231734 159344
rect 295518 159332 295524 159344
rect 295576 159332 295582 159384
rect 295610 159332 295616 159384
rect 295668 159372 295674 159384
rect 342438 159372 342444 159384
rect 295668 159344 342444 159372
rect 295668 159332 295674 159344
rect 342438 159332 342444 159344
rect 342496 159332 342502 159384
rect 346026 159332 346032 159384
rect 346084 159372 346090 159384
rect 382826 159372 382832 159384
rect 346084 159344 382832 159372
rect 346084 159332 346090 159344
rect 382826 159332 382832 159344
rect 382884 159332 382890 159384
rect 383102 159332 383108 159384
rect 383160 159372 383166 159384
rect 411346 159372 411352 159384
rect 383160 159344 411352 159372
rect 383160 159332 383166 159344
rect 411346 159332 411352 159344
rect 411404 159332 411410 159384
rect 414198 159332 414204 159384
rect 414256 159372 414262 159384
rect 435082 159372 435088 159384
rect 414256 159344 435088 159372
rect 414256 159332 414262 159344
rect 435082 159332 435088 159344
rect 435140 159332 435146 159384
rect 448698 159332 448704 159384
rect 448756 159372 448762 159384
rect 461394 159372 461400 159384
rect 448756 159344 461400 159372
rect 448756 159332 448762 159344
rect 461394 159332 461400 159344
rect 461452 159332 461458 159384
rect 469674 159332 469680 159384
rect 469732 159372 469738 159384
rect 477402 159372 477408 159384
rect 469732 159344 477408 159372
rect 469732 159332 469738 159344
rect 477402 159332 477408 159344
rect 477460 159332 477466 159384
rect 478138 159332 478144 159384
rect 478196 159372 478202 159384
rect 483198 159372 483204 159384
rect 478196 159344 483204 159372
rect 478196 159332 478202 159344
rect 483198 159332 483204 159344
rect 483256 159332 483262 159384
rect 518710 159332 518716 159384
rect 518768 159372 518774 159384
rect 523494 159372 523500 159384
rect 518768 159344 523500 159372
rect 518768 159332 518774 159344
rect 523494 159332 523500 159344
rect 523552 159332 523558 159384
rect 73522 159264 73528 159316
rect 73580 159304 73586 159316
rect 80054 159304 80060 159316
rect 73580 159276 80060 159304
rect 73580 159264 73586 159276
rect 80054 159264 80060 159276
rect 80112 159264 80118 159316
rect 83642 159264 83648 159316
rect 83700 159304 83706 159316
rect 166994 159304 167000 159316
rect 83700 159276 167000 159304
rect 83700 159264 83706 159276
rect 166994 159264 167000 159276
rect 167052 159264 167058 159316
rect 170214 159264 170220 159316
rect 170272 159304 170278 159316
rect 195146 159304 195152 159316
rect 170272 159276 195152 159304
rect 170272 159264 170278 159276
rect 195146 159264 195152 159276
rect 195204 159264 195210 159316
rect 195238 159264 195244 159316
rect 195296 159304 195302 159316
rect 201310 159304 201316 159316
rect 195296 159276 201316 159304
rect 195296 159264 195302 159276
rect 201310 159264 201316 159276
rect 201368 159264 201374 159316
rect 201402 159264 201408 159316
rect 201460 159304 201466 159316
rect 212626 159304 212632 159316
rect 201460 159276 212632 159304
rect 201460 159264 201466 159276
rect 212626 159264 212632 159276
rect 212684 159264 212690 159316
rect 214006 159264 214012 159316
rect 214064 159304 214070 159316
rect 281534 159304 281540 159316
rect 214064 159276 281540 159304
rect 214064 159264 214070 159276
rect 281534 159264 281540 159276
rect 281592 159264 281598 159316
rect 282086 159264 282092 159316
rect 282144 159304 282150 159316
rect 334342 159304 334348 159316
rect 282144 159276 334348 159304
rect 282144 159264 282150 159276
rect 334342 159264 334348 159276
rect 334400 159264 334406 159316
rect 335078 159264 335084 159316
rect 335136 159304 335142 159316
rect 373994 159304 374000 159316
rect 335136 159276 374000 159304
rect 335136 159264 335142 159276
rect 373994 159264 374000 159276
rect 374052 159264 374058 159316
rect 374638 159264 374644 159316
rect 374696 159304 374702 159316
rect 382274 159304 382280 159316
rect 374696 159276 382280 159304
rect 374696 159264 374702 159276
rect 382274 159264 382280 159276
rect 382332 159264 382338 159316
rect 388990 159264 388996 159316
rect 389048 159304 389054 159316
rect 404262 159304 404268 159316
rect 389048 159276 404268 159304
rect 389048 159264 389054 159276
rect 404262 159264 404268 159276
rect 404320 159264 404326 159316
rect 457898 159264 457904 159316
rect 457956 159304 457962 159316
rect 464430 159304 464436 159316
rect 457956 159276 464436 159304
rect 457956 159264 457962 159276
rect 464430 159264 464436 159276
rect 464488 159264 464494 159316
rect 80238 159196 80244 159248
rect 80296 159236 80302 159248
rect 91094 159236 91100 159248
rect 80296 159208 91100 159236
rect 80296 159196 80302 159208
rect 91094 159196 91100 159208
rect 91152 159196 91158 159248
rect 100478 159196 100484 159248
rect 100536 159236 100542 159248
rect 184382 159236 184388 159248
rect 100536 159208 184388 159236
rect 100536 159196 100542 159208
rect 184382 159196 184388 159208
rect 184440 159196 184446 159248
rect 187050 159196 187056 159248
rect 187108 159236 187114 159248
rect 214650 159236 214656 159248
rect 187108 159208 214656 159236
rect 187108 159196 187114 159208
rect 214650 159196 214656 159208
rect 214708 159196 214714 159248
rect 218238 159196 218244 159248
rect 218296 159236 218302 159248
rect 284386 159236 284392 159248
rect 218296 159208 284392 159236
rect 218296 159196 218302 159208
rect 284386 159196 284392 159208
rect 284444 159196 284450 159248
rect 287974 159196 287980 159248
rect 288032 159236 288038 159248
rect 338758 159236 338764 159248
rect 288032 159208 338764 159236
rect 288032 159196 288038 159208
rect 338758 159196 338764 159208
rect 338816 159196 338822 159248
rect 339310 159196 339316 159248
rect 339368 159236 339374 159248
rect 377950 159236 377956 159248
rect 339368 159208 377956 159236
rect 339368 159196 339374 159208
rect 377950 159196 377956 159208
rect 378008 159196 378014 159248
rect 385494 159236 385500 159248
rect 379486 159208 385500 159236
rect 86954 159128 86960 159180
rect 87012 159168 87018 159180
rect 87012 159140 162992 159168
rect 87012 159128 87018 159140
rect 93670 159060 93676 159112
rect 93728 159100 93734 159112
rect 162854 159100 162860 159112
rect 93728 159072 162860 159100
rect 93728 159060 93734 159072
rect 162854 159060 162860 159072
rect 162912 159060 162918 159112
rect 162964 159100 162992 159140
rect 163038 159128 163044 159180
rect 163096 159168 163102 159180
rect 172146 159168 172152 159180
rect 163096 159140 172152 159168
rect 163096 159128 163102 159140
rect 172146 159128 172152 159140
rect 172204 159128 172210 159180
rect 173618 159128 173624 159180
rect 173676 159168 173682 159180
rect 193674 159168 193680 159180
rect 173676 159140 193680 159168
rect 173676 159128 173682 159140
rect 193674 159128 193680 159140
rect 193732 159128 193738 159180
rect 193766 159128 193772 159180
rect 193824 159168 193830 159180
rect 218054 159168 218060 159180
rect 193824 159140 218060 159168
rect 193824 159128 193830 159140
rect 218054 159128 218060 159140
rect 218112 159128 218118 159180
rect 224954 159128 224960 159180
rect 225012 159168 225018 159180
rect 290642 159168 290648 159180
rect 225012 159140 290648 159168
rect 225012 159128 225018 159140
rect 290642 159128 290648 159140
rect 290700 159128 290706 159180
rect 293954 159128 293960 159180
rect 294012 159168 294018 159180
rect 295150 159168 295156 159180
rect 294012 159140 295156 159168
rect 294012 159128 294018 159140
rect 295150 159128 295156 159140
rect 295208 159128 295214 159180
rect 302326 159128 302332 159180
rect 302384 159168 302390 159180
rect 302384 159140 340874 159168
rect 302384 159128 302390 159140
rect 169754 159100 169760 159112
rect 162964 159072 169760 159100
rect 169754 159060 169760 159072
rect 169812 159060 169818 159112
rect 171134 159060 171140 159112
rect 171192 159100 171198 159112
rect 173158 159100 173164 159112
rect 171192 159072 173164 159100
rect 171192 159060 171198 159072
rect 173158 159060 173164 159072
rect 173216 159060 173222 159112
rect 180334 159060 180340 159112
rect 180392 159100 180398 159112
rect 204898 159100 204904 159112
rect 180392 159072 204904 159100
rect 180392 159060 180398 159072
rect 204898 159060 204904 159072
rect 204956 159060 204962 159112
rect 220722 159060 220728 159112
rect 220780 159100 220786 159112
rect 283190 159100 283196 159112
rect 220780 159072 283196 159100
rect 220780 159060 220786 159072
rect 283190 159060 283196 159072
rect 283248 159060 283254 159112
rect 284662 159060 284668 159112
rect 284720 159100 284726 159112
rect 285766 159100 285772 159112
rect 284720 159072 285772 159100
rect 284720 159060 284726 159072
rect 285766 159060 285772 159072
rect 285824 159060 285830 159112
rect 288066 159100 288072 159112
rect 287026 159072 288072 159100
rect 107194 158992 107200 159044
rect 107252 159032 107258 159044
rect 183462 159032 183468 159044
rect 107252 159004 183468 159032
rect 107252 158992 107258 159004
rect 183462 158992 183468 159004
rect 183520 158992 183526 159044
rect 183738 158992 183744 159044
rect 183796 159032 183802 159044
rect 195238 159032 195244 159044
rect 183796 159004 195244 159032
rect 183796 158992 183802 159004
rect 195238 158992 195244 159004
rect 195296 158992 195302 159044
rect 203886 158992 203892 159044
rect 203944 159032 203950 159044
rect 213822 159032 213828 159044
rect 203944 159004 213828 159032
rect 203944 158992 203950 159004
rect 213822 158992 213828 159004
rect 213880 158992 213886 159044
rect 214834 158992 214840 159044
rect 214892 159032 214898 159044
rect 222102 159032 222108 159044
rect 214892 159004 222108 159032
rect 214892 158992 214898 159004
rect 222102 158992 222108 159004
rect 222160 158992 222166 159044
rect 224126 158992 224132 159044
rect 224184 159032 224190 159044
rect 287026 159032 287054 159072
rect 288066 159060 288072 159072
rect 288124 159060 288130 159112
rect 288894 159060 288900 159112
rect 288952 159100 288958 159112
rect 338298 159100 338304 159112
rect 288952 159072 338304 159100
rect 288952 159060 288958 159072
rect 338298 159060 338304 159072
rect 338356 159060 338362 159112
rect 338482 159060 338488 159112
rect 338540 159100 338546 159112
rect 339678 159100 339684 159112
rect 338540 159072 339684 159100
rect 338540 159060 338546 159072
rect 339678 159060 339684 159072
rect 339736 159060 339742 159112
rect 340846 159100 340874 159140
rect 341426 159128 341432 159180
rect 341484 159168 341490 159180
rect 345658 159168 345664 159180
rect 341484 159140 345664 159168
rect 341484 159128 341490 159140
rect 345658 159128 345664 159140
rect 345716 159128 345722 159180
rect 345750 159128 345756 159180
rect 345808 159168 345814 159180
rect 351822 159168 351828 159180
rect 345808 159140 351828 159168
rect 345808 159128 345814 159140
rect 351822 159128 351828 159140
rect 351880 159128 351886 159180
rect 351914 159128 351920 159180
rect 351972 159168 351978 159180
rect 379486 159168 379514 159208
rect 385494 159196 385500 159208
rect 385552 159196 385558 159248
rect 385586 159196 385592 159248
rect 385644 159236 385650 159248
rect 398834 159236 398840 159248
rect 385644 159208 398840 159236
rect 385644 159196 385650 159208
rect 398834 159196 398840 159208
rect 398892 159196 398898 159248
rect 457070 159196 457076 159248
rect 457128 159236 457134 159248
rect 464154 159236 464160 159248
rect 457128 159208 464160 159236
rect 457128 159196 457134 159208
rect 464154 159196 464160 159208
rect 464212 159196 464218 159248
rect 388438 159168 388444 159180
rect 351972 159140 379514 159168
rect 383626 159140 388444 159168
rect 351972 159128 351978 159140
rect 349246 159100 349252 159112
rect 340846 159072 349252 159100
rect 349246 159060 349252 159072
rect 349304 159060 349310 159112
rect 349338 159060 349344 159112
rect 349396 159100 349402 159112
rect 349396 159072 374868 159100
rect 349396 159060 349402 159072
rect 224184 159004 287054 159032
rect 224184 158992 224190 159004
rect 298094 158992 298100 159044
rect 298152 159032 298158 159044
rect 300394 159032 300400 159044
rect 298152 159004 300400 159032
rect 298152 158992 298158 159004
rect 300394 158992 300400 159004
rect 300452 158992 300458 159044
rect 307386 158992 307392 159044
rect 307444 159032 307450 159044
rect 345566 159032 345572 159044
rect 307444 159004 345572 159032
rect 307444 158992 307450 159004
rect 345566 158992 345572 159004
rect 345624 158992 345630 159044
rect 345842 158992 345848 159044
rect 345900 159032 345906 159044
rect 349062 159032 349068 159044
rect 345900 159004 349068 159032
rect 345900 158992 345906 159004
rect 349062 158992 349068 159004
rect 349120 158992 349126 159044
rect 351086 158992 351092 159044
rect 351144 159032 351150 159044
rect 374638 159032 374644 159044
rect 351144 159004 374644 159032
rect 351144 158992 351150 159004
rect 374638 158992 374644 159004
rect 374696 158992 374702 159044
rect 374840 159032 374868 159072
rect 378042 159060 378048 159112
rect 378100 159100 378106 159112
rect 383626 159100 383654 159140
rect 388438 159128 388444 159140
rect 388496 159128 388502 159180
rect 392302 159128 392308 159180
rect 392360 159168 392366 159180
rect 404170 159168 404176 159180
rect 392360 159140 404176 159168
rect 392360 159128 392366 159140
rect 404170 159128 404176 159140
rect 404228 159128 404234 159180
rect 461302 159128 461308 159180
rect 461360 159168 461366 159180
rect 468018 159168 468024 159180
rect 461360 159140 468024 159168
rect 461360 159128 461366 159140
rect 468018 159128 468024 159140
rect 468076 159128 468082 159180
rect 378100 159072 383654 159100
rect 378100 159060 378106 159072
rect 395706 159060 395712 159112
rect 395764 159100 395770 159112
rect 405366 159100 405372 159112
rect 395764 159072 405372 159100
rect 395764 159060 395770 159072
rect 405366 159060 405372 159072
rect 405424 159060 405430 159112
rect 405734 159060 405740 159112
rect 405792 159100 405798 159112
rect 409230 159100 409236 159112
rect 405792 159072 409236 159100
rect 405792 159060 405798 159072
rect 409230 159060 409236 159072
rect 409288 159060 409294 159112
rect 460474 159060 460480 159112
rect 460532 159100 460538 159112
rect 466454 159100 466460 159112
rect 460532 159072 466460 159100
rect 460532 159060 460538 159072
rect 466454 159060 466460 159072
rect 466512 159060 466518 159112
rect 472250 159060 472256 159112
rect 472308 159100 472314 159112
rect 479150 159100 479156 159112
rect 472308 159072 479156 159100
rect 472308 159060 472314 159072
rect 479150 159060 479156 159072
rect 479208 159060 479214 159112
rect 378226 159032 378232 159044
rect 374840 159004 378232 159032
rect 378226 158992 378232 159004
rect 378284 158992 378290 159044
rect 447870 158992 447876 159044
rect 447928 159032 447934 159044
rect 460106 159032 460112 159044
rect 447928 159004 460112 159032
rect 447928 158992 447934 159004
rect 460106 158992 460112 159004
rect 460164 158992 460170 159044
rect 462130 158992 462136 159044
rect 462188 159032 462194 159044
rect 467926 159032 467932 159044
rect 462188 159004 467932 159032
rect 462188 158992 462194 159004
rect 467926 158992 467932 159004
rect 467984 158992 467990 159044
rect 473906 158992 473912 159044
rect 473964 159032 473970 159044
rect 480254 159032 480260 159044
rect 473964 159004 480260 159032
rect 473964 158992 473970 159004
rect 480254 158992 480260 159004
rect 480312 158992 480318 159044
rect 96246 158924 96252 158976
rect 96304 158964 96310 158976
rect 121914 158964 121920 158976
rect 96304 158936 121920 158964
rect 96304 158924 96310 158936
rect 121914 158924 121920 158936
rect 121972 158924 121978 158976
rect 124030 158924 124036 158976
rect 124088 158964 124094 158976
rect 193582 158964 193588 158976
rect 124088 158936 193588 158964
rect 124088 158924 124094 158936
rect 193582 158924 193588 158936
rect 193640 158924 193646 158976
rect 193674 158924 193680 158976
rect 193732 158964 193738 158976
rect 197354 158964 197360 158976
rect 193732 158936 197360 158964
rect 193732 158924 193738 158936
rect 197354 158924 197360 158936
rect 197412 158924 197418 158976
rect 200574 158924 200580 158976
rect 200632 158964 200638 158976
rect 224954 158964 224960 158976
rect 200632 158936 224960 158964
rect 200632 158924 200638 158936
rect 224954 158924 224960 158936
rect 225012 158924 225018 158976
rect 237558 158924 237564 158976
rect 237616 158964 237622 158976
rect 299474 158964 299480 158976
rect 237616 158936 299480 158964
rect 237616 158924 237622 158936
rect 299474 158924 299480 158936
rect 299532 158924 299538 158976
rect 314930 158924 314936 158976
rect 314988 158964 314994 158976
rect 357526 158964 357532 158976
rect 314988 158936 357532 158964
rect 314988 158924 314994 158936
rect 357526 158924 357532 158936
rect 357584 158924 357590 158976
rect 361206 158924 361212 158976
rect 361264 158964 361270 158976
rect 361264 158936 367094 158964
rect 361264 158924 361270 158936
rect 102962 158856 102968 158908
rect 103020 158896 103026 158908
rect 125502 158896 125508 158908
rect 103020 158868 125508 158896
rect 103020 158856 103026 158868
rect 125502 158856 125508 158868
rect 125560 158856 125566 158908
rect 126238 158856 126244 158908
rect 126296 158896 126302 158908
rect 129734 158896 129740 158908
rect 126296 158868 129740 158896
rect 126296 158856 126302 158868
rect 129734 158856 129740 158868
rect 129792 158856 129798 158908
rect 130746 158856 130752 158908
rect 130804 158896 130810 158908
rect 195054 158896 195060 158908
rect 130804 158868 195060 158896
rect 130804 158856 130810 158868
rect 195054 158856 195060 158868
rect 195112 158856 195118 158908
rect 195146 158856 195152 158908
rect 195204 158896 195210 158908
rect 198918 158896 198924 158908
rect 195204 158868 198924 158896
rect 195204 158856 195210 158868
rect 198918 158856 198924 158868
rect 198976 158856 198982 158908
rect 208118 158856 208124 158908
rect 208176 158896 208182 158908
rect 212442 158896 212448 158908
rect 208176 158868 212448 158896
rect 208176 158856 208182 158868
rect 212442 158856 212448 158868
rect 212500 158856 212506 158908
rect 230750 158896 230756 158908
rect 214576 158868 230756 158896
rect 109678 158788 109684 158840
rect 109736 158828 109742 158840
rect 132678 158828 132684 158840
rect 109736 158800 132684 158828
rect 109736 158788 109742 158800
rect 132678 158788 132684 158800
rect 132736 158788 132742 158840
rect 133414 158788 133420 158840
rect 133472 158828 133478 158840
rect 158714 158828 158720 158840
rect 133472 158800 158720 158828
rect 133472 158788 133478 158800
rect 158714 158788 158720 158800
rect 158772 158788 158778 158840
rect 163498 158788 163504 158840
rect 163556 158828 163562 158840
rect 195974 158828 195980 158840
rect 163556 158800 195980 158828
rect 163556 158788 163562 158800
rect 195974 158788 195980 158800
rect 196032 158788 196038 158840
rect 207290 158788 207296 158840
rect 207348 158828 207354 158840
rect 214576 158828 214604 158868
rect 230750 158856 230756 158868
rect 230808 158856 230814 158908
rect 241790 158856 241796 158908
rect 241848 158896 241854 158908
rect 303522 158896 303528 158908
rect 241848 158868 303528 158896
rect 241848 158856 241854 158868
rect 303522 158856 303528 158868
rect 303580 158856 303586 158908
rect 305638 158856 305644 158908
rect 305696 158896 305702 158908
rect 307662 158896 307668 158908
rect 305696 158868 307668 158896
rect 305696 158856 305702 158868
rect 307662 158856 307668 158868
rect 307720 158856 307726 158908
rect 310698 158856 310704 158908
rect 310756 158896 310762 158908
rect 312170 158896 312176 158908
rect 310756 158868 312176 158896
rect 310756 158856 310762 158868
rect 312170 158856 312176 158868
rect 312228 158856 312234 158908
rect 312446 158856 312452 158908
rect 312504 158896 312510 158908
rect 313366 158896 313372 158908
rect 312504 158868 313372 158896
rect 312504 158856 312510 158868
rect 313366 158856 313372 158868
rect 313424 158856 313430 158908
rect 322474 158856 322480 158908
rect 322532 158896 322538 158908
rect 365162 158896 365168 158908
rect 322532 158868 365168 158896
rect 322532 158856 322538 158868
rect 365162 158856 365168 158868
rect 365220 158856 365226 158908
rect 207348 158800 214604 158828
rect 207348 158788 207354 158800
rect 217318 158788 217324 158840
rect 217376 158828 217382 158840
rect 220354 158828 220360 158840
rect 217376 158800 220360 158828
rect 217376 158788 217382 158800
rect 220354 158788 220360 158800
rect 220412 158788 220418 158840
rect 238386 158788 238392 158840
rect 238444 158828 238450 158840
rect 242434 158828 242440 158840
rect 238444 158800 242440 158828
rect 238444 158788 238450 158800
rect 242434 158788 242440 158800
rect 242492 158788 242498 158840
rect 261110 158788 261116 158840
rect 261168 158828 261174 158840
rect 317046 158828 317052 158840
rect 261168 158800 317052 158828
rect 261168 158788 261174 158800
rect 317046 158788 317052 158800
rect 317104 158788 317110 158840
rect 319162 158788 319168 158840
rect 319220 158828 319226 158840
rect 321554 158828 321560 158840
rect 319220 158800 321560 158828
rect 319220 158788 319226 158800
rect 321554 158788 321560 158800
rect 321612 158788 321618 158840
rect 327534 158788 327540 158840
rect 327592 158828 327598 158840
rect 330478 158828 330484 158840
rect 327592 158800 330484 158828
rect 327592 158788 327598 158800
rect 330478 158788 330484 158800
rect 330536 158788 330542 158840
rect 363138 158828 363144 158840
rect 330588 158800 363144 158828
rect 90358 158720 90364 158772
rect 90416 158760 90422 158772
rect 92566 158760 92572 158772
rect 90416 158732 92572 158760
rect 90416 158720 90422 158732
rect 92566 158720 92572 158732
rect 92624 158720 92630 158772
rect 92842 158720 92848 158772
rect 92900 158760 92906 158772
rect 114462 158760 114468 158772
rect 92900 158732 114468 158760
rect 92900 158720 92906 158732
rect 114462 158720 114468 158732
rect 114520 158720 114526 158772
rect 119798 158720 119804 158772
rect 119856 158760 119862 158772
rect 147122 158760 147128 158772
rect 119856 158732 147128 158760
rect 119856 158720 119862 158732
rect 147122 158720 147128 158732
rect 147180 158720 147186 158772
rect 147582 158720 147588 158772
rect 147640 158760 147646 158772
rect 149514 158760 149520 158772
rect 147640 158732 149520 158760
rect 147640 158720 147646 158732
rect 149514 158720 149520 158732
rect 149572 158720 149578 158772
rect 153470 158720 153476 158772
rect 153528 158760 153534 158772
rect 179414 158760 179420 158772
rect 153528 158732 179420 158760
rect 153528 158720 153534 158732
rect 179414 158720 179420 158732
rect 179472 158720 179478 158772
rect 194686 158720 194692 158772
rect 194744 158760 194750 158772
rect 203702 158760 203708 158772
rect 194744 158732 203708 158760
rect 194744 158720 194750 158732
rect 203702 158720 203708 158732
rect 203760 158720 203766 158772
rect 210602 158720 210608 158772
rect 210660 158760 210666 158772
rect 215386 158760 215392 158772
rect 210660 158732 215392 158760
rect 210660 158720 210666 158732
rect 215386 158720 215392 158732
rect 215444 158720 215450 158772
rect 221550 158720 221556 158772
rect 221608 158760 221614 158772
rect 224402 158760 224408 158772
rect 221608 158732 224408 158760
rect 221608 158720 221614 158732
rect 224402 158720 224408 158732
rect 224460 158720 224466 158772
rect 240870 158720 240876 158772
rect 240928 158760 240934 158772
rect 243354 158760 243360 158772
rect 240928 158732 243360 158760
rect 240928 158720 240934 158732
rect 243354 158720 243360 158732
rect 243412 158720 243418 158772
rect 254394 158720 254400 158772
rect 254452 158760 254458 158772
rect 255406 158760 255412 158772
rect 254452 158732 255412 158760
rect 254452 158720 254458 158732
rect 255406 158720 255412 158732
rect 255464 158720 255470 158772
rect 258534 158720 258540 158772
rect 258592 158760 258598 158772
rect 260926 158760 260932 158772
rect 258592 158732 260932 158760
rect 258592 158720 258598 158732
rect 260926 158720 260932 158732
rect 260984 158720 260990 158772
rect 264422 158720 264428 158772
rect 264480 158760 264486 158772
rect 266354 158760 266360 158772
rect 264480 158732 266360 158760
rect 264480 158720 264486 158732
rect 266354 158720 266360 158732
rect 266412 158720 266418 158772
rect 267826 158720 267832 158772
rect 267884 158760 267890 158772
rect 320266 158760 320272 158772
rect 267884 158732 320272 158760
rect 267884 158720 267890 158732
rect 320266 158720 320272 158732
rect 320324 158720 320330 158772
rect 321646 158720 321652 158772
rect 321704 158760 321710 158772
rect 321704 158732 330432 158760
rect 321704 158720 321710 158732
rect 81066 158652 81072 158704
rect 81124 158692 81130 158704
rect 180886 158692 180892 158704
rect 81124 158664 180892 158692
rect 81124 158652 81130 158664
rect 180886 158652 180892 158664
rect 180944 158652 180950 158704
rect 181990 158652 181996 158704
rect 182048 158692 182054 158704
rect 256786 158692 256792 158704
rect 182048 158664 256792 158692
rect 182048 158652 182054 158664
rect 256786 158652 256792 158664
rect 256844 158652 256850 158704
rect 330404 158692 330432 158732
rect 330588 158692 330616 158800
rect 363138 158788 363144 158800
rect 363196 158788 363202 158840
rect 367066 158828 367094 158936
rect 369210 158924 369216 158976
rect 369268 158964 369274 158976
rect 384942 158964 384948 158976
rect 369268 158936 384948 158964
rect 369268 158924 369274 158936
rect 384942 158924 384948 158936
rect 385000 158924 385006 158976
rect 416682 158924 416688 158976
rect 416740 158964 416746 158976
rect 419534 158964 419540 158976
rect 416740 158936 419540 158964
rect 416740 158924 416746 158936
rect 419534 158924 419540 158936
rect 419592 158924 419598 158976
rect 456242 158924 456248 158976
rect 456300 158964 456306 158976
rect 463142 158964 463148 158976
rect 456300 158936 463148 158964
rect 456300 158924 456306 158936
rect 463142 158924 463148 158936
rect 463200 158924 463206 158976
rect 466362 158924 466368 158976
rect 466420 158964 466426 158976
rect 472618 158964 472624 158976
rect 466420 158936 472624 158964
rect 466420 158924 466426 158936
rect 472618 158924 472624 158936
rect 472676 158924 472682 158976
rect 475562 158924 475568 158976
rect 475620 158964 475626 158976
rect 481634 158964 481640 158976
rect 475620 158936 481640 158964
rect 475620 158924 475626 158936
rect 481634 158924 481640 158936
rect 481692 158924 481698 158976
rect 386138 158896 386144 158908
rect 383626 158868 386144 158896
rect 374546 158828 374552 158840
rect 367066 158800 374552 158828
rect 374546 158788 374552 158800
rect 374604 158788 374610 158840
rect 374730 158788 374736 158840
rect 374788 158828 374794 158840
rect 383626 158828 383654 158868
rect 386138 158856 386144 158868
rect 386196 158856 386202 158908
rect 391474 158856 391480 158908
rect 391532 158896 391538 158908
rect 394326 158896 394332 158908
rect 391532 158868 394332 158896
rect 391532 158856 391538 158868
rect 394326 158856 394332 158868
rect 394384 158856 394390 158908
rect 412542 158856 412548 158908
rect 412600 158896 412606 158908
rect 412910 158896 412916 158908
rect 412600 158868 412916 158896
rect 412600 158856 412606 158868
rect 412910 158856 412916 158868
rect 412968 158856 412974 158908
rect 420086 158856 420092 158908
rect 420144 158896 420150 158908
rect 423214 158896 423220 158908
rect 420144 158868 423220 158896
rect 420144 158856 420150 158868
rect 423214 158856 423220 158868
rect 423272 158856 423278 158908
rect 454586 158856 454592 158908
rect 454644 158896 454650 158908
rect 461854 158896 461860 158908
rect 454644 158868 461860 158896
rect 454644 158856 454650 158868
rect 461854 158856 461860 158868
rect 461912 158856 461918 158908
rect 465534 158856 465540 158908
rect 465592 158896 465598 158908
rect 472250 158896 472256 158908
rect 465592 158868 472256 158896
rect 465592 158856 465598 158868
rect 472250 158856 472256 158868
rect 472308 158856 472314 158908
rect 474734 158856 474740 158908
rect 474792 158896 474798 158908
rect 481358 158896 481364 158908
rect 474792 158868 481364 158896
rect 474792 158856 474798 158868
rect 481358 158856 481364 158868
rect 481416 158856 481422 158908
rect 482278 158856 482284 158908
rect 482336 158896 482342 158908
rect 487246 158896 487252 158908
rect 482336 158868 487252 158896
rect 482336 158856 482342 158868
rect 487246 158856 487252 158868
rect 487304 158856 487310 158908
rect 508314 158856 508320 158908
rect 508372 158896 508378 158908
rect 510062 158896 510068 158908
rect 508372 158868 510068 158896
rect 508372 158856 508378 158868
rect 510062 158856 510068 158868
rect 510120 158856 510126 158908
rect 374788 158800 383654 158828
rect 374788 158788 374794 158800
rect 384758 158788 384764 158840
rect 384816 158828 384822 158840
rect 389174 158828 389180 158840
rect 384816 158800 389180 158828
rect 384816 158788 384822 158800
rect 389174 158788 389180 158800
rect 389232 158788 389238 158840
rect 455414 158788 455420 158840
rect 455472 158828 455478 158840
rect 462774 158828 462780 158840
rect 455472 158800 462780 158828
rect 455472 158788 455478 158800
rect 462774 158788 462780 158800
rect 462832 158788 462838 158840
rect 464614 158788 464620 158840
rect 464672 158828 464678 158840
rect 471514 158828 471520 158840
rect 464672 158800 471520 158828
rect 464672 158788 464678 158800
rect 471514 158788 471520 158800
rect 471572 158788 471578 158840
rect 476390 158788 476396 158840
rect 476448 158828 476454 158840
rect 482646 158828 482652 158840
rect 476448 158800 482652 158828
rect 476448 158788 476454 158800
rect 482646 158788 482652 158800
rect 482704 158788 482710 158840
rect 505278 158788 505284 158840
rect 505336 158828 505342 158840
rect 507578 158828 507584 158840
rect 505336 158800 507584 158828
rect 505336 158788 505342 158800
rect 507578 158788 507584 158800
rect 507636 158788 507642 158840
rect 330662 158720 330668 158772
rect 330720 158760 330726 158772
rect 367186 158760 367192 158772
rect 330720 158732 367192 158760
rect 330720 158720 330726 158732
rect 367186 158720 367192 158732
rect 367244 158720 367250 158772
rect 367922 158720 367928 158772
rect 367980 158760 367986 158772
rect 386230 158760 386236 158772
rect 367980 158732 386236 158760
rect 367980 158720 367986 158732
rect 386230 158720 386236 158732
rect 386288 158720 386294 158772
rect 388070 158720 388076 158772
rect 388128 158760 388134 158772
rect 390370 158760 390376 158772
rect 388128 158732 390376 158760
rect 388128 158720 388134 158732
rect 390370 158720 390376 158732
rect 390428 158720 390434 158772
rect 409138 158720 409144 158772
rect 409196 158760 409202 158772
rect 410518 158760 410524 158772
rect 409196 158732 410524 158760
rect 409196 158720 409202 158732
rect 410518 158720 410524 158732
rect 410576 158720 410582 158772
rect 413370 158720 413376 158772
rect 413428 158760 413434 158772
rect 419626 158760 419632 158772
rect 413428 158732 419632 158760
rect 413428 158720 413434 158732
rect 419626 158720 419632 158732
rect 419684 158720 419690 158772
rect 452838 158720 452844 158772
rect 452896 158760 452902 158772
rect 459554 158760 459560 158772
rect 452896 158732 459560 158760
rect 452896 158720 452902 158732
rect 459554 158720 459560 158732
rect 459612 158720 459618 158772
rect 462958 158720 462964 158772
rect 463016 158760 463022 158772
rect 469214 158760 469220 158772
rect 463016 158732 469220 158760
rect 463016 158720 463022 158732
rect 469214 158720 469220 158732
rect 469272 158720 469278 158772
rect 481450 158720 481456 158772
rect 481508 158760 481514 158772
rect 486510 158760 486516 158772
rect 481508 158732 486516 158760
rect 481508 158720 481514 158732
rect 486510 158720 486516 158732
rect 486568 158720 486574 158772
rect 505738 158720 505744 158772
rect 505796 158760 505802 158772
rect 506750 158760 506756 158772
rect 505796 158732 506756 158760
rect 505796 158720 505802 158732
rect 506750 158720 506756 158732
rect 506808 158720 506814 158772
rect 507026 158720 507032 158772
rect 507084 158760 507090 158772
rect 508406 158760 508412 158772
rect 507084 158732 508412 158760
rect 507084 158720 507090 158732
rect 508406 158720 508412 158732
rect 508464 158720 508470 158772
rect 509418 158720 509424 158772
rect 509476 158760 509482 158772
rect 511718 158760 511724 158772
rect 509476 158732 511724 158760
rect 509476 158720 509482 158732
rect 511718 158720 511724 158732
rect 511776 158720 511782 158772
rect 514938 158720 514944 158772
rect 514996 158760 515002 158772
rect 518526 158760 518532 158772
rect 514996 158732 518532 158760
rect 514996 158720 515002 158732
rect 518526 158720 518532 158732
rect 518584 158720 518590 158772
rect 330404 158664 330616 158692
rect 67634 158584 67640 158636
rect 67692 158624 67698 158636
rect 170306 158624 170312 158636
rect 67692 158596 170312 158624
rect 67692 158584 67698 158596
rect 170306 158584 170312 158596
rect 170364 158584 170370 158636
rect 171962 158584 171968 158636
rect 172020 158624 172026 158636
rect 250070 158624 250076 158636
rect 172020 158596 250076 158624
rect 172020 158584 172026 158596
rect 250070 158584 250076 158596
rect 250128 158584 250134 158636
rect 74350 158516 74356 158568
rect 74408 158556 74414 158568
rect 74408 158528 173296 158556
rect 74408 158516 74414 158528
rect 71038 158448 71044 158500
rect 71096 158488 71102 158500
rect 173066 158488 173072 158500
rect 71096 158460 173072 158488
rect 71096 158448 71102 158460
rect 173066 158448 173072 158460
rect 173124 158448 173130 158500
rect 173268 158488 173296 158528
rect 175274 158516 175280 158568
rect 175332 158556 175338 158568
rect 252738 158556 252744 158568
rect 175332 158528 252744 158556
rect 175332 158516 175338 158528
rect 252738 158516 252744 158528
rect 252796 158516 252802 158568
rect 175366 158488 175372 158500
rect 173268 158460 175372 158488
rect 175366 158448 175372 158460
rect 175424 158448 175430 158500
rect 178678 158448 178684 158500
rect 178736 158488 178742 158500
rect 255590 158488 255596 158500
rect 178736 158460 255596 158488
rect 178736 158448 178742 158460
rect 255590 158448 255596 158460
rect 255648 158448 255654 158500
rect 60918 158380 60924 158432
rect 60976 158420 60982 158432
rect 164326 158420 164332 158432
rect 60976 158392 164332 158420
rect 60976 158380 60982 158392
rect 164326 158380 164332 158392
rect 164384 158380 164390 158432
rect 165246 158380 165252 158432
rect 165304 158420 165310 158432
rect 245010 158420 245016 158432
rect 165304 158392 245016 158420
rect 165304 158380 165310 158392
rect 245010 158380 245016 158392
rect 245068 158380 245074 158432
rect 64230 158312 64236 158364
rect 64288 158352 64294 158364
rect 167546 158352 167552 158364
rect 64288 158324 167552 158352
rect 64288 158312 64294 158324
rect 167546 158312 167552 158324
rect 167604 158312 167610 158364
rect 168558 158312 168564 158364
rect 168616 158352 168622 158364
rect 247126 158352 247132 158364
rect 168616 158324 247132 158352
rect 168616 158312 168622 158324
rect 247126 158312 247132 158324
rect 247184 158312 247190 158364
rect 54202 158244 54208 158296
rect 54260 158284 54266 158296
rect 160278 158284 160284 158296
rect 54260 158256 160284 158284
rect 54260 158244 54266 158256
rect 160278 158244 160284 158256
rect 160336 158244 160342 158296
rect 161842 158244 161848 158296
rect 161900 158284 161906 158296
rect 242066 158284 242072 158296
rect 161900 158256 242072 158284
rect 161900 158244 161906 158256
rect 242066 158244 242072 158256
rect 242124 158244 242130 158296
rect 47486 158176 47492 158228
rect 47544 158216 47550 158228
rect 155034 158216 155040 158228
rect 47544 158188 155040 158216
rect 47544 158176 47550 158188
rect 155034 158176 155040 158188
rect 155092 158176 155098 158228
rect 155126 158176 155132 158228
rect 155184 158216 155190 158228
rect 237374 158216 237380 158228
rect 155184 158188 237380 158216
rect 155184 158176 155190 158188
rect 237374 158176 237380 158188
rect 237432 158176 237438 158228
rect 256878 158176 256884 158228
rect 256936 158216 256942 158228
rect 315022 158216 315028 158228
rect 256936 158188 315028 158216
rect 256936 158176 256942 158188
rect 315022 158176 315028 158188
rect 315080 158176 315086 158228
rect 50798 158108 50804 158160
rect 50856 158148 50862 158160
rect 157702 158148 157708 158160
rect 50856 158120 157708 158148
rect 50856 158108 50862 158120
rect 157702 158108 157708 158120
rect 157760 158108 157766 158160
rect 158438 158108 158444 158160
rect 158496 158148 158502 158160
rect 238938 158148 238944 158160
rect 158496 158120 238944 158148
rect 158496 158108 158502 158120
rect 238938 158108 238944 158120
rect 238996 158108 239002 158160
rect 246758 158108 246764 158160
rect 246816 158148 246822 158160
rect 306926 158148 306932 158160
rect 246816 158120 306932 158148
rect 246816 158108 246822 158120
rect 306926 158108 306932 158120
rect 306984 158108 306990 158160
rect 37366 158040 37372 158092
rect 37424 158080 37430 158092
rect 146386 158080 146392 158092
rect 37424 158052 146392 158080
rect 37424 158040 37430 158052
rect 146386 158040 146392 158052
rect 146444 158040 146450 158092
rect 148410 158040 148416 158092
rect 148468 158080 148474 158092
rect 231946 158080 231952 158092
rect 148468 158052 231952 158080
rect 148468 158040 148474 158052
rect 231946 158040 231952 158052
rect 232004 158040 232010 158092
rect 243446 158040 243452 158092
rect 243504 158080 243510 158092
rect 304718 158080 304724 158092
rect 243504 158052 304724 158080
rect 243504 158040 243510 158052
rect 304718 158040 304724 158052
rect 304776 158040 304782 158092
rect 382 157972 388 158024
rect 440 158012 446 158024
rect 118878 158012 118884 158024
rect 440 157984 118884 158012
rect 440 157972 446 157984
rect 118878 157972 118884 157984
rect 118936 157972 118942 158024
rect 131574 157972 131580 158024
rect 131632 158012 131638 158024
rect 219342 158012 219348 158024
rect 131632 157984 219348 158012
rect 131632 157972 131638 157984
rect 219342 157972 219348 157984
rect 219400 157972 219406 158024
rect 236730 157972 236736 158024
rect 236788 158012 236794 158024
rect 299658 158012 299664 158024
rect 236788 157984 299664 158012
rect 236788 157972 236794 157984
rect 299658 157972 299664 157984
rect 299716 157972 299722 158024
rect 77754 157904 77760 157956
rect 77812 157944 77818 157956
rect 77812 157916 176056 157944
rect 77812 157904 77818 157916
rect 84470 157836 84476 157888
rect 84528 157876 84534 157888
rect 175918 157876 175924 157888
rect 84528 157848 175924 157876
rect 84528 157836 84534 157848
rect 175918 157836 175924 157848
rect 175976 157836 175982 157888
rect 176028 157876 176056 157916
rect 176194 157904 176200 157956
rect 176252 157944 176258 157956
rect 182266 157944 182272 157956
rect 176252 157916 182272 157944
rect 176252 157904 176258 157916
rect 182266 157904 182272 157916
rect 182324 157904 182330 157956
rect 185394 157904 185400 157956
rect 185452 157944 185458 157956
rect 260466 157944 260472 157956
rect 185452 157916 260472 157944
rect 185452 157904 185458 157916
rect 260466 157904 260472 157916
rect 260524 157904 260530 157956
rect 178034 157876 178040 157888
rect 176028 157848 178040 157876
rect 178034 157836 178040 157848
rect 178092 157836 178098 157888
rect 179414 157836 179420 157888
rect 179472 157876 179478 157888
rect 179472 157848 184888 157876
rect 179472 157836 179478 157848
rect 87782 157768 87788 157820
rect 87840 157808 87846 157820
rect 184750 157808 184756 157820
rect 87840 157780 184756 157808
rect 87840 157768 87846 157780
rect 184750 157768 184756 157780
rect 184808 157768 184814 157820
rect 184860 157808 184888 157848
rect 184934 157836 184940 157888
rect 184992 157876 184998 157888
rect 185946 157876 185952 157888
rect 184992 157848 185952 157876
rect 184992 157836 184998 157848
rect 185946 157836 185952 157848
rect 186004 157836 186010 157888
rect 188798 157836 188804 157888
rect 188856 157876 188862 157888
rect 263042 157876 263048 157888
rect 188856 157848 263048 157876
rect 188856 157836 188862 157848
rect 263042 157836 263048 157848
rect 263100 157836 263106 157888
rect 185210 157808 185216 157820
rect 184860 157780 185216 157808
rect 185210 157768 185216 157780
rect 185268 157768 185274 157820
rect 190638 157808 190644 157820
rect 185504 157780 190644 157808
rect 91186 157700 91192 157752
rect 91244 157740 91250 157752
rect 185302 157740 185308 157752
rect 91244 157712 185308 157740
rect 91244 157700 91250 157712
rect 185302 157700 185308 157712
rect 185360 157700 185366 157752
rect 94590 157632 94596 157684
rect 94648 157672 94654 157684
rect 185504 157672 185532 157780
rect 190638 157768 190644 157780
rect 190696 157768 190702 157820
rect 195514 157768 195520 157820
rect 195572 157808 195578 157820
rect 267734 157808 267740 157820
rect 195572 157780 267740 157808
rect 195572 157768 195578 157780
rect 267734 157768 267740 157780
rect 267792 157768 267798 157820
rect 185670 157700 185676 157752
rect 185728 157740 185734 157752
rect 188522 157740 188528 157752
rect 185728 157712 188528 157740
rect 185728 157700 185734 157712
rect 188522 157700 188528 157712
rect 188580 157700 188586 157752
rect 190454 157700 190460 157752
rect 190512 157740 190518 157752
rect 263686 157740 263692 157752
rect 190512 157712 263692 157740
rect 190512 157700 190518 157712
rect 263686 157700 263692 157712
rect 263744 157700 263750 157752
rect 94648 157644 185532 157672
rect 94648 157632 94654 157644
rect 185578 157632 185584 157684
rect 185636 157672 185642 157684
rect 236086 157672 236092 157684
rect 185636 157644 236092 157672
rect 185636 157632 185642 157644
rect 236086 157632 236092 157644
rect 236144 157632 236150 157684
rect 97902 157564 97908 157616
rect 97960 157604 97966 157616
rect 193306 157604 193312 157616
rect 97960 157576 193312 157604
rect 97960 157564 97966 157576
rect 193306 157564 193312 157576
rect 193364 157564 193370 157616
rect 197354 157564 197360 157616
rect 197412 157604 197418 157616
rect 251450 157604 251456 157616
rect 197412 157576 251456 157604
rect 197412 157564 197418 157576
rect 251450 157564 251456 157576
rect 251508 157564 251514 157616
rect 111334 157496 111340 157548
rect 111392 157536 111398 157548
rect 203426 157536 203432 157548
rect 111392 157508 203432 157536
rect 111392 157496 111398 157508
rect 203426 157496 203432 157508
rect 203484 157496 203490 157548
rect 204898 157496 204904 157548
rect 204956 157536 204962 157548
rect 255866 157536 255872 157548
rect 204956 157508 255872 157536
rect 204956 157496 204962 157508
rect 255866 157496 255872 157508
rect 255924 157496 255930 157548
rect 114738 157428 114744 157480
rect 114796 157468 114802 157480
rect 206554 157468 206560 157480
rect 114796 157440 206560 157468
rect 114796 157428 114802 157440
rect 206554 157428 206560 157440
rect 206612 157428 206618 157480
rect 141694 157360 141700 157412
rect 141752 157400 141758 157412
rect 227070 157400 227076 157412
rect 141752 157372 227076 157400
rect 141752 157360 141758 157372
rect 227070 157360 227076 157372
rect 227128 157360 227134 157412
rect 49142 157292 49148 157344
rect 49200 157332 49206 157344
rect 156414 157332 156420 157344
rect 49200 157304 156420 157332
rect 49200 157292 49206 157304
rect 156414 157292 156420 157304
rect 156472 157292 156478 157344
rect 158714 157292 158720 157344
rect 158772 157332 158778 157344
rect 214466 157332 214472 157344
rect 158772 157304 214472 157332
rect 158772 157292 158778 157304
rect 214466 157292 214472 157304
rect 214524 157292 214530 157344
rect 214558 157292 214564 157344
rect 214616 157332 214622 157344
rect 221366 157332 221372 157344
rect 214616 157304 221372 157332
rect 214616 157292 214622 157304
rect 221366 157292 221372 157304
rect 221424 157292 221430 157344
rect 224218 157292 224224 157344
rect 224276 157332 224282 157344
rect 281626 157332 281632 157344
rect 224276 157304 281632 157332
rect 224276 157292 224282 157304
rect 281626 157292 281632 157304
rect 281684 157292 281690 157344
rect 45738 157224 45744 157276
rect 45796 157264 45802 157276
rect 153838 157264 153844 157276
rect 45796 157236 153844 157264
rect 45796 157224 45802 157236
rect 153838 157224 153844 157236
rect 153896 157224 153902 157276
rect 163774 157224 163780 157276
rect 163832 157264 163838 157276
rect 166442 157264 166448 157276
rect 163832 157236 166448 157264
rect 163832 157224 163838 157236
rect 166442 157224 166448 157236
rect 166500 157224 166506 157276
rect 192110 157224 192116 157276
rect 192168 157264 192174 157276
rect 265158 157264 265164 157276
rect 192168 157236 265164 157264
rect 192168 157224 192174 157236
rect 265158 157224 265164 157236
rect 265216 157224 265222 157276
rect 283834 157224 283840 157276
rect 283892 157264 283898 157276
rect 335538 157264 335544 157276
rect 283892 157236 335544 157264
rect 283892 157224 283898 157236
rect 335538 157224 335544 157236
rect 335596 157224 335602 157276
rect 42426 157156 42432 157208
rect 42484 157196 42490 157208
rect 151262 157196 151268 157208
rect 42484 157168 151268 157196
rect 42484 157156 42490 157168
rect 151262 157156 151268 157168
rect 151320 157156 151326 157208
rect 156506 157156 156512 157208
rect 156564 157196 156570 157208
rect 159082 157196 159088 157208
rect 156564 157168 159088 157196
rect 156564 157156 156570 157168
rect 159082 157156 159088 157168
rect 159140 157156 159146 157208
rect 160094 157156 160100 157208
rect 160152 157196 160158 157208
rect 166166 157196 166172 157208
rect 160152 157168 166172 157196
rect 160152 157156 160158 157168
rect 166166 157156 166172 157168
rect 166224 157156 166230 157208
rect 166258 157156 166264 157208
rect 166316 157196 166322 157208
rect 171134 157196 171140 157208
rect 166316 157168 171140 157196
rect 166316 157156 166322 157168
rect 171134 157156 171140 157168
rect 171192 157156 171198 157208
rect 177022 157156 177028 157208
rect 177080 157196 177086 157208
rect 254026 157196 254032 157208
rect 177080 157168 254032 157196
rect 177080 157156 177086 157168
rect 254026 157156 254032 157168
rect 254084 157156 254090 157208
rect 290550 157156 290556 157208
rect 290608 157196 290614 157208
rect 340046 157196 340052 157208
rect 290608 157168 340052 157196
rect 290608 157156 290614 157168
rect 340046 157156 340052 157168
rect 340104 157156 340110 157208
rect 39022 157088 39028 157140
rect 39080 157128 39086 157140
rect 148778 157128 148784 157140
rect 39080 157100 148784 157128
rect 39080 157088 39086 157100
rect 148778 157088 148784 157100
rect 148836 157088 148842 157140
rect 150066 157088 150072 157140
rect 150124 157128 150130 157140
rect 233510 157128 233516 157140
rect 150124 157100 233516 157128
rect 150124 157088 150130 157100
rect 233510 157088 233516 157100
rect 233568 157088 233574 157140
rect 287146 157088 287152 157140
rect 287204 157128 287210 157140
rect 338114 157128 338120 157140
rect 287204 157100 338120 157128
rect 287204 157088 287210 157100
rect 338114 157088 338120 157100
rect 338172 157088 338178 157140
rect 35710 157020 35716 157072
rect 35768 157060 35774 157072
rect 146202 157060 146208 157072
rect 35768 157032 146208 157060
rect 35768 157020 35774 157032
rect 146202 157020 146208 157032
rect 146260 157020 146266 157072
rect 151722 157020 151728 157072
rect 151780 157060 151786 157072
rect 234798 157060 234804 157072
rect 151780 157032 234804 157060
rect 151780 157020 151786 157032
rect 234798 157020 234804 157032
rect 234856 157020 234862 157072
rect 280430 157020 280436 157072
rect 280488 157060 280494 157072
rect 333054 157060 333060 157072
rect 280488 157032 333060 157060
rect 280488 157020 280494 157032
rect 333054 157020 333060 157032
rect 333112 157020 333118 157072
rect 24762 156952 24768 157004
rect 24820 156992 24826 157004
rect 137370 156992 137376 157004
rect 24820 156964 137376 156992
rect 24820 156952 24826 156964
rect 137370 156952 137376 156964
rect 137428 156952 137434 157004
rect 138290 156952 138296 157004
rect 138348 156992 138354 157004
rect 224126 156992 224132 157004
rect 138348 156964 224132 156992
rect 138348 156952 138354 156964
rect 224126 156952 224132 156964
rect 224184 156952 224190 157004
rect 273714 156952 273720 157004
rect 273772 156992 273778 157004
rect 327902 156992 327908 157004
rect 273772 156964 327908 156992
rect 273772 156952 273778 156964
rect 327902 156952 327908 156964
rect 327960 156952 327966 157004
rect 18046 156884 18052 156936
rect 18104 156924 18110 156936
rect 132494 156924 132500 156936
rect 18104 156896 132500 156924
rect 18104 156884 18110 156896
rect 132494 156884 132500 156896
rect 132552 156884 132558 156936
rect 134886 156884 134892 156936
rect 134944 156924 134950 156936
rect 214558 156924 214564 156936
rect 134944 156896 214564 156924
rect 134944 156884 134950 156896
rect 214558 156884 214564 156896
rect 214616 156884 214622 156936
rect 224954 156884 224960 156936
rect 225012 156924 225018 156936
rect 272058 156924 272064 156936
rect 225012 156896 272064 156924
rect 225012 156884 225018 156896
rect 272058 156884 272064 156896
rect 272116 156884 272122 156936
rect 277118 156884 277124 156936
rect 277176 156924 277182 156936
rect 330478 156924 330484 156936
rect 277176 156896 330484 156924
rect 277176 156884 277182 156896
rect 330478 156884 330484 156896
rect 330536 156884 330542 156936
rect 21358 156816 21364 156868
rect 21416 156856 21422 156868
rect 135254 156856 135260 156868
rect 21416 156828 135260 156856
rect 21416 156816 21422 156828
rect 135254 156816 135260 156828
rect 135312 156816 135318 156868
rect 139118 156816 139124 156868
rect 139176 156856 139182 156868
rect 225138 156856 225144 156868
rect 139176 156828 225144 156856
rect 139176 156816 139182 156828
rect 225138 156816 225144 156828
rect 225196 156816 225202 156868
rect 226610 156816 226616 156868
rect 226668 156856 226674 156868
rect 291930 156856 291936 156868
rect 226668 156828 291936 156856
rect 226668 156816 226674 156828
rect 291930 156816 291936 156828
rect 291988 156816 291994 156868
rect 300670 156816 300676 156868
rect 300728 156856 300734 156868
rect 348050 156856 348056 156868
rect 300728 156828 348056 156856
rect 300728 156816 300734 156828
rect 348050 156816 348056 156828
rect 348108 156816 348114 156868
rect 14642 156748 14648 156800
rect 14700 156788 14706 156800
rect 130102 156788 130108 156800
rect 14700 156760 130108 156788
rect 14700 156748 14706 156760
rect 130102 156748 130108 156760
rect 130160 156748 130166 156800
rect 135806 156748 135812 156800
rect 135864 156788 135870 156800
rect 222562 156788 222568 156800
rect 135864 156760 222568 156788
rect 135864 156748 135870 156760
rect 222562 156748 222568 156760
rect 222620 156748 222626 156800
rect 230014 156748 230020 156800
rect 230072 156788 230078 156800
rect 294046 156788 294052 156800
rect 230072 156760 294052 156788
rect 230072 156748 230078 156760
rect 294046 156748 294052 156760
rect 294104 156748 294110 156800
rect 297266 156748 297272 156800
rect 297324 156788 297330 156800
rect 345106 156788 345112 156800
rect 297324 156760 345112 156788
rect 297324 156748 297330 156760
rect 345106 156748 345112 156760
rect 345164 156748 345170 156800
rect 11238 156680 11244 156732
rect 11296 156720 11302 156732
rect 127526 156720 127532 156732
rect 11296 156692 127532 156720
rect 11296 156680 11302 156692
rect 127526 156680 127532 156692
rect 127584 156680 127590 156732
rect 128170 156680 128176 156732
rect 128228 156720 128234 156732
rect 216766 156720 216772 156732
rect 128228 156692 216772 156720
rect 128228 156680 128234 156692
rect 216766 156680 216772 156692
rect 216824 156680 216830 156732
rect 223206 156680 223212 156732
rect 223264 156720 223270 156732
rect 289354 156720 289360 156732
rect 223264 156692 289360 156720
rect 223264 156680 223270 156692
rect 289354 156680 289360 156692
rect 289412 156680 289418 156732
rect 293862 156680 293868 156732
rect 293920 156720 293926 156732
rect 342530 156720 342536 156732
rect 293920 156692 342536 156720
rect 293920 156680 293926 156692
rect 342530 156680 342536 156692
rect 342588 156680 342594 156732
rect 2038 156612 2044 156664
rect 2096 156652 2102 156664
rect 120442 156652 120448 156664
rect 2096 156624 120448 156652
rect 2096 156612 2102 156624
rect 120442 156612 120448 156624
rect 120500 156612 120506 156664
rect 124858 156612 124864 156664
rect 124916 156652 124922 156664
rect 213914 156652 213920 156664
rect 124916 156624 213920 156652
rect 124916 156612 124922 156624
rect 213914 156612 213920 156624
rect 213972 156612 213978 156664
rect 216490 156612 216496 156664
rect 216548 156652 216554 156664
rect 283098 156652 283104 156664
rect 216548 156624 283104 156652
rect 216548 156612 216554 156624
rect 283098 156612 283104 156624
rect 283156 156612 283162 156664
rect 498286 156612 498292 156664
rect 498344 156652 498350 156664
rect 499298 156652 499304 156664
rect 498344 156624 499304 156652
rect 498344 156612 498350 156624
rect 499298 156612 499304 156624
rect 499356 156612 499362 156664
rect 502334 156612 502340 156664
rect 502392 156652 502398 156664
rect 503346 156652 503352 156664
rect 502392 156624 503352 156652
rect 502392 156612 502398 156624
rect 503346 156612 503352 156624
rect 503404 156612 503410 156664
rect 503714 156612 503720 156664
rect 503772 156652 503778 156664
rect 505002 156652 505008 156664
rect 503772 156624 505008 156652
rect 503772 156612 503778 156624
rect 505002 156612 505008 156624
rect 505060 156612 505066 156664
rect 52454 156544 52460 156596
rect 52512 156584 52518 156596
rect 158990 156584 158996 156596
rect 52512 156556 158996 156584
rect 52512 156544 52518 156556
rect 158990 156544 158996 156556
rect 159048 156544 159054 156596
rect 159082 156544 159088 156596
rect 159140 156584 159146 156596
rect 200758 156584 200764 156596
rect 159140 156556 200764 156584
rect 159140 156544 159146 156556
rect 200758 156544 200764 156556
rect 200816 156544 200822 156596
rect 200942 156544 200948 156596
rect 201000 156584 201006 156596
rect 270494 156584 270500 156596
rect 201000 156556 270500 156584
rect 201000 156544 201006 156556
rect 270494 156544 270500 156556
rect 270552 156544 270558 156596
rect 59262 156476 59268 156528
rect 59320 156516 59326 156528
rect 164142 156516 164148 156528
rect 59320 156488 164148 156516
rect 59320 156476 59326 156488
rect 164142 156476 164148 156488
rect 164200 156476 164206 156528
rect 166166 156476 166172 156528
rect 166224 156516 166230 156528
rect 166224 156488 166396 156516
rect 166224 156476 166230 156488
rect 69290 156408 69296 156460
rect 69348 156448 69354 156460
rect 166258 156448 166264 156460
rect 69348 156420 166264 156448
rect 69348 156408 69354 156420
rect 166258 156408 166264 156420
rect 166316 156408 166322 156460
rect 166368 156448 166396 156488
rect 166442 156476 166448 156528
rect 166500 156516 166506 156528
rect 225046 156516 225052 156528
rect 166500 156488 225052 156516
rect 166500 156476 166506 156488
rect 225046 156476 225052 156488
rect 225104 156476 225110 156528
rect 228358 156448 228364 156460
rect 166368 156420 228364 156448
rect 228358 156408 228364 156420
rect 228416 156408 228422 156460
rect 82814 156340 82820 156392
rect 82872 156380 82878 156392
rect 182082 156380 182088 156392
rect 82872 156352 182088 156380
rect 82872 156340 82878 156352
rect 182082 156340 182088 156352
rect 182140 156340 182146 156392
rect 198826 156340 198832 156392
rect 198884 156380 198890 156392
rect 200942 156380 200948 156392
rect 198884 156352 200948 156380
rect 198884 156340 198890 156352
rect 200942 156340 200948 156352
rect 201000 156340 201006 156392
rect 209774 156340 209780 156392
rect 209832 156380 209838 156392
rect 279050 156380 279056 156392
rect 209832 156352 279056 156380
rect 209832 156340 209838 156352
rect 279050 156340 279056 156352
rect 279108 156340 279114 156392
rect 99558 156272 99564 156324
rect 99616 156312 99622 156324
rect 194962 156312 194968 156324
rect 99616 156284 194968 156312
rect 99616 156272 99622 156284
rect 194962 156272 194968 156284
rect 195020 156272 195026 156324
rect 200758 156272 200764 156324
rect 200816 156312 200822 156324
rect 200816 156284 212672 156312
rect 200816 156272 200822 156284
rect 101306 156204 101312 156256
rect 101364 156244 101370 156256
rect 196250 156244 196256 156256
rect 101364 156216 196256 156244
rect 101364 156204 101370 156216
rect 196250 156204 196256 156216
rect 196308 156204 196314 156256
rect 197446 156204 197452 156256
rect 197504 156244 197510 156256
rect 211614 156244 211620 156256
rect 197504 156216 211620 156244
rect 197504 156204 197510 156216
rect 211614 156204 211620 156216
rect 211672 156204 211678 156256
rect 108022 156136 108028 156188
rect 108080 156176 108086 156188
rect 200666 156176 200672 156188
rect 108080 156148 200672 156176
rect 108080 156136 108086 156148
rect 200666 156136 200672 156148
rect 200724 156136 200730 156188
rect 201034 156176 201040 156188
rect 200776 156148 201040 156176
rect 118142 156068 118148 156120
rect 118200 156108 118206 156120
rect 200776 156108 200804 156148
rect 201034 156136 201040 156148
rect 201092 156136 201098 156188
rect 201218 156136 201224 156188
rect 201276 156176 201282 156188
rect 209130 156176 209136 156188
rect 201276 156148 209136 156176
rect 201276 156136 201282 156148
rect 209130 156136 209136 156148
rect 209188 156136 209194 156188
rect 212644 156176 212672 156284
rect 213178 156272 213184 156324
rect 213236 156312 213242 156324
rect 224218 156312 224224 156324
rect 213236 156284 224224 156312
rect 213236 156272 213242 156284
rect 224218 156272 224224 156284
rect 224276 156272 224282 156324
rect 286226 156312 286232 156324
rect 224328 156284 286232 156312
rect 214466 156204 214472 156256
rect 214524 156244 214530 156256
rect 219986 156244 219992 156256
rect 214524 156216 219992 156244
rect 214524 156204 214530 156216
rect 219986 156204 219992 156216
rect 220044 156204 220050 156256
rect 220078 156204 220084 156256
rect 220136 156244 220142 156256
rect 224328 156244 224356 156284
rect 286226 156272 286232 156284
rect 286284 156272 286290 156324
rect 266906 156244 266912 156256
rect 220136 156216 224356 156244
rect 229066 156216 266912 156244
rect 220136 156204 220142 156216
rect 215478 156176 215484 156188
rect 212644 156148 215484 156176
rect 215478 156136 215484 156148
rect 215536 156136 215542 156188
rect 218054 156136 218060 156188
rect 218112 156176 218118 156188
rect 229066 156176 229094 156216
rect 266906 156204 266912 156216
rect 266964 156204 266970 156256
rect 218112 156148 229094 156176
rect 218112 156136 218118 156148
rect 230750 156136 230756 156188
rect 230808 156176 230814 156188
rect 277118 156176 277124 156188
rect 230808 156148 277124 156176
rect 230808 156136 230814 156148
rect 277118 156136 277124 156148
rect 277176 156136 277182 156188
rect 118200 156080 200804 156108
rect 118200 156068 118206 156080
rect 203058 156068 203064 156120
rect 203116 156108 203122 156120
rect 273898 156108 273904 156120
rect 203116 156080 273904 156108
rect 203116 156068 203122 156080
rect 273898 156068 273904 156080
rect 273956 156068 273962 156120
rect 121454 156000 121460 156052
rect 121512 156040 121518 156052
rect 197446 156040 197452 156052
rect 121512 156012 197452 156040
rect 121512 156000 121518 156012
rect 197446 156000 197452 156012
rect 197504 156000 197510 156052
rect 200942 156000 200948 156052
rect 201000 156040 201006 156052
rect 201402 156040 201408 156052
rect 201000 156012 201408 156040
rect 201000 156000 201006 156012
rect 201402 156000 201408 156012
rect 201460 156000 201466 156052
rect 202230 156000 202236 156052
rect 202288 156040 202294 156052
rect 273254 156040 273260 156052
rect 202288 156012 273260 156040
rect 202288 156000 202294 156012
rect 273254 156000 273260 156012
rect 273312 156000 273318 156052
rect 145006 155932 145012 155984
rect 145064 155972 145070 155984
rect 229646 155972 229652 155984
rect 145064 155944 229652 155972
rect 145064 155932 145070 155944
rect 229646 155932 229652 155944
rect 229704 155932 229710 155984
rect 66806 155864 66812 155916
rect 66864 155904 66870 155916
rect 82906 155904 82912 155916
rect 66864 155876 82912 155904
rect 66864 155864 66870 155876
rect 82906 155864 82912 155876
rect 82964 155864 82970 155916
rect 88702 155864 88708 155916
rect 88760 155904 88766 155916
rect 186406 155904 186412 155916
rect 88760 155876 186412 155904
rect 88760 155864 88766 155876
rect 186406 155864 186412 155876
rect 186464 155864 186470 155916
rect 189166 155904 189172 155916
rect 186700 155876 189172 155904
rect 60090 155796 60096 155848
rect 60148 155836 60154 155848
rect 79318 155836 79324 155848
rect 60148 155808 79324 155836
rect 60148 155796 60154 155808
rect 79318 155796 79324 155808
rect 79376 155796 79382 155848
rect 92014 155796 92020 155848
rect 92072 155836 92078 155848
rect 186700 155836 186728 155876
rect 189166 155864 189172 155876
rect 189224 155864 189230 155916
rect 194318 155904 194324 155916
rect 192864 155876 194324 155904
rect 92072 155808 186728 155836
rect 92072 155796 92078 155808
rect 186774 155796 186780 155848
rect 186832 155836 186838 155848
rect 192864 155836 192892 155876
rect 194318 155864 194324 155876
rect 194376 155864 194382 155916
rect 196342 155864 196348 155916
rect 196400 155904 196406 155916
rect 268838 155904 268844 155916
rect 196400 155876 268844 155904
rect 196400 155864 196406 155876
rect 268838 155864 268844 155876
rect 268896 155864 268902 155916
rect 296438 155864 296444 155916
rect 296496 155904 296502 155916
rect 345198 155904 345204 155916
rect 296496 155876 345204 155904
rect 296496 155864 296502 155876
rect 345198 155864 345204 155876
rect 345256 155864 345262 155916
rect 186832 155808 192892 155836
rect 186832 155796 186838 155808
rect 192938 155796 192944 155848
rect 192996 155836 193002 155848
rect 266262 155836 266268 155848
rect 192996 155808 266268 155836
rect 192996 155796 193002 155808
rect 266262 155796 266268 155808
rect 266320 155796 266326 155848
rect 293034 155796 293040 155848
rect 293092 155836 293098 155848
rect 342346 155836 342352 155848
rect 293092 155808 342352 155836
rect 293092 155796 293098 155808
rect 342346 155796 342352 155808
rect 342404 155796 342410 155848
rect 12158 155728 12164 155780
rect 12216 155768 12222 155780
rect 110322 155768 110328 155780
rect 12216 155740 110328 155768
rect 12216 155728 12222 155740
rect 110322 155728 110328 155740
rect 110380 155728 110386 155780
rect 112254 155728 112260 155780
rect 112312 155768 112318 155780
rect 204622 155768 204628 155780
rect 112312 155740 204628 155768
rect 112312 155728 112318 155740
rect 204622 155728 204628 155740
rect 204680 155728 204686 155780
rect 206462 155728 206468 155780
rect 206520 155768 206526 155780
rect 276106 155768 276112 155780
rect 206520 155740 276112 155768
rect 206520 155728 206526 155740
rect 276106 155728 276112 155740
rect 276164 155728 276170 155780
rect 289722 155728 289728 155780
rect 289780 155768 289786 155780
rect 339586 155768 339592 155780
rect 289780 155740 339592 155768
rect 289780 155728 289786 155740
rect 339586 155728 339592 155740
rect 339644 155728 339650 155780
rect 46566 155660 46572 155712
rect 46624 155700 46630 155712
rect 75086 155700 75092 155712
rect 46624 155672 75092 155700
rect 46624 155660 46630 155672
rect 75086 155660 75092 155672
rect 75144 155660 75150 155712
rect 81894 155660 81900 155712
rect 81952 155700 81958 155712
rect 180978 155700 180984 155712
rect 81952 155672 180984 155700
rect 81952 155660 81958 155672
rect 180978 155660 180984 155672
rect 181036 155660 181042 155712
rect 186222 155660 186228 155712
rect 186280 155700 186286 155712
rect 260834 155700 260840 155712
rect 186280 155672 260840 155700
rect 186280 155660 186286 155672
rect 260834 155660 260840 155672
rect 260892 155660 260898 155712
rect 270310 155660 270316 155712
rect 270368 155700 270374 155712
rect 325326 155700 325332 155712
rect 270368 155672 325332 155700
rect 270368 155660 270374 155672
rect 325326 155660 325332 155672
rect 325384 155660 325390 155712
rect 344370 155660 344376 155712
rect 344428 155700 344434 155712
rect 381814 155700 381820 155712
rect 344428 155672 381820 155700
rect 344428 155660 344434 155672
rect 381814 155660 381820 155672
rect 381872 155660 381878 155712
rect 53374 155592 53380 155644
rect 53432 155632 53438 155644
rect 66622 155632 66628 155644
rect 53432 155604 66628 155632
rect 53432 155592 53438 155604
rect 66622 155592 66628 155604
rect 66680 155592 66686 155644
rect 71866 155592 71872 155644
rect 71924 155632 71930 155644
rect 172698 155632 172704 155644
rect 71924 155604 172704 155632
rect 71924 155592 71930 155604
rect 172698 155592 172704 155604
rect 172756 155592 172762 155644
rect 176286 155592 176292 155644
rect 176344 155632 176350 155644
rect 253382 155632 253388 155644
rect 176344 155604 253388 155632
rect 176344 155592 176350 155604
rect 253382 155592 253388 155604
rect 253440 155592 253446 155644
rect 266998 155592 267004 155644
rect 267056 155632 267062 155644
rect 322106 155632 322112 155644
rect 267056 155604 322112 155632
rect 267056 155592 267062 155604
rect 322106 155592 322112 155604
rect 322164 155592 322170 155644
rect 340966 155592 340972 155644
rect 341024 155632 341030 155644
rect 378134 155632 378140 155644
rect 341024 155604 378140 155632
rect 341024 155592 341030 155604
rect 378134 155592 378140 155604
rect 378192 155592 378198 155644
rect 39850 155524 39856 155576
rect 39908 155564 39914 155576
rect 68922 155564 68928 155576
rect 39908 155536 68928 155564
rect 39908 155524 39914 155536
rect 68922 155524 68928 155536
rect 68980 155524 68986 155576
rect 75178 155524 75184 155576
rect 75236 155564 75242 155576
rect 176378 155564 176384 155576
rect 75236 155536 176384 155564
rect 75236 155524 75242 155536
rect 176378 155524 176384 155536
rect 176436 155524 176442 155576
rect 179506 155524 179512 155576
rect 179564 155564 179570 155576
rect 255682 155564 255688 155576
rect 179564 155536 255688 155564
rect 179564 155524 179570 155536
rect 255682 155524 255688 155536
rect 255740 155524 255746 155576
rect 263594 155524 263600 155576
rect 263652 155564 263658 155576
rect 320174 155564 320180 155576
rect 263652 155536 320180 155564
rect 263652 155524 263658 155536
rect 320174 155524 320180 155536
rect 320232 155524 320238 155576
rect 337654 155524 337660 155576
rect 337712 155564 337718 155576
rect 375558 155564 375564 155576
rect 337712 155536 375564 155564
rect 337712 155524 337718 155536
rect 375558 155524 375564 155536
rect 375616 155524 375622 155576
rect 65150 155456 65156 155508
rect 65208 155496 65214 155508
rect 168650 155496 168656 155508
rect 65208 155468 168656 155496
rect 65208 155456 65214 155468
rect 168650 155456 168656 155468
rect 168708 155456 168714 155508
rect 169386 155456 169392 155508
rect 169444 155496 169450 155508
rect 248230 155496 248236 155508
rect 169444 155468 248236 155496
rect 169444 155456 169450 155468
rect 248230 155456 248236 155468
rect 248288 155456 248294 155508
rect 260282 155456 260288 155508
rect 260340 155496 260346 155508
rect 317598 155496 317604 155508
rect 260340 155468 317604 155496
rect 260340 155456 260346 155468
rect 317598 155456 317604 155468
rect 317656 155456 317662 155508
rect 333422 155456 333428 155508
rect 333480 155496 333486 155508
rect 373442 155496 373448 155508
rect 333480 155468 373448 155496
rect 333480 155456 333486 155468
rect 373442 155456 373448 155468
rect 373500 155456 373506 155508
rect 7926 155388 7932 155440
rect 7984 155428 7990 155440
rect 124674 155428 124680 155440
rect 7984 155400 124680 155428
rect 7984 155388 7990 155400
rect 124674 155388 124680 155400
rect 124732 155388 124738 155440
rect 149238 155388 149244 155440
rect 149296 155428 149302 155440
rect 232866 155428 232872 155440
rect 149296 155400 232872 155428
rect 149296 155388 149302 155400
rect 232866 155388 232872 155400
rect 232924 155388 232930 155440
rect 253566 155388 253572 155440
rect 253624 155428 253630 155440
rect 312446 155428 312452 155440
rect 253624 155400 312452 155428
rect 253624 155388 253630 155400
rect 312446 155388 312452 155400
rect 312504 155388 312510 155440
rect 330110 155388 330116 155440
rect 330168 155428 330174 155440
rect 370866 155428 370872 155440
rect 330168 155400 370872 155428
rect 330168 155388 330174 155400
rect 370866 155388 370872 155400
rect 370924 155388 370930 155440
rect 8754 155320 8760 155372
rect 8812 155360 8818 155372
rect 125686 155360 125692 155372
rect 8812 155332 125692 155360
rect 8812 155320 8818 155332
rect 125686 155320 125692 155332
rect 125744 155320 125750 155372
rect 145834 155320 145840 155372
rect 145892 155360 145898 155372
rect 229186 155360 229192 155372
rect 145892 155332 229192 155360
rect 145892 155320 145898 155332
rect 229186 155320 229192 155332
rect 229244 155320 229250 155372
rect 250162 155320 250168 155372
rect 250220 155360 250226 155372
rect 309870 155360 309876 155372
rect 250220 155332 309876 155360
rect 250220 155320 250226 155332
rect 309870 155320 309876 155332
rect 309928 155320 309934 155372
rect 319990 155320 319996 155372
rect 320048 155360 320054 155372
rect 363230 155360 363236 155372
rect 320048 155332 363236 155360
rect 320048 155320 320054 155332
rect 363230 155320 363236 155332
rect 363288 155320 363294 155372
rect 4522 155252 4528 155304
rect 4580 155292 4586 155304
rect 122006 155292 122012 155304
rect 4580 155264 122012 155292
rect 4580 155252 4586 155264
rect 122006 155252 122012 155264
rect 122064 155252 122070 155304
rect 142522 155252 142528 155304
rect 142580 155292 142586 155304
rect 227806 155292 227812 155304
rect 142580 155264 227812 155292
rect 142580 155252 142586 155264
rect 227806 155252 227812 155264
rect 227864 155252 227870 155304
rect 233326 155252 233332 155304
rect 233384 155292 233390 155304
rect 297082 155292 297088 155304
rect 233384 155264 297088 155292
rect 233384 155252 233390 155264
rect 297082 155252 297088 155264
rect 297140 155252 297146 155304
rect 299750 155252 299756 155304
rect 299808 155292 299814 155304
rect 347866 155292 347872 155304
rect 299808 155264 347872 155292
rect 299808 155252 299814 155264
rect 347866 155252 347872 155264
rect 347924 155252 347930 155304
rect 373810 155252 373816 155304
rect 373868 155292 373874 155304
rect 404078 155292 404084 155304
rect 373868 155264 404084 155292
rect 373868 155252 373874 155264
rect 404078 155252 404084 155264
rect 404136 155252 404142 155304
rect 5350 155184 5356 155236
rect 5408 155224 5414 155236
rect 123018 155224 123024 155236
rect 5408 155196 123024 155224
rect 5408 155184 5414 155196
rect 123018 155184 123024 155196
rect 123076 155184 123082 155236
rect 128998 155184 129004 155236
rect 129056 155224 129062 155236
rect 217410 155224 217416 155236
rect 129056 155196 217416 155224
rect 129056 155184 129062 155196
rect 217410 155184 217416 155196
rect 217468 155184 217474 155236
rect 240042 155184 240048 155236
rect 240100 155224 240106 155236
rect 302510 155224 302516 155236
rect 240100 155196 302516 155224
rect 240100 155184 240106 155196
rect 302510 155184 302516 155196
rect 302568 155184 302574 155236
rect 306558 155184 306564 155236
rect 306616 155224 306622 155236
rect 352466 155224 352472 155236
rect 306616 155196 352472 155224
rect 306616 155184 306622 155196
rect 352466 155184 352472 155196
rect 352524 155184 352530 155236
rect 370406 155184 370412 155236
rect 370464 155224 370470 155236
rect 401686 155224 401692 155236
rect 370464 155196 401692 155224
rect 370464 155184 370470 155196
rect 401686 155184 401692 155196
rect 401744 155184 401750 155236
rect 89530 155116 89536 155168
rect 89588 155156 89594 155168
rect 187234 155156 187240 155168
rect 89588 155128 187240 155156
rect 89588 155116 89594 155128
rect 187234 155116 187240 155128
rect 187292 155116 187298 155168
rect 189626 155116 189632 155168
rect 189684 155156 189690 155168
rect 263686 155156 263692 155168
rect 189684 155128 263692 155156
rect 189684 155116 189690 155128
rect 263686 155116 263692 155128
rect 263744 155116 263750 155168
rect 98730 155048 98736 155100
rect 98788 155088 98794 155100
rect 186498 155088 186504 155100
rect 98788 155060 186504 155088
rect 98788 155048 98794 155060
rect 186498 155048 186504 155060
rect 186556 155048 186562 155100
rect 186866 155048 186872 155100
rect 186924 155088 186930 155100
rect 191190 155088 191196 155100
rect 186924 155060 191196 155088
rect 186924 155048 186930 155060
rect 191190 155048 191196 155060
rect 191248 155048 191254 155100
rect 195974 155048 195980 155100
rect 196032 155088 196038 155100
rect 196986 155088 196992 155100
rect 196032 155060 196992 155088
rect 196032 155048 196038 155060
rect 196986 155048 196992 155060
rect 197044 155048 197050 155100
rect 199654 155048 199660 155100
rect 199712 155088 199718 155100
rect 271414 155088 271420 155100
rect 199712 155060 271420 155088
rect 199712 155048 199718 155060
rect 271414 155048 271420 155060
rect 271472 155048 271478 155100
rect 303154 155048 303160 155100
rect 303212 155088 303218 155100
rect 350350 155088 350356 155100
rect 303212 155060 350356 155088
rect 303212 155048 303218 155060
rect 350350 155048 350356 155060
rect 350408 155048 350414 155100
rect 95418 154980 95424 155032
rect 95476 155020 95482 155032
rect 190822 155020 190828 155032
rect 95476 154992 190828 155020
rect 95476 154980 95482 154992
rect 190822 154980 190828 154992
rect 190880 154980 190886 155032
rect 190914 154980 190920 155032
rect 190972 155020 190978 155032
rect 200114 155020 200120 155032
rect 190972 154992 200120 155020
rect 190972 154980 190978 154992
rect 200114 154980 200120 154992
rect 200172 154980 200178 155032
rect 207014 154980 207020 155032
rect 207072 155020 207078 155032
rect 269482 155020 269488 155032
rect 207072 154992 269488 155020
rect 207072 154980 207078 154992
rect 269482 154980 269488 154992
rect 269540 154980 269546 155032
rect 15470 154912 15476 154964
rect 15528 154952 15534 154964
rect 109034 154952 109040 154964
rect 15528 154924 109040 154952
rect 15528 154912 15534 154924
rect 109034 154912 109040 154924
rect 109092 154912 109098 154964
rect 122282 154912 122288 154964
rect 122340 154952 122346 154964
rect 190730 154952 190736 154964
rect 122340 154924 190736 154952
rect 122340 154912 122346 154924
rect 190730 154912 190736 154924
rect 190788 154912 190794 154964
rect 191006 154912 191012 154964
rect 191064 154952 191070 154964
rect 211246 154952 211252 154964
rect 191064 154924 211252 154952
rect 191064 154912 191070 154924
rect 211246 154912 211252 154924
rect 211304 154912 211310 154964
rect 214650 154912 214656 154964
rect 214708 154952 214714 154964
rect 261386 154952 261392 154964
rect 214708 154924 261392 154952
rect 214708 154912 214714 154924
rect 261386 154912 261392 154924
rect 261444 154912 261450 154964
rect 106366 154844 106372 154896
rect 106424 154884 106430 154896
rect 190914 154884 190920 154896
rect 106424 154856 190920 154884
rect 106424 154844 106430 154856
rect 190914 154844 190920 154856
rect 190972 154844 190978 154896
rect 191190 154844 191196 154896
rect 191248 154884 191254 154896
rect 245838 154884 245844 154896
rect 191248 154856 245844 154884
rect 191248 154844 191254 154856
rect 245838 154844 245844 154856
rect 245896 154844 245902 154896
rect 125778 154776 125784 154828
rect 125836 154816 125842 154828
rect 214834 154816 214840 154828
rect 125836 154788 214840 154816
rect 125836 154776 125842 154788
rect 214834 154776 214840 154788
rect 214892 154776 214898 154828
rect 110506 154708 110512 154760
rect 110564 154748 110570 154760
rect 139302 154748 139308 154760
rect 110564 154720 139308 154748
rect 110564 154708 110570 154720
rect 139302 154708 139308 154720
rect 139360 154708 139366 154760
rect 151814 154708 151820 154760
rect 151872 154748 151878 154760
rect 153102 154748 153108 154760
rect 151872 154720 153108 154748
rect 151872 154708 151878 154720
rect 153102 154708 153108 154720
rect 153160 154708 153166 154760
rect 155954 154708 155960 154760
rect 156012 154748 156018 154760
rect 238018 154748 238024 154760
rect 156012 154720 238024 154748
rect 156012 154708 156018 154720
rect 238018 154708 238024 154720
rect 238076 154708 238082 154760
rect 280264 154720 283788 154748
rect 109126 154640 109132 154692
rect 109184 154680 109190 154692
rect 133046 154680 133052 154692
rect 109184 154652 133052 154680
rect 109184 154640 109190 154652
rect 133046 154640 133052 154652
rect 133104 154640 133110 154692
rect 157334 154680 157340 154692
rect 142080 154652 142844 154680
rect 118602 154572 118608 154624
rect 118660 154612 118666 154624
rect 119982 154612 119988 154624
rect 118660 154584 119988 154612
rect 118660 154572 118666 154584
rect 119982 154572 119988 154584
rect 120040 154572 120046 154624
rect 137094 154572 137100 154624
rect 137152 154612 137158 154624
rect 138014 154612 138020 154624
rect 137152 154584 138020 154612
rect 137152 154572 137158 154584
rect 138014 154572 138020 154584
rect 138072 154572 138078 154624
rect 51074 154504 51080 154556
rect 51132 154544 51138 154556
rect 142080 154544 142108 154652
rect 142154 154572 142160 154624
rect 142212 154612 142218 154624
rect 142212 154584 142752 154612
rect 142212 154572 142218 154584
rect 51132 154516 142108 154544
rect 51132 154504 51138 154516
rect 44174 154436 44180 154488
rect 44232 154476 44238 154488
rect 142338 154476 142344 154488
rect 44232 154448 142344 154476
rect 44232 154436 44238 154448
rect 142338 154436 142344 154448
rect 142396 154436 142402 154488
rect 142430 154436 142436 154488
rect 142488 154436 142494 154488
rect 142724 154476 142752 154584
rect 142816 154544 142844 154652
rect 157306 154640 157340 154680
rect 157392 154640 157398 154692
rect 162670 154640 162676 154692
rect 162728 154680 162734 154692
rect 243078 154680 243084 154692
rect 162728 154652 243084 154680
rect 162728 154640 162734 154652
rect 243078 154640 243084 154652
rect 243136 154640 243142 154692
rect 157306 154612 157334 154640
rect 157168 154584 157334 154612
rect 157168 154544 157196 154584
rect 159358 154572 159364 154624
rect 159416 154612 159422 154624
rect 240594 154612 240600 154624
rect 159416 154584 240600 154612
rect 159416 154572 159422 154584
rect 240594 154572 240600 154584
rect 240652 154572 240658 154624
rect 142816 154516 157196 154544
rect 157242 154504 157248 154556
rect 157300 154544 157306 154556
rect 212902 154544 212908 154556
rect 157300 154516 212908 154544
rect 157300 154504 157306 154516
rect 212902 154504 212908 154516
rect 212960 154504 212966 154556
rect 218330 154504 218336 154556
rect 218388 154544 218394 154556
rect 280264 154544 280292 154720
rect 283650 154544 283656 154556
rect 218388 154516 280292 154544
rect 283024 154516 283656 154544
rect 218388 154504 218394 154516
rect 190914 154476 190920 154488
rect 142724 154448 190920 154476
rect 190914 154436 190920 154448
rect 190972 154436 190978 154488
rect 191006 154436 191012 154488
rect 191064 154476 191070 154488
rect 201218 154476 201224 154488
rect 191064 154448 201224 154476
rect 191064 154436 191070 154448
rect 201218 154436 201224 154448
rect 201276 154436 201282 154488
rect 201310 154436 201316 154488
rect 201368 154476 201374 154488
rect 207934 154476 207940 154488
rect 201368 154448 207940 154476
rect 201368 154436 201374 154448
rect 207934 154436 207940 154448
rect 207992 154436 207998 154488
rect 215294 154436 215300 154488
rect 215352 154476 215358 154488
rect 283024 154476 283052 154516
rect 283650 154504 283656 154516
rect 283708 154504 283714 154556
rect 283760 154544 283788 154720
rect 285582 154544 285588 154556
rect 283760 154516 285588 154544
rect 285582 154504 285588 154516
rect 285640 154504 285646 154556
rect 285674 154504 285680 154556
rect 285732 154544 285738 154556
rect 337470 154544 337476 154556
rect 285732 154516 337476 154544
rect 285732 154504 285738 154516
rect 337470 154504 337476 154516
rect 337528 154504 337534 154556
rect 353662 154504 353668 154556
rect 353720 154544 353726 154556
rect 388898 154544 388904 154556
rect 353720 154516 388904 154544
rect 353720 154504 353726 154516
rect 388898 154504 388904 154516
rect 388956 154504 388962 154556
rect 215352 154448 283052 154476
rect 215352 154436 215358 154448
rect 283282 154436 283288 154488
rect 283340 154476 283346 154488
rect 334894 154476 334900 154488
rect 283340 154448 334900 154476
rect 283340 154436 283346 154448
rect 334894 154436 334900 154448
rect 334952 154436 334958 154488
rect 349522 154436 349528 154488
rect 349580 154476 349586 154488
rect 386322 154476 386328 154488
rect 349580 154448 386328 154476
rect 349580 154436 349586 154448
rect 386322 154436 386328 154448
rect 386380 154436 386386 154488
rect 390646 154436 390652 154488
rect 390704 154476 390710 154488
rect 417142 154476 417148 154488
rect 390704 154448 417148 154476
rect 390704 154436 390710 154448
rect 417142 154436 417148 154448
rect 417200 154436 417206 154488
rect 114462 154368 114468 154420
rect 114520 154408 114526 154420
rect 118602 154408 118608 154420
rect 114520 154380 118608 154408
rect 114520 154368 114526 154380
rect 118602 154368 118608 154380
rect 118660 154368 118666 154420
rect 118694 154368 118700 154420
rect 118752 154408 118758 154420
rect 119890 154408 119896 154420
rect 118752 154380 119896 154408
rect 118752 154368 118758 154380
rect 119890 154368 119896 154380
rect 119948 154368 119954 154420
rect 119982 154368 119988 154420
rect 120040 154408 120046 154420
rect 142448 154408 142476 154436
rect 120040 154380 142476 154408
rect 120040 154368 120046 154380
rect 142614 154368 142620 154420
rect 142672 154408 142678 154420
rect 189810 154408 189816 154420
rect 142672 154380 189816 154408
rect 142672 154368 142678 154380
rect 189810 154368 189816 154380
rect 189868 154368 189874 154420
rect 191190 154368 191196 154420
rect 191248 154408 191254 154420
rect 202046 154408 202052 154420
rect 191248 154380 202052 154408
rect 191248 154368 191254 154380
rect 202046 154368 202052 154380
rect 202104 154368 202110 154420
rect 204990 154368 204996 154420
rect 205048 154408 205054 154420
rect 275830 154408 275836 154420
rect 205048 154380 275836 154408
rect 205048 154368 205054 154380
rect 275830 154368 275836 154380
rect 275888 154368 275894 154420
rect 276198 154368 276204 154420
rect 276256 154408 276262 154420
rect 329926 154408 329932 154420
rect 276256 154380 329932 154408
rect 276256 154368 276262 154380
rect 329926 154368 329932 154380
rect 329984 154368 329990 154420
rect 346394 154368 346400 154420
rect 346452 154408 346458 154420
rect 383746 154408 383752 154420
rect 346452 154380 383752 154408
rect 346452 154368 346458 154380
rect 383746 154368 383752 154380
rect 383804 154368 383810 154420
rect 397362 154368 397368 154420
rect 397420 154408 397426 154420
rect 422386 154408 422392 154420
rect 397420 154380 422392 154408
rect 397420 154368 397426 154380
rect 422386 154368 422392 154380
rect 422444 154368 422450 154420
rect 34514 154300 34520 154352
rect 34572 154340 34578 154352
rect 34572 154312 142660 154340
rect 34572 154300 34578 154312
rect 142632 154284 142660 154312
rect 142706 154300 142712 154352
rect 142764 154340 142770 154352
rect 201126 154340 201132 154352
rect 142764 154312 201132 154340
rect 142764 154300 142770 154312
rect 201126 154300 201132 154312
rect 201184 154300 201190 154352
rect 201218 154300 201224 154352
rect 201276 154340 201282 154352
rect 202690 154340 202696 154352
rect 201276 154312 202696 154340
rect 201276 154300 201282 154312
rect 202690 154300 202696 154312
rect 202748 154300 202754 154352
rect 208394 154300 208400 154352
rect 208452 154340 208458 154352
rect 278406 154340 278412 154352
rect 208452 154312 278412 154340
rect 208452 154300 208458 154312
rect 278406 154300 278412 154312
rect 278464 154300 278470 154352
rect 278866 154300 278872 154352
rect 278924 154340 278930 154352
rect 332410 154340 332416 154352
rect 278924 154312 332416 154340
rect 278924 154300 278930 154312
rect 332410 154300 332416 154312
rect 332468 154300 332474 154352
rect 343542 154300 343548 154352
rect 343600 154340 343606 154352
rect 381170 154340 381176 154352
rect 343600 154312 381176 154340
rect 343600 154300 343606 154312
rect 381170 154300 381176 154312
rect 381228 154300 381234 154352
rect 393314 154300 393320 154352
rect 393372 154340 393378 154352
rect 419718 154340 419724 154352
rect 393372 154312 419724 154340
rect 393372 154300 393378 154312
rect 419718 154300 419724 154312
rect 419776 154300 419782 154352
rect 37918 154232 37924 154284
rect 37976 154272 37982 154284
rect 37976 154244 142292 154272
rect 37976 154232 37982 154244
rect 27246 154164 27252 154216
rect 27304 154204 27310 154216
rect 136910 154204 136916 154216
rect 27304 154176 136916 154204
rect 27304 154164 27310 154176
rect 136910 154164 136916 154176
rect 136968 154164 136974 154216
rect 142154 154204 142160 154216
rect 137112 154176 142160 154204
rect 23474 154096 23480 154148
rect 23532 154136 23538 154148
rect 137002 154136 137008 154148
rect 23532 154108 137008 154136
rect 23532 154096 23538 154108
rect 137002 154096 137008 154108
rect 137060 154096 137066 154148
rect 13814 154028 13820 154080
rect 13872 154068 13878 154080
rect 129274 154068 129280 154080
rect 13872 154040 129280 154068
rect 13872 154028 13878 154040
rect 129274 154028 129280 154040
rect 129332 154028 129338 154080
rect 137112 154068 137140 154176
rect 142154 154164 142160 154176
rect 142212 154164 142218 154216
rect 142264 154204 142292 154244
rect 142614 154232 142620 154284
rect 142672 154232 142678 154284
rect 142890 154232 142896 154284
rect 142948 154272 142954 154284
rect 150618 154272 150624 154284
rect 142948 154244 150624 154272
rect 142948 154232 142954 154244
rect 150618 154232 150624 154244
rect 150676 154232 150682 154284
rect 152366 154232 152372 154284
rect 152424 154272 152430 154284
rect 163498 154272 163504 154284
rect 152424 154244 163504 154272
rect 152424 154232 152430 154244
rect 163498 154232 163504 154244
rect 163556 154232 163562 154284
rect 176654 154232 176660 154284
rect 176712 154272 176718 154284
rect 179690 154272 179696 154284
rect 176712 154244 179696 154272
rect 176712 154232 176718 154244
rect 179690 154232 179696 154244
rect 179748 154232 179754 154284
rect 182174 154232 182180 154284
rect 182232 154272 182238 154284
rect 258534 154272 258540 154284
rect 182232 154244 258540 154272
rect 182232 154232 182238 154244
rect 258534 154232 258540 154244
rect 258592 154232 258598 154284
rect 262214 154232 262220 154284
rect 262272 154272 262278 154284
rect 319530 154272 319536 154284
rect 262272 154244 319536 154272
rect 262272 154232 262278 154244
rect 319530 154232 319536 154244
rect 319588 154232 319594 154284
rect 339494 154232 339500 154284
rect 339552 154272 339558 154284
rect 378594 154272 378600 154284
rect 339552 154244 378600 154272
rect 339552 154232 339558 154244
rect 378594 154232 378600 154244
rect 378652 154232 378658 154284
rect 386506 154232 386512 154284
rect 386564 154272 386570 154284
rect 414566 154272 414572 154284
rect 386564 154244 414572 154272
rect 386564 154232 386570 154244
rect 414566 154232 414572 154244
rect 414624 154232 414630 154284
rect 147582 154204 147588 154216
rect 142264 154176 147588 154204
rect 147582 154164 147588 154176
rect 147640 154164 147646 154216
rect 147766 154164 147772 154216
rect 147824 154204 147830 154216
rect 157242 154204 157248 154216
rect 147824 154176 157248 154204
rect 147824 154164 147830 154176
rect 157242 154164 157248 154176
rect 157300 154164 157306 154216
rect 157334 154164 157340 154216
rect 157392 154204 157398 154216
rect 158346 154204 158352 154216
rect 157392 154176 158352 154204
rect 157392 154164 157398 154176
rect 158346 154164 158352 154176
rect 158404 154164 158410 154216
rect 161474 154164 161480 154216
rect 161532 154204 161538 154216
rect 166074 154204 166080 154216
rect 161532 154176 166080 154204
rect 161532 154164 161538 154176
rect 166074 154164 166080 154176
rect 166132 154164 166138 154216
rect 172514 154164 172520 154216
rect 172572 154204 172578 154216
rect 250806 154204 250812 154216
rect 172572 154176 250812 154204
rect 172572 154164 172578 154176
rect 250806 154164 250812 154176
rect 250864 154164 250870 154216
rect 255314 154164 255320 154216
rect 255372 154204 255378 154216
rect 314378 154204 314384 154216
rect 255372 154176 314384 154204
rect 255372 154164 255378 154176
rect 314378 154164 314384 154176
rect 314436 154164 314442 154216
rect 336826 154164 336832 154216
rect 336884 154204 336890 154216
rect 376018 154204 376024 154216
rect 336884 154176 376024 154204
rect 336884 154164 336890 154176
rect 376018 154164 376024 154176
rect 376076 154164 376082 154216
rect 383654 154164 383660 154216
rect 383712 154204 383718 154216
rect 411990 154204 411996 154216
rect 383712 154176 411996 154204
rect 383712 154164 383718 154176
rect 411990 154164 411996 154176
rect 412048 154164 412054 154216
rect 142246 154136 142252 154148
rect 129476 154040 137140 154068
rect 137204 154108 142252 154136
rect 9674 153960 9680 154012
rect 9732 154000 9738 154012
rect 126882 154000 126888 154012
rect 9732 153972 126888 154000
rect 9732 153960 9738 153972
rect 126882 153960 126888 153972
rect 126940 153960 126946 154012
rect 127618 153960 127624 154012
rect 127676 154000 127682 154012
rect 129366 154000 129372 154012
rect 127676 153972 129372 154000
rect 127676 153960 127682 153972
rect 129366 153960 129372 153972
rect 129424 153960 129430 154012
rect 7098 153892 7104 153944
rect 7156 153932 7162 153944
rect 124306 153932 124312 153944
rect 7156 153904 124312 153932
rect 7156 153892 7162 153904
rect 124306 153892 124312 153904
rect 124364 153892 124370 153944
rect 125502 153892 125508 153944
rect 125560 153932 125566 153944
rect 129476 153932 129504 154040
rect 129642 153960 129648 154012
rect 129700 154000 129706 154012
rect 137204 154000 137232 154108
rect 142246 154096 142252 154108
rect 142304 154096 142310 154148
rect 142614 154096 142620 154148
rect 142672 154136 142678 154148
rect 145558 154136 145564 154148
rect 142672 154108 145564 154136
rect 142672 154096 142678 154108
rect 145558 154096 145564 154108
rect 145616 154096 145622 154148
rect 147122 154096 147128 154148
rect 147180 154136 147186 154148
rect 147180 154108 157334 154136
rect 147180 154096 147186 154108
rect 137278 154028 137284 154080
rect 137336 154068 137342 154080
rect 139762 154068 139768 154080
rect 137336 154040 139768 154068
rect 137336 154028 137342 154040
rect 139762 154028 139768 154040
rect 139820 154028 139826 154080
rect 139854 154028 139860 154080
rect 139912 154068 139918 154080
rect 142430 154068 142436 154080
rect 139912 154040 142436 154068
rect 139912 154028 139918 154040
rect 142430 154028 142436 154040
rect 142488 154028 142494 154080
rect 142522 154028 142528 154080
rect 142580 154068 142586 154080
rect 153194 154068 153200 154080
rect 142580 154040 153200 154068
rect 142580 154028 142586 154040
rect 153194 154028 153200 154040
rect 153252 154028 153258 154080
rect 153286 154028 153292 154080
rect 153344 154068 153350 154080
rect 155954 154068 155960 154080
rect 153344 154040 155960 154068
rect 153344 154028 153350 154040
rect 155954 154028 155960 154040
rect 156012 154028 156018 154080
rect 157306 154068 157334 154108
rect 160186 154096 160192 154148
rect 160244 154136 160250 154148
rect 160244 154108 162900 154136
rect 160244 154096 160250 154108
rect 161566 154068 161572 154080
rect 157306 154040 161572 154068
rect 161566 154028 161572 154040
rect 161624 154028 161630 154080
rect 162872 154068 162900 154108
rect 165614 154096 165620 154148
rect 165672 154136 165678 154148
rect 245654 154136 245660 154148
rect 165672 154108 245660 154136
rect 165672 154096 165678 154108
rect 245654 154096 245660 154108
rect 245712 154096 245718 154148
rect 245930 154096 245936 154148
rect 245988 154136 245994 154148
rect 306650 154136 306656 154148
rect 245988 154108 306656 154136
rect 245988 154096 245994 154108
rect 306650 154096 306656 154108
rect 306708 154096 306714 154148
rect 326706 154096 326712 154148
rect 326764 154136 326770 154148
rect 368290 154136 368296 154148
rect 326764 154108 368296 154136
rect 326764 154096 326770 154108
rect 368290 154096 368296 154108
rect 368348 154096 368354 154148
rect 376846 154096 376852 154148
rect 376904 154136 376910 154148
rect 406838 154136 406844 154148
rect 376904 154108 406844 154136
rect 376904 154096 376910 154108
rect 406838 154096 406844 154108
rect 406896 154096 406902 154148
rect 241238 154068 241244 154080
rect 162872 154040 241244 154068
rect 241238 154028 241244 154040
rect 241296 154028 241302 154080
rect 248598 154028 248604 154080
rect 248656 154068 248662 154080
rect 309226 154068 309232 154080
rect 248656 154040 309232 154068
rect 248656 154028 248662 154040
rect 309226 154028 309232 154040
rect 309284 154028 309290 154080
rect 323302 154028 323308 154080
rect 323360 154068 323366 154080
rect 365806 154068 365812 154080
rect 323360 154040 365812 154068
rect 323360 154028 323366 154040
rect 365806 154028 365812 154040
rect 365864 154028 365870 154080
rect 380158 154028 380164 154080
rect 380216 154068 380222 154080
rect 409414 154068 409420 154080
rect 380216 154040 409420 154068
rect 380216 154028 380222 154040
rect 409414 154028 409420 154040
rect 409472 154028 409478 154080
rect 219894 154000 219900 154012
rect 129700 153972 137232 154000
rect 137296 153972 219900 154000
rect 129700 153960 129706 153972
rect 125560 153904 129504 153932
rect 125560 153892 125566 153904
rect 132402 153892 132408 153944
rect 132460 153932 132466 153944
rect 137296 153932 137324 153972
rect 219894 153960 219900 153972
rect 219952 153960 219958 154012
rect 222378 153960 222384 154012
rect 222436 154000 222442 154012
rect 288710 154000 288716 154012
rect 222436 153972 288716 154000
rect 222436 153960 222442 153972
rect 288710 153960 288716 153972
rect 288768 153960 288774 154012
rect 316034 153960 316040 154012
rect 316092 154000 316098 154012
rect 360654 154000 360660 154012
rect 316092 153972 360660 154000
rect 316092 153960 316098 153972
rect 360654 153960 360660 153972
rect 360712 153960 360718 154012
rect 367094 153960 367100 154012
rect 367152 154000 367158 154012
rect 399110 154000 399116 154012
rect 367152 153972 399116 154000
rect 367152 153960 367158 153972
rect 399110 153960 399116 153972
rect 399168 153960 399174 154012
rect 132460 153904 137324 153932
rect 132460 153892 132466 153904
rect 138014 153892 138020 153944
rect 138072 153932 138078 153944
rect 138072 153904 142936 153932
rect 138072 153892 138078 153904
rect 474 153824 480 153876
rect 532 153864 538 153876
rect 119798 153864 119804 153876
rect 532 153836 119804 153864
rect 532 153824 538 153836
rect 119798 153824 119804 153836
rect 119856 153824 119862 153876
rect 119890 153824 119896 153876
rect 119948 153864 119954 153876
rect 142798 153864 142804 153876
rect 119948 153836 142804 153864
rect 119948 153824 119954 153836
rect 142798 153824 142804 153836
rect 142856 153824 142862 153876
rect 142908 153864 142936 153904
rect 142982 153892 142988 153944
rect 143040 153932 143046 153944
rect 223206 153932 223212 153944
rect 143040 153904 223212 153932
rect 143040 153892 143046 153904
rect 223206 153892 223212 153904
rect 223264 153892 223270 153944
rect 225230 153892 225236 153944
rect 225288 153932 225294 153944
rect 291286 153932 291292 153944
rect 225288 153904 291292 153932
rect 225288 153892 225294 153904
rect 291286 153892 291292 153904
rect 291344 153892 291350 153944
rect 313274 153892 313280 153944
rect 313332 153932 313338 153944
rect 357894 153932 357900 153944
rect 313332 153904 357900 153932
rect 313332 153892 313338 153904
rect 357894 153892 357900 153904
rect 357952 153892 357958 153944
rect 363046 153892 363052 153944
rect 363104 153932 363110 153944
rect 396534 153932 396540 153944
rect 363104 153904 396540 153932
rect 363104 153892 363110 153904
rect 396534 153892 396540 153904
rect 396592 153892 396598 153944
rect 401594 153892 401600 153944
rect 401652 153932 401658 153944
rect 425514 153932 425520 153944
rect 401652 153904 425520 153932
rect 401652 153892 401658 153904
rect 425514 153892 425520 153904
rect 425572 153892 425578 153944
rect 152458 153864 152464 153876
rect 142908 153836 152464 153864
rect 152458 153824 152464 153836
rect 152516 153824 152522 153876
rect 154482 153824 154488 153876
rect 154540 153864 154546 153876
rect 154540 153836 155908 153864
rect 154540 153824 154546 153836
rect 48314 153756 48320 153808
rect 48372 153796 48378 153808
rect 155770 153796 155776 153808
rect 48372 153768 155776 153796
rect 48372 153756 48378 153768
rect 155770 153756 155776 153768
rect 155828 153756 155834 153808
rect 155880 153796 155908 153836
rect 155954 153824 155960 153876
rect 156012 153864 156018 153876
rect 235442 153864 235448 153876
rect 156012 153836 235448 153864
rect 156012 153824 156018 153836
rect 235442 153824 235448 153836
rect 235500 153824 235506 153876
rect 241882 153824 241888 153876
rect 241940 153864 241946 153876
rect 304074 153864 304080 153876
rect 241940 153836 304080 153864
rect 241940 153824 241946 153836
rect 304074 153824 304080 153836
rect 304132 153824 304138 153876
rect 309134 153824 309140 153876
rect 309192 153864 309198 153876
rect 355502 153864 355508 153876
rect 309192 153836 355508 153864
rect 309192 153824 309198 153836
rect 355502 153824 355508 153836
rect 355560 153824 355566 153876
rect 356238 153824 356244 153876
rect 356296 153864 356302 153876
rect 391474 153864 391480 153876
rect 356296 153836 391480 153864
rect 356296 153824 356302 153836
rect 391474 153824 391480 153836
rect 391532 153824 391538 153876
rect 397454 153824 397460 153876
rect 397512 153864 397518 153876
rect 422938 153864 422944 153876
rect 397512 153836 422944 153864
rect 397512 153824 397518 153836
rect 422938 153824 422944 153836
rect 422996 153824 423002 153876
rect 218054 153796 218060 153808
rect 155880 153768 218060 153796
rect 218054 153756 218060 153768
rect 218112 153756 218118 153808
rect 231854 153756 231860 153808
rect 231912 153796 231918 153808
rect 296438 153796 296444 153808
rect 231912 153768 296444 153796
rect 231912 153756 231918 153768
rect 296438 153756 296444 153768
rect 296496 153756 296502 153808
rect 360378 153756 360384 153808
rect 360436 153796 360442 153808
rect 394050 153796 394056 153808
rect 360436 153768 394056 153796
rect 360436 153756 360442 153768
rect 394050 153756 394056 153768
rect 394108 153756 394114 153808
rect 61102 153688 61108 153740
rect 61160 153728 61166 153740
rect 161474 153728 161480 153740
rect 61160 153700 161480 153728
rect 61160 153688 61166 153700
rect 161474 153688 161480 153700
rect 161532 153688 161538 153740
rect 161566 153688 161572 153740
rect 161624 153728 161630 153740
rect 210418 153728 210424 153740
rect 161624 153700 210424 153728
rect 161624 153688 161630 153700
rect 210418 153688 210424 153700
rect 210476 153688 210482 153740
rect 235074 153688 235080 153740
rect 235132 153728 235138 153740
rect 299014 153728 299020 153740
rect 235132 153700 299020 153728
rect 235132 153688 235138 153700
rect 299014 153688 299020 153700
rect 299072 153688 299078 153740
rect 57974 153620 57980 153672
rect 58032 153660 58038 153672
rect 152366 153660 152372 153672
rect 58032 153632 152372 153660
rect 58032 153620 58038 153632
rect 152366 153620 152372 153632
rect 152424 153620 152430 153672
rect 152458 153620 152464 153672
rect 152516 153660 152522 153672
rect 191006 153660 191012 153672
rect 152516 153632 191012 153660
rect 152516 153620 152522 153632
rect 191006 153620 191012 153632
rect 191064 153620 191070 153672
rect 191742 153620 191748 153672
rect 191800 153660 191806 153672
rect 195882 153660 195888 153672
rect 191800 153632 195888 153660
rect 191800 153620 191806 153632
rect 195882 153620 195888 153632
rect 195940 153620 195946 153672
rect 195974 153620 195980 153672
rect 196032 153660 196038 153672
rect 209774 153660 209780 153672
rect 196032 153632 209780 153660
rect 196032 153620 196038 153632
rect 209774 153620 209780 153632
rect 209832 153620 209838 153672
rect 229094 153620 229100 153672
rect 229152 153660 229158 153672
rect 293862 153660 293868 153672
rect 229152 153632 293868 153660
rect 229152 153620 229158 153632
rect 293862 153620 293868 153632
rect 293920 153620 293926 153672
rect 78674 153552 78680 153604
rect 78732 153592 78738 153604
rect 179598 153592 179604 153604
rect 78732 153564 179604 153592
rect 78732 153552 78738 153564
rect 179598 153552 179604 153564
rect 179656 153552 179662 153604
rect 179690 153552 179696 153604
rect 179748 153592 179754 153604
rect 230934 153592 230940 153604
rect 179748 153564 230940 153592
rect 179748 153552 179754 153564
rect 230934 153552 230940 153564
rect 230992 153552 230998 153604
rect 238846 153552 238852 153604
rect 238904 153592 238910 153604
rect 301590 153592 301596 153604
rect 238904 153564 301596 153592
rect 238904 153552 238910 153564
rect 301590 153552 301596 153564
rect 301648 153552 301654 153604
rect 102134 153484 102140 153536
rect 102192 153524 102198 153536
rect 196894 153524 196900 153536
rect 102192 153496 196900 153524
rect 102192 153484 102198 153496
rect 196894 153484 196900 153496
rect 196952 153484 196958 153536
rect 196986 153484 196992 153536
rect 197044 153524 197050 153536
rect 200850 153524 200856 153536
rect 197044 153496 200856 153524
rect 197044 153484 197050 153496
rect 200850 153484 200856 153496
rect 200908 153484 200914 153536
rect 201126 153484 201132 153536
rect 201184 153524 201190 153536
rect 205266 153524 205272 153536
rect 201184 153496 205272 153524
rect 201184 153484 201190 153496
rect 205266 153484 205272 153496
rect 205324 153484 205330 153536
rect 205358 153484 205364 153536
rect 205416 153524 205422 153536
rect 248874 153524 248880 153536
rect 205416 153496 248880 153524
rect 205416 153484 205422 153496
rect 248874 153484 248880 153496
rect 248932 153484 248938 153536
rect 252646 153484 252652 153536
rect 252704 153524 252710 153536
rect 311802 153524 311808 153536
rect 252704 153496 311808 153524
rect 252704 153484 252710 153496
rect 311802 153484 311808 153496
rect 311860 153484 311866 153536
rect 104894 153416 104900 153468
rect 104952 153456 104958 153468
rect 199470 153456 199476 153468
rect 104952 153428 199476 153456
rect 104952 153416 104958 153428
rect 199470 153416 199476 153428
rect 199528 153416 199534 153468
rect 207842 153456 207848 153468
rect 200684 153428 207848 153456
rect 108298 153348 108304 153400
rect 108356 153388 108362 153400
rect 191190 153388 191196 153400
rect 108356 153360 191196 153388
rect 108356 153348 108362 153360
rect 191190 153348 191196 153360
rect 191248 153348 191254 153400
rect 191282 153348 191288 153400
rect 191340 153388 191346 153400
rect 197538 153388 197544 153400
rect 191340 153360 197544 153388
rect 191340 153348 191346 153360
rect 197538 153348 197544 153360
rect 197596 153348 197602 153400
rect 198918 153348 198924 153400
rect 198976 153388 198982 153400
rect 200574 153388 200580 153400
rect 198976 153360 200580 153388
rect 198976 153348 198982 153360
rect 200574 153348 200580 153360
rect 200632 153348 200638 153400
rect 115934 153280 115940 153332
rect 115992 153320 115998 153332
rect 200684 153320 200712 153428
rect 207842 153416 207848 153428
rect 207900 153416 207906 153468
rect 207934 153416 207940 153468
rect 207992 153456 207998 153468
rect 259178 153456 259184 153468
rect 207992 153428 259184 153456
rect 207992 153416 207998 153428
rect 259178 153416 259184 153428
rect 259236 153416 259242 153468
rect 265434 153416 265440 153468
rect 265492 153456 265498 153468
rect 322014 153456 322020 153468
rect 265492 153428 322020 153456
rect 265492 153416 265498 153428
rect 322014 153416 322020 153428
rect 322072 153416 322078 153468
rect 200758 153348 200764 153400
rect 200816 153388 200822 153400
rect 205358 153388 205364 153400
rect 200816 153360 205364 153388
rect 200816 153348 200822 153360
rect 205358 153348 205364 153360
rect 205416 153348 205422 153400
rect 243722 153388 243728 153400
rect 205468 153360 243728 153388
rect 115992 153292 200712 153320
rect 115992 153280 115998 153292
rect 200850 153280 200856 153332
rect 200908 153320 200914 153332
rect 205468 153320 205496 153360
rect 243722 153348 243728 153360
rect 243780 153348 243786 153400
rect 259454 153348 259460 153400
rect 259512 153388 259518 153400
rect 316954 153388 316960 153400
rect 259512 153360 316960 153388
rect 259512 153348 259518 153360
rect 316954 153348 316960 153360
rect 317012 153348 317018 153400
rect 238662 153320 238668 153332
rect 200908 153292 205496 153320
rect 205606 153292 238668 153320
rect 200908 153280 200914 153292
rect 41598 153212 41604 153264
rect 41656 153252 41662 153264
rect 142706 153252 142712 153264
rect 41656 153224 142712 153252
rect 41656 153212 41662 153224
rect 142706 153212 142712 153224
rect 142764 153212 142770 153264
rect 142798 153212 142804 153264
rect 142856 153252 142862 153264
rect 195974 153252 195980 153264
rect 142856 153224 195980 153252
rect 142856 153212 142862 153224
rect 195974 153212 195980 153224
rect 196032 153212 196038 153264
rect 196066 153212 196072 153264
rect 196124 153252 196130 153264
rect 205606 153252 205634 153292
rect 238662 153280 238668 153292
rect 238720 153280 238726 153332
rect 272886 153280 272892 153332
rect 272944 153320 272950 153332
rect 327258 153320 327264 153332
rect 272944 153292 327264 153320
rect 272944 153280 272950 153292
rect 327258 153280 327264 153292
rect 327316 153280 327322 153332
rect 196124 153224 205634 153252
rect 196124 153212 196130 153224
rect 269206 153212 269212 153264
rect 269264 153252 269270 153264
rect 324682 153252 324688 153264
rect 269264 153224 324688 153252
rect 269264 153212 269270 153224
rect 324682 153212 324688 153224
rect 324740 153212 324746 153264
rect 23290 153144 23296 153196
rect 23348 153184 23354 153196
rect 110966 153184 110972 153196
rect 23348 153156 110972 153184
rect 23348 153144 23354 153156
rect 110966 153144 110972 153156
rect 111024 153144 111030 153196
rect 113174 153144 113180 153196
rect 113232 153184 113238 153196
rect 205910 153184 205916 153196
rect 113232 153156 205916 153184
rect 113232 153144 113238 153156
rect 205910 153144 205916 153156
rect 205968 153144 205974 153196
rect 215386 153144 215392 153196
rect 215444 153184 215450 153196
rect 279694 153184 279700 153196
rect 215444 153156 279700 153184
rect 215444 153144 215450 153156
rect 279694 153144 279700 153156
rect 279752 153144 279758 153196
rect 285490 153144 285496 153196
rect 285548 153184 285554 153196
rect 336826 153184 336832 153196
rect 285548 153156 336832 153184
rect 285548 153144 285554 153156
rect 336826 153144 336832 153156
rect 336884 153144 336890 153196
rect 339678 153144 339684 153196
rect 339736 153184 339742 153196
rect 377306 153184 377312 153196
rect 339736 153156 377312 153184
rect 339736 153144 339742 153156
rect 377306 153144 377312 153156
rect 377364 153144 377370 153196
rect 378226 153144 378232 153196
rect 378284 153184 378290 153196
rect 379882 153184 379888 153196
rect 378284 153156 379888 153184
rect 378284 153144 378290 153156
rect 379882 153144 379888 153156
rect 379940 153144 379946 153196
rect 385494 153144 385500 153196
rect 385552 153184 385558 153196
rect 387610 153184 387616 153196
rect 385552 153156 387616 153184
rect 385552 153144 385558 153156
rect 387610 153144 387616 153156
rect 387668 153144 387674 153196
rect 389174 153144 389180 153196
rect 389232 153184 389238 153196
rect 393498 153184 393504 153196
rect 389232 153156 393504 153184
rect 389232 153144 389238 153156
rect 393498 153144 393504 153156
rect 393556 153144 393562 153196
rect 395522 153144 395528 153196
rect 395580 153184 395586 153196
rect 397822 153184 397828 153196
rect 395580 153156 397828 153184
rect 395580 153144 395586 153156
rect 397822 153144 397828 153156
rect 397880 153144 397886 153196
rect 397914 153144 397920 153196
rect 397972 153184 397978 153196
rect 415210 153184 415216 153196
rect 397972 153156 415216 153184
rect 397972 153144 397978 153156
rect 415210 153144 415216 153156
rect 415268 153144 415274 153196
rect 418154 153144 418160 153196
rect 418212 153184 418218 153196
rect 437566 153184 437572 153196
rect 418212 153156 437572 153184
rect 418212 153144 418218 153156
rect 437566 153144 437572 153156
rect 437624 153144 437630 153196
rect 437842 153144 437848 153196
rect 437900 153184 437906 153196
rect 446398 153184 446404 153196
rect 437900 153156 446404 153184
rect 437900 153144 437906 153156
rect 446398 153144 446404 153156
rect 446456 153144 446462 153196
rect 456794 153144 456800 153196
rect 456852 153184 456858 153196
rect 459462 153184 459468 153196
rect 456852 153156 459468 153184
rect 456852 153144 456858 153156
rect 459462 153144 459468 153156
rect 459520 153144 459526 153196
rect 461854 153144 461860 153196
rect 461912 153184 461918 153196
rect 465902 153184 465908 153196
rect 461912 153156 465908 153184
rect 461912 153144 461918 153156
rect 465902 153144 465908 153156
rect 465960 153144 465966 153196
rect 466454 153144 466460 153196
rect 466512 153184 466518 153196
rect 470410 153184 470416 153196
rect 466512 153156 470416 153184
rect 466512 153144 466518 153156
rect 470410 153144 470416 153156
rect 470468 153144 470474 153196
rect 471514 153144 471520 153196
rect 471572 153184 471578 153196
rect 473630 153184 473636 153196
rect 471572 153156 473636 153184
rect 471572 153144 471578 153156
rect 473630 153144 473636 153156
rect 473688 153144 473694 153196
rect 474826 153144 474832 153196
rect 474884 153184 474890 153196
rect 476942 153184 476948 153196
rect 474884 153156 476948 153184
rect 474884 153144 474890 153156
rect 476942 153144 476948 153156
rect 477000 153144 477006 153196
rect 485682 153144 485688 153196
rect 485740 153184 485746 153196
rect 489638 153184 489644 153196
rect 485740 153156 489644 153184
rect 485740 153144 485746 153156
rect 489638 153144 489644 153156
rect 489696 153144 489702 153196
rect 490742 153144 490748 153196
rect 490800 153184 490806 153196
rect 493502 153184 493508 153196
rect 490800 153156 493508 153184
rect 490800 153144 490806 153156
rect 493502 153144 493508 153156
rect 493560 153144 493566 153196
rect 494054 153144 494060 153196
rect 494112 153184 494118 153196
rect 496078 153184 496084 153196
rect 494112 153156 496084 153184
rect 494112 153144 494118 153156
rect 496078 153144 496084 153156
rect 496136 153144 496142 153196
rect 496630 153144 496636 153196
rect 496688 153184 496694 153196
rect 498010 153184 498016 153196
rect 496688 153156 498016 153184
rect 496688 153144 496694 153156
rect 498010 153144 498016 153156
rect 498068 153144 498074 153196
rect 512270 153144 512276 153196
rect 512328 153184 512334 153196
rect 514846 153184 514852 153196
rect 512328 153156 514852 153184
rect 512328 153144 512334 153156
rect 514846 153144 514852 153156
rect 514904 153144 514910 153196
rect 80054 153076 80060 153128
rect 80112 153116 80118 153128
rect 175090 153116 175096 153128
rect 80112 153088 175096 153116
rect 80112 153076 80118 153088
rect 175090 153076 175096 153088
rect 175148 153076 175154 153128
rect 180794 153076 180800 153128
rect 180852 153116 180858 153128
rect 257246 153116 257252 153128
rect 180852 153088 257252 153116
rect 180852 153076 180858 153088
rect 257246 153076 257252 153088
rect 257304 153076 257310 153128
rect 264974 153076 264980 153128
rect 265032 153116 265038 153128
rect 321462 153116 321468 153128
rect 265032 153088 321468 153116
rect 265032 153076 265038 153088
rect 321462 153076 321468 153088
rect 321520 153076 321526 153128
rect 324314 153076 324320 153128
rect 324372 153116 324378 153128
rect 367002 153116 367008 153128
rect 324372 153088 367008 153116
rect 324372 153076 324378 153088
rect 367002 153076 367008 153088
rect 367060 153076 367066 153128
rect 367186 153076 367192 153128
rect 367244 153116 367250 153128
rect 368934 153116 368940 153128
rect 367244 153088 368940 153116
rect 367244 153076 367250 153088
rect 368934 153076 368940 153088
rect 368992 153076 368998 153128
rect 382182 153076 382188 153128
rect 382240 153116 382246 153128
rect 410702 153116 410708 153128
rect 382240 153088 410708 153116
rect 382240 153076 382246 153088
rect 410702 153076 410708 153088
rect 410760 153076 410766 153128
rect 412910 153076 412916 153128
rect 412968 153116 412974 153128
rect 422202 153116 422208 153128
rect 412968 153088 422208 153116
rect 412968 153076 412974 153088
rect 422202 153076 422208 153088
rect 422260 153076 422266 153128
rect 422294 153076 422300 153128
rect 422352 153116 422358 153128
rect 423122 153116 423128 153128
rect 422352 153088 423128 153116
rect 422352 153076 422358 153088
rect 423122 153076 423128 153088
rect 423180 153076 423186 153128
rect 425146 153076 425152 153128
rect 425204 153116 425210 153128
rect 434622 153116 434628 153128
rect 425204 153088 434628 153116
rect 425204 153076 425210 153088
rect 434622 153076 434628 153088
rect 434680 153076 434686 153128
rect 434714 153076 434720 153128
rect 434772 153116 434778 153128
rect 443914 153116 443920 153128
rect 434772 153088 443920 153116
rect 434772 153076 434778 153088
rect 443914 153076 443920 153088
rect 443972 153076 443978 153128
rect 444006 153076 444012 153128
rect 444064 153116 444070 153128
rect 450538 153116 450544 153128
rect 444064 153088 450544 153116
rect 444064 153076 444070 153088
rect 450538 153076 450544 153088
rect 450596 153076 450602 153128
rect 462774 153076 462780 153128
rect 462832 153116 462838 153128
rect 466546 153116 466552 153128
rect 462832 153088 466552 153116
rect 462832 153076 462838 153088
rect 466546 153076 466552 153088
rect 466604 153076 466610 153128
rect 466638 153076 466644 153128
rect 466696 153116 466702 153128
rect 469766 153116 469772 153128
rect 466696 153088 469772 153116
rect 466696 153076 466702 153088
rect 469766 153076 469772 153088
rect 469824 153076 469830 153128
rect 472250 153076 472256 153128
rect 472308 153116 472314 153128
rect 474274 153116 474280 153128
rect 472308 153088 474280 153116
rect 472308 153076 472314 153088
rect 474274 153076 474280 153088
rect 474332 153076 474338 153128
rect 476114 153076 476120 153128
rect 476172 153116 476178 153128
rect 478138 153116 478144 153128
rect 476172 153088 478144 153116
rect 476172 153076 476178 153088
rect 478138 153076 478144 153088
rect 478196 153076 478202 153128
rect 484026 153076 484032 153128
rect 484084 153116 484090 153128
rect 488442 153116 488448 153128
rect 484084 153088 488448 153116
rect 484084 153076 484090 153088
rect 488442 153076 488448 153088
rect 488500 153076 488506 153128
rect 492398 153076 492404 153128
rect 492456 153116 492462 153128
rect 494790 153116 494796 153128
rect 492456 153088 494796 153116
rect 492456 153076 492462 153088
rect 494790 153076 494796 153088
rect 494848 153076 494854 153128
rect 494974 153076 494980 153128
rect 495032 153116 495038 153128
rect 496722 153116 496728 153128
rect 495032 153088 496728 153116
rect 495032 153076 495038 153088
rect 496722 153076 496728 153088
rect 496780 153076 496786 153128
rect 496814 153076 496820 153128
rect 496872 153116 496878 153128
rect 498654 153116 498660 153128
rect 496872 153088 498660 153116
rect 496872 153076 496878 153088
rect 498654 153076 498660 153088
rect 498712 153076 498718 153128
rect 510982 153076 510988 153128
rect 511040 153116 511046 153128
rect 513466 153116 513472 153128
rect 511040 153088 513472 153116
rect 511040 153076 511046 153088
rect 513466 153076 513472 153088
rect 513524 153076 513530 153128
rect 513558 153076 513564 153128
rect 513616 153116 513622 153128
rect 516134 153116 516140 153128
rect 513616 153088 516140 153116
rect 513616 153076 513622 153088
rect 516134 153076 516140 153088
rect 516192 153076 516198 153128
rect 103514 153008 103520 153060
rect 103572 153048 103578 153060
rect 198182 153048 198188 153060
rect 103572 153020 198188 153048
rect 103572 153008 103578 153020
rect 198182 153008 198188 153020
rect 198240 153008 198246 153060
rect 203702 153008 203708 153060
rect 203760 153048 203766 153060
rect 267550 153048 267556 153060
rect 203760 153020 267556 153048
rect 203760 153008 203766 153020
rect 267550 153008 267556 153020
rect 267608 153008 267614 153060
rect 272150 153008 272156 153060
rect 272208 153048 272214 153060
rect 326614 153048 326620 153060
rect 272208 153020 326620 153048
rect 272208 153008 272214 153020
rect 326614 153008 326620 153020
rect 326672 153008 326678 153060
rect 330938 153008 330944 153060
rect 330996 153048 331002 153060
rect 371510 153048 371516 153060
rect 330996 153020 371516 153048
rect 330996 153008 331002 153020
rect 371510 153008 371516 153020
rect 371568 153008 371574 153060
rect 372614 153008 372620 153060
rect 372672 153048 372678 153060
rect 403618 153048 403624 153060
rect 372672 153020 403624 153048
rect 372672 153008 372678 153020
rect 403618 153008 403624 153020
rect 403676 153008 403682 153060
rect 405826 153008 405832 153060
rect 405884 153048 405890 153060
rect 408770 153048 408776 153060
rect 405884 153020 408776 153048
rect 405884 153008 405890 153020
rect 408770 153008 408776 153020
rect 408828 153008 408834 153060
rect 410518 153008 410524 153060
rect 410576 153048 410582 153060
rect 431126 153048 431132 153060
rect 410576 153020 431132 153048
rect 410576 153008 410582 153020
rect 431126 153008 431132 153020
rect 431184 153008 431190 153060
rect 431954 153008 431960 153060
rect 432012 153048 432018 153060
rect 441982 153048 441988 153060
rect 432012 153020 441988 153048
rect 432012 153008 432018 153020
rect 441982 153008 441988 153020
rect 442040 153008 442046 153060
rect 442074 153008 442080 153060
rect 442132 153048 442138 153060
rect 447410 153048 447416 153060
rect 442132 153020 447416 153048
rect 442132 153008 442138 153020
rect 447410 153008 447416 153020
rect 447468 153008 447474 153060
rect 463142 153008 463148 153060
rect 463200 153048 463206 153060
rect 467190 153048 467196 153060
rect 463200 153020 467196 153048
rect 463200 153008 463206 153020
rect 467190 153008 467196 153020
rect 467248 153008 467254 153060
rect 472618 153008 472624 153060
rect 472676 153048 472682 153060
rect 474918 153048 474924 153060
rect 472676 153020 474924 153048
rect 472676 153008 472682 153020
rect 474918 153008 474924 153020
rect 474976 153008 474982 153060
rect 484486 153008 484492 153060
rect 484544 153048 484550 153060
rect 488994 153048 489000 153060
rect 484544 153020 489000 153048
rect 484544 153008 484550 153020
rect 488994 153008 489000 153020
rect 489052 153008 489058 153060
rect 492674 153008 492680 153060
rect 492732 153048 492738 153060
rect 495434 153048 495440 153060
rect 492732 153020 495440 153048
rect 492732 153008 492738 153020
rect 495434 153008 495440 153020
rect 495492 153008 495498 153060
rect 495526 153008 495532 153060
rect 495584 153048 495590 153060
rect 497366 153048 497372 153060
rect 495584 153020 497372 153048
rect 495584 153008 495590 153020
rect 497366 153008 497372 153020
rect 497424 153008 497430 153060
rect 511626 153008 511632 153060
rect 511684 153048 511690 153060
rect 514294 153048 514300 153060
rect 511684 153020 514300 153048
rect 511684 153008 511690 153020
rect 514294 153008 514300 153020
rect 514352 153008 514358 153060
rect 92566 152940 92572 152992
rect 92624 152980 92630 152992
rect 187878 152980 187884 152992
rect 92624 152952 187884 152980
rect 92624 152940 92630 152952
rect 187878 152940 187884 152952
rect 187936 152940 187942 152992
rect 195054 152940 195060 152992
rect 195112 152980 195118 152992
rect 218698 152980 218704 152992
rect 195112 152952 218704 152980
rect 195112 152940 195118 152952
rect 218698 152940 218704 152952
rect 218756 152940 218762 152992
rect 220354 152940 220360 152992
rect 220412 152980 220418 152992
rect 284846 152980 284852 152992
rect 220412 152952 284852 152980
rect 220412 152940 220418 152952
rect 284846 152940 284852 152952
rect 284904 152940 284910 152992
rect 288066 152940 288072 152992
rect 288124 152980 288130 152992
rect 289998 152980 290004 152992
rect 288124 152952 290004 152980
rect 288124 152940 288130 152952
rect 289998 152940 290004 152952
rect 290056 152940 290062 152992
rect 292206 152940 292212 152992
rect 292264 152980 292270 152992
rect 341978 152980 341984 152992
rect 292264 152952 341984 152980
rect 292264 152940 292270 152952
rect 341978 152940 341984 152952
rect 342036 152940 342042 152992
rect 342254 152940 342260 152992
rect 342312 152980 342318 152992
rect 343910 152980 343916 152992
rect 342312 152952 343916 152980
rect 342312 152940 342318 152952
rect 343910 152940 343916 152952
rect 343968 152940 343974 152992
rect 345290 152940 345296 152992
rect 345348 152980 345354 152992
rect 382458 152980 382464 152992
rect 345348 152952 382464 152980
rect 345348 152940 345354 152952
rect 382458 152940 382464 152952
rect 382516 152940 382522 152992
rect 384942 152940 384948 152992
rect 385000 152980 385006 152992
rect 392118 152980 392124 152992
rect 385000 152952 392124 152980
rect 385000 152940 385006 152952
rect 392118 152940 392124 152952
rect 392176 152940 392182 152992
rect 394878 152940 394884 152992
rect 394936 152980 394942 152992
rect 415302 152980 415308 152992
rect 394936 152952 415308 152980
rect 394936 152940 394942 152952
rect 415302 152940 415308 152952
rect 415360 152940 415366 152992
rect 415394 152940 415400 152992
rect 415452 152980 415458 152992
rect 415452 152952 418154 152980
rect 415452 152940 415458 152952
rect 71406 152872 71412 152924
rect 71464 152912 71470 152924
rect 92474 152912 92480 152924
rect 71464 152884 92480 152912
rect 71464 152872 71470 152884
rect 92474 152872 92480 152884
rect 92532 152872 92538 152924
rect 96614 152872 96620 152924
rect 96672 152912 96678 152924
rect 193030 152912 193036 152924
rect 96672 152884 193036 152912
rect 96672 152872 96678 152884
rect 193030 152872 193036 152884
rect 193088 152872 193094 152924
rect 212442 152872 212448 152924
rect 212500 152912 212506 152924
rect 277762 152912 277768 152924
rect 212500 152884 277768 152912
rect 212500 152872 212506 152884
rect 277762 152872 277768 152884
rect 277820 152872 277826 152924
rect 278774 152872 278780 152924
rect 278832 152912 278838 152924
rect 331766 152912 331772 152924
rect 278832 152884 331772 152912
rect 278832 152872 278838 152884
rect 331766 152872 331772 152884
rect 331824 152872 331830 152924
rect 332594 152872 332600 152924
rect 332652 152912 332658 152924
rect 372798 152912 372804 152924
rect 332652 152884 372804 152912
rect 332652 152872 332658 152884
rect 372798 152872 372804 152884
rect 372856 152872 372862 152924
rect 375466 152872 375472 152924
rect 375524 152912 375530 152924
rect 405550 152912 405556 152924
rect 375524 152884 405556 152912
rect 375524 152872 375530 152884
rect 405550 152872 405556 152884
rect 405608 152872 405614 152924
rect 406654 152872 406660 152924
rect 406712 152912 406718 152924
rect 417602 152912 417608 152924
rect 406712 152884 417608 152912
rect 406712 152872 406718 152884
rect 417602 152872 417608 152884
rect 417660 152872 417666 152924
rect 418126 152912 418154 152952
rect 421006 152940 421012 152992
rect 421064 152980 421070 152992
rect 421064 152952 436508 152980
rect 421064 152940 421070 152952
rect 436370 152912 436376 152924
rect 418126 152884 436376 152912
rect 436370 152872 436376 152884
rect 436428 152872 436434 152924
rect 436480 152912 436508 152952
rect 437566 152940 437572 152992
rect 437624 152980 437630 152992
rect 438302 152980 438308 152992
rect 437624 152952 438308 152980
rect 437624 152940 437630 152952
rect 438302 152940 438308 152952
rect 438360 152940 438366 152992
rect 439038 152980 439044 152992
rect 438412 152952 439044 152980
rect 438412 152912 438440 152952
rect 439038 152940 439044 152952
rect 439096 152940 439102 152992
rect 440326 152940 440332 152992
rect 440384 152980 440390 152992
rect 455690 152980 455696 152992
rect 440384 152952 455696 152980
rect 440384 152940 440390 152952
rect 455690 152940 455696 152952
rect 455748 152940 455754 152992
rect 464154 152940 464160 152992
rect 464212 152980 464218 152992
rect 467834 152980 467840 152992
rect 464212 152952 467840 152980
rect 464212 152940 464218 152952
rect 467834 152940 467840 152952
rect 467892 152940 467898 152992
rect 471422 152940 471428 152992
rect 471480 152980 471486 152992
rect 472986 152980 472992 152992
rect 471480 152952 472992 152980
rect 471480 152940 471486 152952
rect 472986 152940 472992 152952
rect 473044 152940 473050 152992
rect 473354 152940 473360 152992
rect 473412 152980 473418 152992
rect 475562 152980 475568 152992
rect 473412 152952 475568 152980
rect 473412 152940 473418 152952
rect 475562 152940 475568 152952
rect 475620 152940 475626 152992
rect 483106 152940 483112 152992
rect 483164 152980 483170 152992
rect 487798 152980 487804 152992
rect 483164 152952 487804 152980
rect 483164 152940 483170 152952
rect 487798 152940 487804 152952
rect 487856 152940 487862 152992
rect 491570 152940 491576 152992
rect 491628 152980 491634 152992
rect 494146 152980 494152 152992
rect 491628 152952 494152 152980
rect 491628 152940 491634 152952
rect 494146 152940 494152 152952
rect 494204 152940 494210 152992
rect 512914 152940 512920 152992
rect 512972 152980 512978 152992
rect 515950 152980 515956 152992
rect 512972 152952 515956 152980
rect 512972 152940 512978 152952
rect 515950 152940 515956 152952
rect 516008 152940 516014 152992
rect 436480 152884 438440 152912
rect 438854 152872 438860 152924
rect 438912 152912 438918 152924
rect 454402 152912 454408 152924
rect 438912 152884 454408 152912
rect 438912 152872 438918 152884
rect 454402 152872 454408 152884
rect 454460 152872 454466 152924
rect 464430 152872 464436 152924
rect 464488 152912 464494 152924
rect 468386 152912 468392 152924
rect 464488 152884 468392 152912
rect 464488 152872 464494 152884
rect 468386 152872 468392 152884
rect 468444 152872 468450 152924
rect 489914 152872 489920 152924
rect 489972 152912 489978 152924
rect 492858 152912 492864 152924
rect 489972 152884 492864 152912
rect 489972 152872 489978 152884
rect 492858 152872 492864 152884
rect 492916 152872 492922 152924
rect 514202 152872 514208 152924
rect 514260 152912 514266 152924
rect 517422 152912 517428 152924
rect 514260 152884 517428 152912
rect 514260 152872 514266 152884
rect 517422 152872 517428 152884
rect 517480 152872 517486 152924
rect 33134 152804 33140 152856
rect 33192 152844 33198 152856
rect 138014 152844 138020 152856
rect 33192 152816 138020 152844
rect 33192 152804 33198 152816
rect 138014 152804 138020 152816
rect 138072 152804 138078 152856
rect 138106 152804 138112 152856
rect 138164 152844 138170 152856
rect 141694 152844 141700 152856
rect 138164 152816 141700 152844
rect 138164 152804 138170 152816
rect 141694 152804 141700 152816
rect 141752 152804 141758 152856
rect 146570 152804 146576 152856
rect 146628 152844 146634 152856
rect 167362 152844 167368 152856
rect 146628 152816 167368 152844
rect 146628 152804 146634 152816
rect 167362 152804 167368 152816
rect 167420 152804 167426 152856
rect 173894 152804 173900 152856
rect 173952 152844 173958 152856
rect 252094 152844 252100 152856
rect 173952 152816 252100 152844
rect 173952 152804 173958 152816
rect 252094 152804 252100 152816
rect 252152 152804 252158 152856
rect 255406 152804 255412 152856
rect 255464 152844 255470 152856
rect 313090 152844 313096 152856
rect 255464 152816 313096 152844
rect 255464 152804 255470 152816
rect 313090 152804 313096 152816
rect 313148 152804 313154 152856
rect 317046 152804 317052 152856
rect 317104 152844 317110 152856
rect 318242 152844 318248 152856
rect 317104 152816 318248 152844
rect 317104 152804 317110 152816
rect 318242 152804 318248 152816
rect 318300 152804 318306 152856
rect 320266 152804 320272 152856
rect 320324 152844 320330 152856
rect 323118 152844 323124 152856
rect 320324 152816 323124 152844
rect 320324 152804 320330 152816
rect 323118 152804 323124 152816
rect 323176 152804 323182 152856
rect 324222 152804 324228 152856
rect 324280 152844 324286 152856
rect 366358 152844 366364 152856
rect 324280 152816 366364 152844
rect 324280 152804 324286 152816
rect 366358 152804 366364 152816
rect 366416 152804 366422 152856
rect 371326 152804 371332 152856
rect 371384 152844 371390 152856
rect 402330 152844 402336 152856
rect 371384 152816 402336 152844
rect 371384 152804 371390 152816
rect 402330 152804 402336 152816
rect 402388 152804 402394 152856
rect 411254 152804 411260 152856
rect 411312 152844 411318 152856
rect 433150 152844 433156 152856
rect 411312 152816 433156 152844
rect 411312 152804 411318 152816
rect 433150 152804 433156 152816
rect 433208 152804 433214 152856
rect 434346 152804 434352 152856
rect 434404 152844 434410 152856
rect 444006 152844 444012 152856
rect 434404 152816 444012 152844
rect 434404 152804 434410 152816
rect 444006 152804 444012 152816
rect 444064 152804 444070 152856
rect 446674 152844 446680 152856
rect 444116 152816 446680 152844
rect 26418 152736 26424 152788
rect 26476 152776 26482 152788
rect 139118 152776 139124 152788
rect 26476 152748 139124 152776
rect 26476 152736 26482 152748
rect 139118 152736 139124 152748
rect 139176 152736 139182 152788
rect 140774 152736 140780 152788
rect 140832 152776 140838 152788
rect 144270 152776 144276 152788
rect 140832 152748 144276 152776
rect 140832 152736 140838 152748
rect 144270 152736 144276 152748
rect 144328 152736 144334 152788
rect 144362 152736 144368 152788
rect 144420 152776 144426 152788
rect 162210 152776 162216 152788
rect 144420 152748 162216 152776
rect 144420 152736 144426 152748
rect 162210 152736 162216 152748
rect 162268 152736 162274 152788
rect 164418 152736 164424 152788
rect 164476 152776 164482 152788
rect 244366 152776 244372 152788
rect 164476 152748 244372 152776
rect 164476 152736 164482 152748
rect 244366 152736 244372 152748
rect 244424 152736 244430 152788
rect 257706 152736 257712 152788
rect 257764 152776 257770 152788
rect 315666 152776 315672 152788
rect 257764 152748 315672 152776
rect 257764 152736 257770 152748
rect 315666 152736 315672 152748
rect 315724 152736 315730 152788
rect 317414 152736 317420 152788
rect 317472 152776 317478 152788
rect 361298 152776 361304 152788
rect 317472 152748 361304 152776
rect 317472 152736 317478 152748
rect 361298 152736 361304 152748
rect 361356 152736 361362 152788
rect 361574 152736 361580 152788
rect 361632 152776 361638 152788
rect 395338 152776 395344 152788
rect 361632 152748 395344 152776
rect 361632 152736 361638 152748
rect 395338 152736 395344 152748
rect 395396 152736 395402 152788
rect 398834 152736 398840 152788
rect 398892 152776 398898 152788
rect 403802 152776 403808 152788
rect 398892 152748 403808 152776
rect 398892 152736 398898 152748
rect 403802 152736 403808 152748
rect 403860 152736 403866 152788
rect 404354 152736 404360 152788
rect 404412 152776 404418 152788
rect 427998 152776 428004 152788
rect 404412 152748 428004 152776
rect 404412 152736 404418 152748
rect 427998 152736 428004 152748
rect 428056 152736 428062 152788
rect 429286 152736 429292 152788
rect 429344 152776 429350 152788
rect 444116 152776 444144 152816
rect 446674 152804 446680 152816
rect 446732 152804 446738 152856
rect 446766 152804 446772 152856
rect 446824 152844 446830 152856
rect 452470 152844 452476 152856
rect 446824 152816 452476 152844
rect 446824 152804 446830 152816
rect 452470 152804 452476 152816
rect 452528 152804 452534 152856
rect 465074 152804 465080 152856
rect 465132 152844 465138 152856
rect 469122 152844 469128 152856
rect 465132 152816 469128 152844
rect 465132 152804 465138 152816
rect 469122 152804 469128 152816
rect 469180 152804 469186 152856
rect 510338 152804 510344 152856
rect 510396 152844 510402 152856
rect 511994 152844 512000 152856
rect 510396 152816 512000 152844
rect 510396 152804 510402 152816
rect 511994 152804 512000 152816
rect 512052 152804 512058 152856
rect 429344 152748 444144 152776
rect 429344 152736 429350 152748
rect 444466 152736 444472 152788
rect 444524 152776 444530 152788
rect 444524 152748 444880 152776
rect 444524 152736 444530 152748
rect 28166 152668 28172 152720
rect 28224 152708 28230 152720
rect 141050 152708 141056 152720
rect 28224 152680 141056 152708
rect 28224 152668 28230 152680
rect 141050 152668 141056 152680
rect 141108 152668 141114 152720
rect 142798 152668 142804 152720
rect 142856 152708 142862 152720
rect 149422 152708 149428 152720
rect 142856 152680 149428 152708
rect 142856 152668 142862 152680
rect 149422 152668 149428 152680
rect 149480 152668 149486 152720
rect 149514 152668 149520 152720
rect 149572 152708 149578 152720
rect 231578 152708 231584 152720
rect 149572 152680 231584 152708
rect 149572 152668 149578 152680
rect 231578 152668 231584 152680
rect 231636 152668 231642 152720
rect 240318 152668 240324 152720
rect 240376 152708 240382 152720
rect 241882 152708 241888 152720
rect 240376 152680 241888 152708
rect 240376 152668 240382 152680
rect 241882 152668 241888 152680
rect 241940 152668 241946 152720
rect 251174 152668 251180 152720
rect 251232 152708 251238 152720
rect 311158 152708 311164 152720
rect 251232 152680 311164 152708
rect 251232 152668 251238 152680
rect 311158 152668 311164 152680
rect 311216 152668 311222 152720
rect 312170 152668 312176 152720
rect 312228 152708 312234 152720
rect 356146 152708 356152 152720
rect 312228 152680 356152 152708
rect 312228 152668 312234 152680
rect 356146 152668 356152 152680
rect 356204 152668 356210 152720
rect 358814 152668 358820 152720
rect 358872 152708 358878 152720
rect 393406 152708 393412 152720
rect 358872 152680 393412 152708
rect 358872 152668 358878 152680
rect 393406 152668 393412 152680
rect 393464 152668 393470 152720
rect 393498 152668 393504 152720
rect 393556 152708 393562 152720
rect 398098 152708 398104 152720
rect 393556 152680 398104 152708
rect 393556 152668 393562 152680
rect 398098 152668 398104 152680
rect 398156 152668 398162 152720
rect 399202 152668 399208 152720
rect 399260 152708 399266 152720
rect 417326 152708 417332 152720
rect 399260 152680 417332 152708
rect 399260 152668 399266 152680
rect 417326 152668 417332 152680
rect 417384 152668 417390 152720
rect 421650 152708 421656 152720
rect 417436 152680 421656 152708
rect 22186 152600 22192 152652
rect 22244 152640 22250 152652
rect 135898 152640 135904 152652
rect 22244 152612 135904 152640
rect 22244 152600 22250 152612
rect 135898 152600 135904 152612
rect 135956 152600 135962 152652
rect 151906 152640 151912 152652
rect 137986 152612 151912 152640
rect 19334 152532 19340 152584
rect 19392 152572 19398 152584
rect 133966 152572 133972 152584
rect 19392 152544 133972 152572
rect 19392 152532 19398 152544
rect 133966 152532 133972 152544
rect 134024 152532 134030 152584
rect 136634 152532 136640 152584
rect 136692 152572 136698 152584
rect 137986 152572 138014 152612
rect 151906 152600 151912 152612
rect 151964 152600 151970 152652
rect 153562 152600 153568 152652
rect 153620 152640 153626 152652
rect 236730 152640 236736 152652
rect 153620 152612 236736 152640
rect 153620 152600 153626 152612
rect 236730 152600 236736 152612
rect 236788 152600 236794 152652
rect 247034 152600 247040 152652
rect 247092 152640 247098 152652
rect 307938 152640 307944 152652
rect 247092 152612 307944 152640
rect 247092 152600 247098 152612
rect 307938 152600 307944 152612
rect 307996 152600 308002 152652
rect 311526 152600 311532 152652
rect 311584 152640 311590 152652
rect 320818 152640 320824 152652
rect 311584 152612 320824 152640
rect 311584 152600 311590 152612
rect 320818 152600 320824 152612
rect 320876 152600 320882 152652
rect 320910 152600 320916 152652
rect 320968 152640 320974 152652
rect 361942 152640 361948 152652
rect 320968 152612 361948 152640
rect 320968 152600 320974 152612
rect 361942 152600 361948 152612
rect 362000 152600 362006 152652
rect 368474 152600 368480 152652
rect 368532 152640 368538 152652
rect 400398 152640 400404 152652
rect 368532 152612 400404 152640
rect 368532 152600 368538 152612
rect 400398 152600 400404 152612
rect 400456 152600 400462 152652
rect 413922 152640 413928 152652
rect 403452 152612 413928 152640
rect 136692 152544 138014 152572
rect 136692 152532 136698 152544
rect 138106 152532 138112 152584
rect 138164 152572 138170 152584
rect 144270 152572 144276 152584
rect 138164 152544 144276 152572
rect 138164 152532 138170 152544
rect 144270 152532 144276 152544
rect 144328 152532 144334 152584
rect 144362 152532 144368 152584
rect 144420 152572 144426 152584
rect 226426 152572 226432 152584
rect 144420 152544 226432 152572
rect 144420 152532 144426 152544
rect 226426 152532 226432 152544
rect 226484 152532 226490 152584
rect 234154 152532 234160 152584
rect 234212 152572 234218 152584
rect 297726 152572 297732 152584
rect 234212 152544 297732 152572
rect 234212 152532 234218 152544
rect 297726 152532 297732 152544
rect 297784 152532 297790 152584
rect 303614 152532 303620 152584
rect 303672 152572 303678 152584
rect 350994 152572 351000 152584
rect 303672 152544 351000 152572
rect 303672 152532 303678 152544
rect 350994 152532 351000 152544
rect 351052 152532 351058 152584
rect 351914 152532 351920 152584
rect 351972 152572 351978 152584
rect 353478 152572 353484 152584
rect 351972 152544 353484 152572
rect 351972 152532 351978 152544
rect 353478 152532 353484 152544
rect 353536 152532 353542 152584
rect 354490 152532 354496 152584
rect 354548 152572 354554 152584
rect 389542 152572 389548 152584
rect 354548 152544 389548 152572
rect 354548 152532 354554 152544
rect 389542 152532 389548 152544
rect 389600 152532 389606 152584
rect 390370 152532 390376 152584
rect 390428 152572 390434 152584
rect 397914 152572 397920 152584
rect 390428 152544 397920 152572
rect 390428 152532 390434 152544
rect 397914 152532 397920 152544
rect 397972 152532 397978 152584
rect 398006 152532 398012 152584
rect 398064 152572 398070 152584
rect 403342 152572 403348 152584
rect 398064 152544 403348 152572
rect 398064 152532 398070 152544
rect 403342 152532 403348 152544
rect 403400 152532 403406 152584
rect 2866 152464 2872 152516
rect 2924 152504 2930 152516
rect 121086 152504 121092 152516
rect 2924 152476 121092 152504
rect 2924 152464 2930 152476
rect 121086 152464 121092 152476
rect 121144 152464 121150 152516
rect 126974 152464 126980 152516
rect 127032 152504 127038 152516
rect 216122 152504 216128 152516
rect 127032 152476 216128 152504
rect 127032 152464 127038 152476
rect 216122 152464 216128 152476
rect 216180 152464 216186 152516
rect 227714 152464 227720 152516
rect 227772 152504 227778 152516
rect 293218 152504 293224 152516
rect 227772 152476 293224 152504
rect 227772 152464 227778 152476
rect 293218 152464 293224 152476
rect 293276 152464 293282 152516
rect 298646 152464 298652 152516
rect 298704 152504 298710 152516
rect 347130 152504 347136 152516
rect 298704 152476 347136 152504
rect 298704 152464 298710 152476
rect 347130 152464 347136 152476
rect 347188 152464 347194 152516
rect 348142 152464 348148 152516
rect 348200 152504 348206 152516
rect 385034 152504 385040 152516
rect 348200 152476 385040 152504
rect 348200 152464 348206 152476
rect 385034 152464 385040 152476
rect 385092 152464 385098 152516
rect 386414 152464 386420 152516
rect 386472 152504 386478 152516
rect 403452 152504 403480 152612
rect 413922 152600 413928 152612
rect 413980 152600 413986 152652
rect 414014 152600 414020 152652
rect 414072 152640 414078 152652
rect 417436 152640 417464 152680
rect 421650 152668 421656 152680
rect 421708 152668 421714 152720
rect 426342 152708 426348 152720
rect 421852 152680 426348 152708
rect 414072 152612 417464 152640
rect 414072 152600 414078 152612
rect 417602 152600 417608 152652
rect 417660 152640 417666 152652
rect 421742 152640 421748 152652
rect 417660 152612 421748 152640
rect 417660 152600 417666 152612
rect 421742 152600 421748 152612
rect 421800 152600 421806 152652
rect 403526 152532 403532 152584
rect 403584 152572 403590 152584
rect 419074 152572 419080 152584
rect 403584 152544 419080 152572
rect 403584 152532 403590 152544
rect 419074 152532 419080 152544
rect 419132 152532 419138 152584
rect 421852 152572 421880 152680
rect 426342 152668 426348 152680
rect 426400 152668 426406 152720
rect 426434 152668 426440 152720
rect 426492 152708 426498 152720
rect 444742 152708 444748 152720
rect 426492 152680 444748 152708
rect 426492 152668 426498 152680
rect 444742 152668 444748 152680
rect 444800 152668 444806 152720
rect 444852 152708 444880 152748
rect 444926 152736 444932 152788
rect 444984 152776 444990 152788
rect 451182 152776 451188 152788
rect 444984 152748 451188 152776
rect 444984 152736 444990 152748
rect 451182 152736 451188 152748
rect 451240 152736 451246 152788
rect 458174 152708 458180 152720
rect 444852 152680 458180 152708
rect 458174 152668 458180 152680
rect 458232 152668 458238 152720
rect 421926 152600 421932 152652
rect 421984 152640 421990 152652
rect 429194 152640 429200 152652
rect 421984 152612 426204 152640
rect 421984 152600 421990 152612
rect 426066 152572 426072 152584
rect 419184 152544 421880 152572
rect 422128 152544 426072 152572
rect 410058 152504 410064 152516
rect 386472 152476 403480 152504
rect 403636 152476 410064 152504
rect 386472 152464 386478 152476
rect 66622 152396 66628 152448
rect 66680 152436 66686 152448
rect 159634 152436 159640 152448
rect 66680 152408 159640 152436
rect 66680 152396 66686 152408
rect 159634 152396 159640 152408
rect 159692 152396 159698 152448
rect 173158 152396 173164 152448
rect 173216 152436 173222 152448
rect 249518 152436 249524 152448
rect 173216 152408 249524 152436
rect 173216 152396 173222 152408
rect 249518 152396 249524 152408
rect 249576 152396 249582 152448
rect 260926 152396 260932 152448
rect 260984 152436 260990 152448
rect 316310 152436 316316 152448
rect 260984 152408 316316 152436
rect 260984 152396 260990 152408
rect 316310 152396 316316 152408
rect 316368 152396 316374 152448
rect 317506 152396 317512 152448
rect 317564 152436 317570 152448
rect 320634 152436 320640 152448
rect 317564 152408 320640 152436
rect 317564 152396 317570 152408
rect 320634 152396 320640 152408
rect 320692 152396 320698 152448
rect 320726 152396 320732 152448
rect 320784 152436 320790 152448
rect 325970 152436 325976 152448
rect 320784 152408 325976 152436
rect 320784 152396 320790 152408
rect 325970 152396 325976 152408
rect 326028 152396 326034 152448
rect 326062 152396 326068 152448
rect 326120 152436 326126 152448
rect 367646 152436 367652 152448
rect 326120 152408 367652 152436
rect 326120 152396 326126 152408
rect 367646 152396 367652 152408
rect 367704 152396 367710 152448
rect 380986 152396 380992 152448
rect 381044 152436 381050 152448
rect 403636 152436 403664 152476
rect 410058 152464 410064 152476
rect 410116 152464 410122 152516
rect 413830 152464 413836 152516
rect 413888 152504 413894 152516
rect 416498 152504 416504 152516
rect 413888 152476 416504 152504
rect 413888 152464 413894 152476
rect 416498 152464 416504 152476
rect 416556 152464 416562 152516
rect 418614 152464 418620 152516
rect 418672 152504 418678 152516
rect 419184 152504 419212 152544
rect 418672 152476 419212 152504
rect 418672 152464 418678 152476
rect 419534 152464 419540 152516
rect 419592 152504 419598 152516
rect 421926 152504 421932 152516
rect 419592 152476 421932 152504
rect 419592 152464 419598 152476
rect 421926 152464 421932 152476
rect 421984 152464 421990 152516
rect 381044 152408 403664 152436
rect 381044 152396 381050 152408
rect 403710 152396 403716 152448
rect 403768 152436 403774 152448
rect 412634 152436 412640 152448
rect 403768 152408 412640 152436
rect 403768 152396 403774 152408
rect 412634 152396 412640 152408
rect 412692 152396 412698 152448
rect 415302 152396 415308 152448
rect 415360 152436 415366 152448
rect 420362 152436 420368 152448
rect 415360 152408 420368 152436
rect 415360 152396 415366 152408
rect 420362 152396 420368 152408
rect 420420 152396 420426 152448
rect 33594 152328 33600 152380
rect 33652 152368 33658 152380
rect 109678 152368 109684 152380
rect 33652 152340 109684 152368
rect 33652 152328 33658 152340
rect 109678 152328 109684 152340
rect 109736 152328 109742 152380
rect 109770 152328 109776 152380
rect 109828 152368 109834 152380
rect 110506 152368 110512 152380
rect 109828 152340 110512 152368
rect 109828 152328 109834 152340
rect 110506 152328 110512 152340
rect 110564 152328 110570 152380
rect 120074 152328 120080 152380
rect 120132 152368 120138 152380
rect 211062 152368 211068 152380
rect 120132 152340 211068 152368
rect 120132 152328 120138 152340
rect 211062 152328 211068 152340
rect 211120 152328 211126 152380
rect 224402 152328 224408 152380
rect 224460 152368 224466 152380
rect 288066 152368 288072 152380
rect 224460 152340 288072 152368
rect 224460 152328 224466 152340
rect 288066 152328 288072 152340
rect 288124 152328 288130 152380
rect 291378 152328 291384 152380
rect 291436 152368 291442 152380
rect 341334 152368 341340 152380
rect 291436 152340 341340 152368
rect 291436 152328 291442 152340
rect 341334 152328 341340 152340
rect 341392 152328 341398 152380
rect 343818 152328 343824 152380
rect 343876 152368 343882 152380
rect 349798 152368 349804 152380
rect 343876 152340 349804 152368
rect 343876 152328 343882 152340
rect 349798 152328 349804 152340
rect 349856 152328 349862 152380
rect 349890 152328 349896 152380
rect 349948 152368 349954 152380
rect 385678 152368 385684 152380
rect 349948 152340 385684 152368
rect 349948 152328 349954 152340
rect 385678 152328 385684 152340
rect 385736 152328 385742 152380
rect 386230 152328 386236 152380
rect 386288 152368 386294 152380
rect 399754 152368 399760 152380
rect 386288 152340 399760 152368
rect 386288 152328 386294 152340
rect 399754 152328 399760 152340
rect 399812 152328 399818 152380
rect 402422 152328 402428 152380
rect 402480 152368 402486 152380
rect 422128 152368 422156 152544
rect 426066 152532 426072 152544
rect 426124 152532 426130 152584
rect 426176 152572 426204 152612
rect 426452 152612 429200 152640
rect 426452 152572 426480 152612
rect 429194 152600 429200 152612
rect 429252 152600 429258 152652
rect 429378 152600 429384 152652
rect 429436 152640 429442 152652
rect 429436 152612 441614 152640
rect 429436 152600 429442 152612
rect 426176 152544 426480 152572
rect 426526 152532 426532 152584
rect 426584 152572 426590 152584
rect 438946 152572 438952 152584
rect 426584 152544 438952 152572
rect 426584 152532 426590 152544
rect 438946 152532 438952 152544
rect 439004 152532 439010 152584
rect 439038 152532 439044 152584
rect 439096 152572 439102 152584
rect 440878 152572 440884 152584
rect 439096 152544 440884 152572
rect 439096 152532 439102 152544
rect 440878 152532 440884 152544
rect 440936 152532 440942 152584
rect 441586 152572 441614 152612
rect 441982 152600 441988 152652
rect 442040 152640 442046 152652
rect 446122 152640 446128 152652
rect 442040 152612 446128 152640
rect 442040 152600 442046 152612
rect 446122 152600 446128 152612
rect 446180 152600 446186 152652
rect 446398 152600 446404 152652
rect 446456 152640 446462 152652
rect 453758 152640 453764 152652
rect 446456 152612 453764 152640
rect 446456 152600 446462 152612
rect 453758 152600 453764 152612
rect 453816 152600 453822 152652
rect 447318 152572 447324 152584
rect 441586 152544 447324 152572
rect 447318 152532 447324 152544
rect 447376 152532 447382 152584
rect 447410 152532 447416 152584
rect 447468 152572 447474 152584
rect 456978 152572 456984 152584
rect 447468 152544 456984 152572
rect 447468 152532 447474 152544
rect 456978 152532 456984 152544
rect 457036 152532 457042 152584
rect 422846 152464 422852 152516
rect 422904 152504 422910 152516
rect 435726 152504 435732 152516
rect 422904 152476 435732 152504
rect 422904 152464 422910 152476
rect 435726 152464 435732 152476
rect 435784 152464 435790 152516
rect 436922 152464 436928 152516
rect 436980 152504 436986 152516
rect 446766 152504 446772 152516
rect 436980 152476 446772 152504
rect 436980 152464 436986 152476
rect 446766 152464 446772 152476
rect 446824 152464 446830 152516
rect 459554 152464 459560 152516
rect 459612 152504 459618 152516
rect 464614 152504 464620 152516
rect 459612 152476 464620 152504
rect 459612 152464 459618 152476
rect 464614 152464 464620 152476
rect 464672 152464 464678 152516
rect 422202 152396 422208 152448
rect 422260 152436 422266 152448
rect 422260 152408 422892 152436
rect 422260 152396 422266 152408
rect 402480 152340 422156 152368
rect 422864 152368 422892 152408
rect 423030 152396 423036 152448
rect 423088 152436 423094 152448
rect 442166 152436 442172 152448
rect 423088 152408 442172 152436
rect 423088 152396 423094 152408
rect 442166 152396 442172 152408
rect 442224 152396 442230 152448
rect 442994 152396 443000 152448
rect 443052 152436 443058 152448
rect 457622 152436 457628 152448
rect 443052 152408 457628 152436
rect 443052 152396 443058 152408
rect 457622 152396 457628 152408
rect 457680 152396 457686 152448
rect 424410 152368 424416 152380
rect 422864 152340 424416 152368
rect 402480 152328 402486 152340
rect 424410 152328 424416 152340
rect 424468 152328 424474 152380
rect 424502 152328 424508 152380
rect 424560 152368 424566 152380
rect 426894 152368 426900 152380
rect 424560 152340 426900 152368
rect 424560 152328 424566 152340
rect 426894 152328 426900 152340
rect 426952 152328 426958 152380
rect 427814 152328 427820 152380
rect 427872 152368 427878 152380
rect 446030 152368 446036 152380
rect 427872 152340 446036 152368
rect 427872 152328 427878 152340
rect 446030 152328 446036 152340
rect 446088 152328 446094 152380
rect 446122 152328 446128 152380
rect 446180 152368 446186 152380
rect 449250 152368 449256 152380
rect 446180 152340 449256 152368
rect 446180 152328 446186 152340
rect 449250 152328 449256 152340
rect 449308 152328 449314 152380
rect 91094 152260 91100 152312
rect 91152 152300 91158 152312
rect 180242 152300 180248 152312
rect 91152 152272 180248 152300
rect 91152 152260 91158 152272
rect 180242 152260 180248 152272
rect 180300 152260 180306 152312
rect 187970 152260 187976 152312
rect 188028 152300 188034 152312
rect 262398 152300 262404 152312
rect 188028 152272 262404 152300
rect 188028 152260 188034 152272
rect 262398 152260 262404 152272
rect 262456 152260 262462 152312
rect 266354 152260 266360 152312
rect 266412 152300 266418 152312
rect 320910 152300 320916 152312
rect 266412 152272 320916 152300
rect 266412 152260 266418 152272
rect 320910 152260 320916 152272
rect 320968 152260 320974 152312
rect 331214 152260 331220 152312
rect 331272 152300 331278 152312
rect 372154 152300 372160 152312
rect 331272 152272 372160 152300
rect 331272 152260 331278 152272
rect 372154 152260 372160 152272
rect 372212 152260 372218 152312
rect 382274 152260 382280 152312
rect 382332 152300 382338 152312
rect 386966 152300 386972 152312
rect 382332 152272 386972 152300
rect 382332 152260 382338 152272
rect 386966 152260 386972 152272
rect 387024 152260 387030 152312
rect 393130 152260 393136 152312
rect 393188 152300 393194 152312
rect 398006 152300 398012 152312
rect 393188 152272 398012 152300
rect 393188 152260 393194 152272
rect 398006 152260 398012 152272
rect 398064 152260 398070 152312
rect 398098 152260 398104 152312
rect 398156 152300 398162 152312
rect 403710 152300 403716 152312
rect 398156 152272 403716 152300
rect 398156 152260 398162 152272
rect 403710 152260 403716 152272
rect 403768 152260 403774 152312
rect 403802 152260 403808 152312
rect 403860 152300 403866 152312
rect 413278 152300 413284 152312
rect 403860 152272 413284 152300
rect 403860 152260 403866 152272
rect 413278 152260 413284 152272
rect 413336 152260 413342 152312
rect 414290 152260 414296 152312
rect 414348 152300 414354 152312
rect 422846 152300 422852 152312
rect 414348 152272 422852 152300
rect 414348 152260 414354 152272
rect 422846 152260 422852 152272
rect 422904 152260 422910 152312
rect 423122 152260 423128 152312
rect 423180 152300 423186 152312
rect 441522 152300 441528 152312
rect 423180 152272 441528 152300
rect 423180 152260 423186 152272
rect 441522 152260 441528 152272
rect 441580 152260 441586 152312
rect 441614 152260 441620 152312
rect 441672 152300 441678 152312
rect 456334 152300 456340 152312
rect 441672 152272 456340 152300
rect 441672 152260 441678 152272
rect 456334 152260 456340 152272
rect 456392 152260 456398 152312
rect 19794 152192 19800 152244
rect 19852 152232 19858 152244
rect 97902 152232 97908 152244
rect 19852 152204 97908 152232
rect 19852 152192 19858 152204
rect 97902 152192 97908 152204
rect 97960 152192 97966 152244
rect 109034 152192 109040 152244
rect 109092 152232 109098 152244
rect 130746 152232 130752 152244
rect 109092 152204 130752 152232
rect 109092 152192 109098 152204
rect 130746 152192 130752 152204
rect 130804 152192 130810 152244
rect 134058 152192 134064 152244
rect 134116 152232 134122 152244
rect 221274 152232 221280 152244
rect 134116 152204 221280 152232
rect 134116 152192 134122 152204
rect 221274 152192 221280 152204
rect 221332 152192 221338 152244
rect 222102 152192 222108 152244
rect 222160 152232 222166 152244
rect 282914 152232 282920 152244
rect 222160 152204 282920 152232
rect 222160 152192 222166 152204
rect 282914 152192 282920 152204
rect 282972 152192 282978 152244
rect 285766 152192 285772 152244
rect 285824 152232 285830 152244
rect 336182 152232 336188 152244
rect 285824 152204 336188 152232
rect 285824 152192 285830 152204
rect 336182 152192 336188 152204
rect 336240 152192 336246 152244
rect 342438 152192 342444 152244
rect 342496 152232 342502 152244
rect 344554 152232 344560 152244
rect 342496 152204 344560 152232
rect 342496 152192 342502 152204
rect 344554 152192 344560 152204
rect 344612 152192 344618 152244
rect 349154 152192 349160 152244
rect 349212 152232 349218 152244
rect 349890 152232 349896 152244
rect 349212 152204 349896 152232
rect 349212 152192 349218 152204
rect 349890 152192 349896 152204
rect 349948 152192 349954 152244
rect 352006 152192 352012 152244
rect 352064 152232 352070 152244
rect 388254 152232 388260 152244
rect 352064 152204 388260 152232
rect 352064 152192 352070 152204
rect 388254 152192 388260 152204
rect 388312 152192 388318 152244
rect 394326 152192 394332 152244
rect 394384 152232 394390 152244
rect 417786 152232 417792 152244
rect 394384 152204 417792 152232
rect 394384 152192 394390 152204
rect 417786 152192 417792 152204
rect 417844 152192 417850 152244
rect 417878 152192 417884 152244
rect 417936 152232 417942 152244
rect 424318 152232 424324 152244
rect 417936 152204 424324 152232
rect 417936 152192 417942 152204
rect 424318 152192 424324 152204
rect 424376 152192 424382 152244
rect 425974 152192 425980 152244
rect 426032 152232 426038 152244
rect 444098 152232 444104 152244
rect 426032 152204 444104 152232
rect 426032 152192 426038 152204
rect 444098 152192 444104 152204
rect 444156 152192 444162 152244
rect 445294 152192 445300 152244
rect 445352 152232 445358 152244
rect 458818 152232 458824 152244
rect 445352 152204 458824 152232
rect 445352 152192 445358 152204
rect 458818 152192 458824 152204
rect 458876 152192 458882 152244
rect 9490 152124 9496 152176
rect 9548 152164 9554 152176
rect 82814 152164 82820 152176
rect 9548 152136 82820 152164
rect 9548 152124 9554 152136
rect 82814 152124 82820 152136
rect 82872 152124 82878 152176
rect 82906 152124 82912 152176
rect 82964 152164 82970 152176
rect 169938 152164 169944 152176
rect 82964 152136 169944 152164
rect 82964 152124 82970 152136
rect 169938 152124 169944 152136
rect 169996 152124 170002 152176
rect 172146 152124 172152 152176
rect 172204 152164 172210 152176
rect 190454 152164 190460 152176
rect 172204 152136 190460 152164
rect 172204 152124 172210 152136
rect 190454 152124 190460 152136
rect 190512 152124 190518 152176
rect 193582 152124 193588 152176
rect 193640 152164 193646 152176
rect 213546 152164 213552 152176
rect 193640 152136 213552 152164
rect 193640 152124 193646 152136
rect 213546 152124 213552 152136
rect 213604 152124 213610 152176
rect 225322 152124 225328 152176
rect 225380 152164 225386 152176
rect 229002 152164 229008 152176
rect 225380 152136 229008 152164
rect 225380 152124 225386 152136
rect 229002 152124 229008 152136
rect 229060 152124 229066 152176
rect 244458 152124 244464 152176
rect 244516 152164 244522 152176
rect 306006 152164 306012 152176
rect 244516 152136 306012 152164
rect 244516 152124 244522 152136
rect 306006 152124 306012 152136
rect 306064 152124 306070 152176
rect 320818 152124 320824 152176
rect 320876 152164 320882 152176
rect 356790 152164 356796 152176
rect 320876 152136 356796 152164
rect 320876 152124 320882 152136
rect 356790 152124 356796 152136
rect 356848 152124 356854 152176
rect 357526 152124 357532 152176
rect 357584 152164 357590 152176
rect 359366 152164 359372 152176
rect 357584 152136 359372 152164
rect 357584 152124 357590 152136
rect 359366 152124 359372 152136
rect 359424 152124 359430 152176
rect 365714 152124 365720 152176
rect 365772 152164 365778 152176
rect 398466 152164 398472 152176
rect 365772 152136 398472 152164
rect 365772 152124 365778 152136
rect 398466 152124 398472 152136
rect 398524 152124 398530 152176
rect 398558 152124 398564 152176
rect 398616 152164 398622 152176
rect 408126 152164 408132 152176
rect 398616 152136 408132 152164
rect 398616 152124 398622 152136
rect 408126 152124 408132 152136
rect 408184 152124 408190 152176
rect 409230 152124 409236 152176
rect 409288 152164 409294 152176
rect 428642 152164 428648 152176
rect 409288 152136 428648 152164
rect 409288 152124 409294 152136
rect 428642 152124 428648 152136
rect 428700 152124 428706 152176
rect 430666 152124 430672 152176
rect 430724 152164 430730 152176
rect 447962 152164 447968 152176
rect 430724 152136 447968 152164
rect 430724 152124 430730 152136
rect 447962 152124 447968 152136
rect 448020 152124 448026 152176
rect 79318 152056 79324 152108
rect 79376 152096 79382 152108
rect 164786 152096 164792 152108
rect 79376 152068 164792 152096
rect 79376 152056 79382 152068
rect 164786 152056 164792 152068
rect 164844 152056 164850 152108
rect 166994 152056 167000 152108
rect 167052 152096 167058 152108
rect 182726 152096 182732 152108
rect 167052 152068 182732 152096
rect 167052 152056 167058 152068
rect 182726 152056 182732 152068
rect 182784 152056 182790 152108
rect 183462 152056 183468 152108
rect 183520 152096 183526 152108
rect 200758 152096 200764 152108
rect 183520 152068 200764 152096
rect 183520 152056 183526 152068
rect 200758 152056 200764 152068
rect 200816 152056 200822 152108
rect 213822 152056 213828 152108
rect 213880 152096 213886 152108
rect 274542 152096 274548 152108
rect 213880 152068 274548 152096
rect 213880 152056 213886 152068
rect 274542 152056 274548 152068
rect 274600 152056 274606 152108
rect 277394 152056 277400 152108
rect 277452 152096 277458 152108
rect 331122 152096 331128 152108
rect 277452 152068 331128 152096
rect 277452 152056 277458 152068
rect 331122 152056 331128 152068
rect 331180 152056 331186 152108
rect 335354 152056 335360 152108
rect 335412 152096 335418 152108
rect 375374 152096 375380 152108
rect 335412 152068 375380 152096
rect 335412 152056 335418 152068
rect 375374 152056 375380 152068
rect 375432 152056 375438 152108
rect 378778 152056 378784 152108
rect 378836 152096 378842 152108
rect 384390 152096 384396 152108
rect 378836 152068 384396 152096
rect 378836 152056 378842 152068
rect 384390 152056 384396 152068
rect 384448 152056 384454 152108
rect 388438 152056 388444 152108
rect 388496 152096 388502 152108
rect 407482 152096 407488 152108
rect 388496 152068 407488 152096
rect 388496 152056 388502 152068
rect 407482 152056 407488 152068
rect 407540 152056 407546 152108
rect 408494 152056 408500 152108
rect 408552 152096 408558 152108
rect 423582 152096 423588 152108
rect 408552 152068 423588 152096
rect 408552 152056 408558 152068
rect 423582 152056 423588 152068
rect 423640 152056 423646 152108
rect 424410 152056 424416 152108
rect 424468 152096 424474 152108
rect 433794 152096 433800 152108
rect 424468 152068 433800 152096
rect 424468 152056 424474 152068
rect 433794 152056 433800 152068
rect 433852 152056 433858 152108
rect 433886 152056 433892 152108
rect 433944 152096 433950 152108
rect 449894 152096 449900 152108
rect 433944 152068 449900 152096
rect 433944 152056 433950 152068
rect 449894 152056 449900 152068
rect 449952 152056 449958 152108
rect 516686 152056 516692 152108
rect 516744 152096 516750 152108
rect 520274 152096 520280 152108
rect 516744 152068 520280 152096
rect 516744 152056 516750 152068
rect 520274 152056 520280 152068
rect 520332 152056 520338 152108
rect 68922 151988 68928 152040
rect 68980 152028 68986 152040
rect 142798 152028 142804 152040
rect 68980 152000 142804 152028
rect 68980 151988 68986 152000
rect 142798 151988 142804 152000
rect 142856 151988 142862 152040
rect 143166 151988 143172 152040
rect 143224 152028 143230 152040
rect 146938 152028 146944 152040
rect 143224 152000 146944 152028
rect 143224 151988 143230 152000
rect 146938 151988 146944 152000
rect 146996 151988 147002 152040
rect 156322 151988 156328 152040
rect 156380 152028 156386 152040
rect 172514 152028 172520 152040
rect 156380 152000 172520 152028
rect 156380 151988 156386 152000
rect 172514 151988 172520 152000
rect 172572 151988 172578 152040
rect 191466 151988 191472 152040
rect 191524 152028 191530 152040
rect 208486 152028 208492 152040
rect 191524 152000 208492 152028
rect 191524 151988 191530 152000
rect 208486 151988 208492 152000
rect 208544 151988 208550 152040
rect 242434 151988 242440 152040
rect 242492 152028 242498 152040
rect 300946 152028 300952 152040
rect 242492 152000 300952 152028
rect 242492 151988 242498 152000
rect 300946 151988 300952 152000
rect 301004 151988 301010 152040
rect 304166 151988 304172 152040
rect 304224 152028 304230 152040
rect 351638 152028 351644 152040
rect 304224 152000 351644 152028
rect 304224 151988 304230 152000
rect 351638 151988 351644 152000
rect 351696 151988 351702 152040
rect 354674 151988 354680 152040
rect 354732 152028 354738 152040
rect 390186 152028 390192 152040
rect 354732 152000 390192 152028
rect 354732 151988 354738 152000
rect 390186 151988 390192 152000
rect 390244 151988 390250 152040
rect 397178 152028 397184 152040
rect 393424 152000 397184 152028
rect 75086 151920 75092 151972
rect 75144 151960 75150 151972
rect 154482 151960 154488 151972
rect 75144 151932 154488 151960
rect 75144 151920 75150 151932
rect 154482 151920 154488 151932
rect 154540 151920 154546 151972
rect 162486 151920 162492 151972
rect 162544 151960 162550 151972
rect 177666 151960 177672 151972
rect 162544 151932 177672 151960
rect 162544 151920 162550 151932
rect 177666 151920 177672 151932
rect 177724 151920 177730 151972
rect 184382 151920 184388 151972
rect 184440 151960 184446 151972
rect 195606 151960 195612 151972
rect 184440 151932 195612 151960
rect 184440 151920 184446 151932
rect 195606 151920 195612 151932
rect 195664 151920 195670 151972
rect 243354 151920 243360 151972
rect 243412 151960 243418 151972
rect 302878 151960 302884 151972
rect 243412 151932 302884 151960
rect 243412 151920 243418 151932
rect 302878 151920 302884 151932
rect 302936 151920 302942 151972
rect 307662 151920 307668 151972
rect 307720 151960 307726 151972
rect 352282 151960 352288 151972
rect 307720 151932 352288 151960
rect 307720 151920 307726 151932
rect 352282 151920 352288 151932
rect 352340 151920 352346 151972
rect 364610 151920 364616 151972
rect 364668 151960 364674 151972
rect 393424 151960 393452 152000
rect 397178 151988 397184 152000
rect 397236 151988 397242 152040
rect 404906 152028 404912 152040
rect 398806 152000 404912 152028
rect 398806 151960 398834 152000
rect 404906 151988 404912 152000
rect 404964 151988 404970 152040
rect 405366 151988 405372 152040
rect 405424 152028 405430 152040
rect 421006 152028 421012 152040
rect 405424 152000 421012 152028
rect 405424 151988 405430 152000
rect 421006 151988 421012 152000
rect 421064 151988 421070 152040
rect 434438 152028 434444 152040
rect 421116 152000 434444 152028
rect 364668 151932 393452 151960
rect 393976 151932 398834 151960
rect 364668 151920 364674 151932
rect 30190 151852 30196 151904
rect 30248 151892 30254 151904
rect 110322 151892 110328 151904
rect 30248 151864 110328 151892
rect 30248 151852 30254 151864
rect 110322 151852 110328 151864
rect 110380 151852 110386 151904
rect 110506 151852 110512 151904
rect 110564 151892 110570 151904
rect 138474 151892 138480 151904
rect 110564 151864 138480 151892
rect 110564 151852 110570 151864
rect 138474 151852 138480 151864
rect 138532 151852 138538 151904
rect 139302 151852 139308 151904
rect 139360 151892 139366 151904
rect 203334 151892 203340 151904
rect 139360 151864 203340 151892
rect 139360 151852 139366 151864
rect 203334 151852 203340 151864
rect 203392 151852 203398 151904
rect 212626 151852 212632 151904
rect 212684 151892 212690 151904
rect 272702 151892 272708 151904
rect 212684 151864 272708 151892
rect 212684 151852 212690 151864
rect 272702 151852 272708 151864
rect 272760 151852 272766 151904
rect 320726 151892 320732 151904
rect 277366 151864 320732 151892
rect 74810 151784 74816 151836
rect 74868 151824 74874 151836
rect 81342 151824 81348 151836
rect 74868 151796 81348 151824
rect 74868 151784 74874 151796
rect 81342 151784 81348 151796
rect 81400 151784 81406 151836
rect 105814 151784 105820 151836
rect 105872 151824 105878 151836
rect 110230 151824 110236 151836
rect 105872 151796 110236 151824
rect 105872 151784 105878 151796
rect 110230 151784 110236 151796
rect 110288 151784 110294 151836
rect 110414 151784 110420 151836
rect 110472 151824 110478 151836
rect 128170 151824 128176 151836
rect 110472 151796 128176 151824
rect 110472 151784 110478 151796
rect 128170 151784 128176 151796
rect 128228 151784 128234 151836
rect 129734 151784 129740 151836
rect 129792 151824 129798 151836
rect 146846 151824 146852 151836
rect 129792 151796 146852 151824
rect 129792 151784 129798 151796
rect 146846 151784 146852 151796
rect 146904 151784 146910 151836
rect 146938 151784 146944 151836
rect 146996 151824 147002 151836
rect 157058 151824 157064 151836
rect 146996 151796 157064 151824
rect 146996 151784 147002 151796
rect 157058 151784 157064 151796
rect 157116 151784 157122 151836
rect 169754 151784 169760 151836
rect 169812 151824 169818 151836
rect 185302 151824 185308 151836
rect 169812 151796 185308 151824
rect 169812 151784 169818 151796
rect 185302 151784 185308 151796
rect 185360 151784 185366 151836
rect 271874 151784 271880 151836
rect 271932 151824 271938 151836
rect 277366 151824 277394 151864
rect 320726 151852 320732 151864
rect 320784 151852 320790 151904
rect 321554 151852 321560 151904
rect 321612 151892 321618 151904
rect 362586 151892 362592 151904
rect 321612 151864 362592 151892
rect 321612 151852 321618 151864
rect 362586 151852 362592 151864
rect 362644 151852 362650 151904
rect 363138 151852 363144 151904
rect 363196 151892 363202 151904
rect 364518 151892 364524 151904
rect 363196 151864 364524 151892
rect 363196 151852 363202 151864
rect 364518 151852 364524 151864
rect 364576 151852 364582 151904
rect 388162 151852 388168 151904
rect 388220 151892 388226 151904
rect 393976 151892 394004 151932
rect 404170 151920 404176 151972
rect 404228 151960 404234 151972
rect 418430 151960 418436 151972
rect 404228 151932 418436 151960
rect 404228 151920 404234 151932
rect 418430 151920 418436 151932
rect 418488 151920 418494 151972
rect 419626 151920 419632 151972
rect 419684 151960 419690 151972
rect 421116 151960 421144 152000
rect 434438 151988 434444 152000
rect 434496 151988 434502 152040
rect 434622 151988 434628 152040
rect 434680 152028 434686 152040
rect 443454 152028 443460 152040
rect 434680 152000 443460 152028
rect 434680 151988 434686 152000
rect 443454 151988 443460 152000
rect 443512 151988 443518 152040
rect 446306 151988 446312 152040
rect 446364 152028 446370 152040
rect 460014 152028 460020 152040
rect 446364 152000 460020 152028
rect 446364 151988 446370 152000
rect 460014 151988 460020 152000
rect 460072 151988 460078 152040
rect 485774 151988 485780 152040
rect 485832 152028 485838 152040
rect 490282 152028 490288 152040
rect 485832 152000 490288 152028
rect 485832 151988 485838 152000
rect 490282 151988 490288 152000
rect 490340 151988 490346 152040
rect 419684 151932 421144 151960
rect 419684 151920 419690 151932
rect 423214 151920 423220 151972
rect 423272 151960 423278 151972
rect 439590 151960 439596 151972
rect 423272 151932 439596 151960
rect 423272 151920 423278 151932
rect 439590 151920 439596 151932
rect 439648 151920 439654 151972
rect 440234 151920 440240 151972
rect 440292 151960 440298 151972
rect 455046 151960 455052 151972
rect 440292 151932 455052 151960
rect 440292 151920 440298 151932
rect 455046 151920 455052 151932
rect 455104 151920 455110 151972
rect 469214 151920 469220 151972
rect 469272 151960 469278 151972
rect 472342 151960 472348 151972
rect 469272 151932 472348 151960
rect 469272 151920 469278 151932
rect 472342 151920 472348 151932
rect 472400 151920 472406 151972
rect 488534 151920 488540 151972
rect 488592 151960 488598 151972
rect 492214 151960 492220 151972
rect 488592 151932 492220 151960
rect 488592 151920 488598 151932
rect 492214 151920 492220 151932
rect 492272 151920 492278 151972
rect 509050 151920 509056 151972
rect 509108 151960 509114 151972
rect 510890 151960 510896 151972
rect 509108 151932 510896 151960
rect 509108 151920 509114 151932
rect 510890 151920 510896 151932
rect 510948 151920 510954 151972
rect 517422 151920 517428 151972
rect 517480 151960 517486 151972
rect 521562 151960 521568 151972
rect 517480 151932 521568 151960
rect 517480 151920 517486 151932
rect 521562 151920 521568 151932
rect 521620 151920 521626 151972
rect 388220 151864 394004 151892
rect 388220 151852 388226 151864
rect 396166 151852 396172 151904
rect 396224 151892 396230 151904
rect 402974 151892 402980 151904
rect 396224 151864 402980 151892
rect 396224 151852 396230 151864
rect 402974 151852 402980 151864
rect 403032 151852 403038 151904
rect 416590 151852 416596 151904
rect 416648 151892 416654 151904
rect 426802 151892 426808 151904
rect 416648 151864 426808 151892
rect 416648 151852 416654 151864
rect 426802 151852 426808 151864
rect 426860 151852 426866 151904
rect 426894 151852 426900 151904
rect 426952 151892 426958 151904
rect 437014 151892 437020 151904
rect 426952 151864 437020 151892
rect 426952 151852 426958 151864
rect 437014 151852 437020 151864
rect 437072 151852 437078 151904
rect 437474 151852 437480 151904
rect 437532 151892 437538 151904
rect 453114 151892 453120 151904
rect 437532 151864 453120 151892
rect 437532 151852 437538 151864
rect 453114 151852 453120 151864
rect 453172 151852 453178 151904
rect 468018 151852 468024 151904
rect 468076 151892 468082 151904
rect 471054 151892 471060 151904
rect 468076 151864 471060 151892
rect 468076 151852 468082 151864
rect 471054 151852 471060 151864
rect 471112 151852 471118 151904
rect 487338 151852 487344 151904
rect 487396 151892 487402 151904
rect 490926 151892 490932 151904
rect 487396 151864 490932 151892
rect 487396 151852 487402 151864
rect 490926 151852 490932 151864
rect 490984 151852 490990 151904
rect 507762 151852 507768 151904
rect 507820 151892 507826 151904
rect 509510 151892 509516 151904
rect 507820 151864 509516 151892
rect 507820 151852 507826 151864
rect 509510 151852 509516 151864
rect 509568 151852 509574 151904
rect 516042 151852 516048 151904
rect 516100 151892 516106 151904
rect 519906 151892 519912 151904
rect 516100 151864 519912 151892
rect 516100 151852 516106 151864
rect 519906 151852 519912 151864
rect 519964 151852 519970 151904
rect 271932 151796 277394 151824
rect 271932 151784 271938 151796
rect 283190 151784 283196 151836
rect 283248 151824 283254 151836
rect 287422 151824 287428 151836
rect 283248 151796 287428 151824
rect 283248 151784 283254 151796
rect 287422 151784 287428 151796
rect 287480 151784 287486 151836
rect 300394 151784 300400 151836
rect 300452 151824 300458 151836
rect 346486 151824 346492 151836
rect 300452 151796 342852 151824
rect 300452 151784 300458 151796
rect 81710 151716 81716 151768
rect 81768 151756 81774 151768
rect 112806 151756 112812 151768
rect 81768 151728 112812 151756
rect 81768 151716 81774 151728
rect 112806 151716 112812 151728
rect 112864 151716 112870 151768
rect 342824 151756 342852 151796
rect 344020 151796 346492 151824
rect 344020 151756 344048 151796
rect 346486 151784 346492 151796
rect 346544 151784 346550 151836
rect 349798 151784 349804 151836
rect 349856 151824 349862 151836
rect 380526 151824 380532 151836
rect 349856 151796 380532 151824
rect 349856 151784 349862 151796
rect 380526 151784 380532 151796
rect 380584 151784 380590 151836
rect 386138 151784 386144 151836
rect 386196 151824 386202 151836
rect 394694 151824 394700 151836
rect 386196 151796 394700 151824
rect 386196 151784 386202 151796
rect 394694 151784 394700 151796
rect 394752 151784 394758 151836
rect 404262 151784 404268 151836
rect 404320 151824 404326 151836
rect 415854 151824 415860 151836
rect 404320 151796 415860 151824
rect 404320 151784 404326 151796
rect 415854 151784 415860 151796
rect 415912 151784 415918 151836
rect 417326 151784 417332 151836
rect 417384 151824 417390 151836
rect 424226 151824 424232 151836
rect 417384 151796 424232 151824
rect 417384 151784 417390 151796
rect 424226 151784 424232 151796
rect 424284 151784 424290 151836
rect 424318 151784 424324 151836
rect 424376 151824 424382 151836
rect 431862 151824 431868 151836
rect 424376 151796 431868 151824
rect 424376 151784 424382 151796
rect 431862 151784 431868 151796
rect 431920 151784 431926 151836
rect 436094 151784 436100 151836
rect 436152 151824 436158 151836
rect 451826 151824 451832 151836
rect 436152 151796 437428 151824
rect 436152 151784 436158 151796
rect 342824 151728 344048 151756
rect 437400 151756 437428 151796
rect 438412 151796 451832 151824
rect 438412 151756 438440 151796
rect 451826 151784 451832 151796
rect 451884 151784 451890 151836
rect 467926 151784 467932 151836
rect 467984 151824 467990 151836
rect 471698 151824 471704 151836
rect 467984 151796 471704 151824
rect 467984 151784 467990 151796
rect 471698 151784 471704 151796
rect 471756 151784 471762 151836
rect 488166 151784 488172 151836
rect 488224 151824 488230 151836
rect 491570 151824 491576 151836
rect 488224 151796 491576 151824
rect 488224 151784 488230 151796
rect 491570 151784 491576 151796
rect 491628 151784 491634 151836
rect 499114 151784 499120 151836
rect 499172 151824 499178 151836
rect 499942 151824 499948 151836
rect 499172 151796 499948 151824
rect 499172 151784 499178 151796
rect 499942 151784 499948 151796
rect 500000 151784 500006 151836
rect 515490 151784 515496 151836
rect 515548 151824 515554 151836
rect 518986 151824 518992 151836
rect 515548 151796 518992 151824
rect 515548 151784 515554 151796
rect 518986 151784 518992 151796
rect 519044 151784 519050 151836
rect 437400 151728 438440 151756
rect 43898 151648 43904 151700
rect 43956 151688 43962 151700
rect 111426 151688 111432 151700
rect 43956 151660 111432 151688
rect 43956 151648 43962 151660
rect 111426 151648 111432 151660
rect 111484 151648 111490 151700
rect 40494 151580 40500 151632
rect 40552 151620 40558 151632
rect 111334 151620 111340 151632
rect 40552 151592 111340 151620
rect 40552 151580 40558 151592
rect 111334 151580 111340 151592
rect 111392 151580 111398 151632
rect 36998 151512 37004 151564
rect 37056 151552 37062 151564
rect 111058 151552 111064 151564
rect 37056 151524 111064 151552
rect 37056 151512 37062 151524
rect 111058 151512 111064 151524
rect 111116 151512 111122 151564
rect 26694 151444 26700 151496
rect 26752 151484 26758 151496
rect 116946 151484 116952 151496
rect 26752 151456 116952 151484
rect 26752 151444 26758 151456
rect 116946 151444 116952 151456
rect 117004 151444 117010 151496
rect 16390 151376 16396 151428
rect 16448 151416 16454 151428
rect 116762 151416 116768 151428
rect 16448 151388 116768 151416
rect 16448 151376 16454 151388
rect 116762 151376 116768 151388
rect 116820 151376 116826 151428
rect 12986 151308 12992 151360
rect 13044 151348 13050 151360
rect 116670 151348 116676 151360
rect 13044 151320 116676 151348
rect 13044 151308 13050 151320
rect 116670 151308 116676 151320
rect 116728 151308 116734 151360
rect 68002 151240 68008 151292
rect 68060 151280 68066 151292
rect 112714 151280 112720 151292
rect 68060 151252 112720 151280
rect 68060 151240 68066 151252
rect 112714 151240 112720 151252
rect 112772 151240 112778 151292
rect 64506 151172 64512 151224
rect 64564 151212 64570 151224
rect 112622 151212 112628 151224
rect 64564 151184 112628 151212
rect 64564 151172 64570 151184
rect 112622 151172 112628 151184
rect 112680 151172 112686 151224
rect 61102 151104 61108 151156
rect 61160 151144 61166 151156
rect 112530 151144 112536 151156
rect 61160 151116 112536 151144
rect 61160 151104 61166 151116
rect 112530 151104 112536 151116
rect 112588 151104 112594 151156
rect 57698 151036 57704 151088
rect 57756 151076 57762 151088
rect 111702 151076 111708 151088
rect 57756 151048 111708 151076
rect 57756 151036 57762 151048
rect 111702 151036 111708 151048
rect 111760 151036 111766 151088
rect 54202 150968 54208 151020
rect 54260 151008 54266 151020
rect 112438 151008 112444 151020
rect 54260 150980 112444 151008
rect 54260 150968 54266 150980
rect 112438 150968 112444 150980
rect 112496 150968 112502 151020
rect 50798 150900 50804 150952
rect 50856 150940 50862 150952
rect 111610 150940 111616 150952
rect 50856 150912 111616 150940
rect 50856 150900 50862 150912
rect 111610 150900 111616 150912
rect 111668 150900 111674 150952
rect 47302 150832 47308 150884
rect 47360 150872 47366 150884
rect 111518 150872 111524 150884
rect 47360 150844 111524 150872
rect 47360 150832 47366 150844
rect 111518 150832 111524 150844
rect 111576 150832 111582 150884
rect 98914 150764 98920 150816
rect 98972 150804 98978 150816
rect 116026 150804 116032 150816
rect 98972 150776 116032 150804
rect 98972 150764 98978 150776
rect 116026 150764 116032 150776
rect 116084 150764 116090 150816
rect 95510 150696 95516 150748
rect 95568 150736 95574 150748
rect 115290 150736 115296 150748
rect 95568 150708 115296 150736
rect 95568 150696 95574 150708
rect 115290 150696 115296 150708
rect 115348 150696 115354 150748
rect 92014 150628 92020 150680
rect 92072 150668 92078 150680
rect 113082 150668 113088 150680
rect 92072 150640 113088 150668
rect 92072 150628 92078 150640
rect 113082 150628 113088 150640
rect 113140 150628 113146 150680
rect 88610 150560 88616 150612
rect 88668 150600 88674 150612
rect 112990 150600 112996 150612
rect 88668 150572 112996 150600
rect 88668 150560 88674 150572
rect 112990 150560 112996 150572
rect 113048 150560 113054 150612
rect 85206 150492 85212 150544
rect 85264 150532 85270 150544
rect 115198 150532 115204 150544
rect 85264 150504 115204 150532
rect 85264 150492 85270 150504
rect 115198 150492 115204 150504
rect 115256 150492 115262 150544
rect 102318 150424 102324 150476
rect 102376 150464 102382 150476
rect 116118 150464 116124 150476
rect 102376 150436 116124 150464
rect 102376 150424 102382 150436
rect 116118 150424 116124 150436
rect 116176 150424 116182 150476
rect 78306 150288 78312 150340
rect 78364 150328 78370 150340
rect 112898 150328 112904 150340
rect 78364 150300 112904 150328
rect 78364 150288 78370 150300
rect 112898 150288 112904 150300
rect 112956 150288 112962 150340
rect 110322 150220 110328 150272
rect 110380 150260 110386 150272
rect 117130 150260 117136 150272
rect 110380 150232 117136 150260
rect 110380 150220 110386 150232
rect 117130 150220 117136 150232
rect 117188 150220 117194 150272
rect 97902 150152 97908 150204
rect 97960 150192 97966 150204
rect 116854 150192 116860 150204
rect 97960 150164 116860 150192
rect 97960 150152 97966 150164
rect 116854 150152 116860 150164
rect 116912 150152 116918 150204
rect 122834 150152 122840 150204
rect 122892 150192 122898 150204
rect 123708 150192 123714 150204
rect 122892 150164 123714 150192
rect 122892 150152 122898 150164
rect 123708 150152 123714 150164
rect 123766 150152 123772 150204
rect 146386 150152 146392 150204
rect 146444 150192 146450 150204
rect 147536 150192 147542 150204
rect 146444 150164 147542 150192
rect 146444 150152 146450 150164
rect 147536 150152 147542 150164
rect 147594 150152 147600 150204
rect 164326 150152 164332 150204
rect 164384 150192 164390 150204
rect 165476 150192 165482 150204
rect 164384 150164 165482 150192
rect 164384 150152 164390 150164
rect 165476 150152 165482 150164
rect 165534 150152 165540 150204
rect 168374 150152 168380 150204
rect 168432 150192 168438 150204
rect 169340 150192 169346 150204
rect 168432 150164 169346 150192
rect 168432 150152 168438 150164
rect 169340 150152 169346 150164
rect 169398 150152 169404 150204
rect 171134 150152 171140 150204
rect 171192 150192 171198 150204
rect 171916 150192 171922 150204
rect 171192 150164 171922 150192
rect 171192 150152 171198 150164
rect 171916 150152 171922 150164
rect 171974 150152 171980 150204
rect 172698 150152 172704 150204
rect 172756 150192 172762 150204
rect 173848 150192 173854 150204
rect 172756 150164 173854 150192
rect 172756 150152 172762 150164
rect 173848 150152 173854 150164
rect 173906 150152 173912 150204
rect 182266 150152 182272 150204
rect 182324 150192 182330 150204
rect 183416 150192 183422 150204
rect 182324 150164 183422 150192
rect 182324 150152 182330 150164
rect 183416 150152 183422 150164
rect 183474 150152 183480 150204
rect 190822 150152 190828 150204
rect 190880 150192 190886 150204
rect 191788 150192 191794 150204
rect 190880 150164 191794 150192
rect 190880 150152 190886 150164
rect 191788 150152 191794 150164
rect 191846 150152 191852 150204
rect 211246 150152 211252 150204
rect 211304 150192 211310 150204
rect 212304 150192 212310 150204
rect 211304 150164 212310 150192
rect 211304 150152 211310 150164
rect 212304 150152 212310 150164
rect 212362 150152 212368 150204
rect 225046 150152 225052 150204
rect 225104 150192 225110 150204
rect 225828 150192 225834 150204
rect 225104 150164 225834 150192
rect 225104 150152 225110 150164
rect 225828 150152 225834 150164
rect 225886 150152 225892 150204
rect 229186 150152 229192 150204
rect 229244 150192 229250 150204
rect 230336 150192 230342 150204
rect 229244 150164 230342 150192
rect 229244 150152 229250 150164
rect 230336 150152 230342 150164
rect 230394 150152 230400 150204
rect 233234 150152 233240 150204
rect 233292 150192 233298 150204
rect 234200 150192 234206 150204
rect 233292 150164 234206 150192
rect 233292 150152 233298 150164
rect 234200 150152 234206 150164
rect 234258 150152 234264 150204
rect 238938 150152 238944 150204
rect 238996 150192 239002 150204
rect 239996 150192 240002 150204
rect 238996 150164 240002 150192
rect 238996 150152 239002 150164
rect 239996 150152 240002 150164
rect 240054 150152 240060 150204
rect 253934 150152 253940 150204
rect 253992 150192 253998 150204
rect 254716 150192 254722 150204
rect 253992 150164 254722 150192
rect 253992 150152 253998 150164
rect 254716 150152 254722 150164
rect 254774 150152 254780 150204
rect 256786 150152 256792 150204
rect 256844 150192 256850 150204
rect 257936 150192 257942 150204
rect 256844 150164 257942 150192
rect 256844 150152 256850 150164
rect 257936 150152 257942 150164
rect 257994 150152 258000 150204
rect 263594 150152 263600 150204
rect 263652 150192 263658 150204
rect 264376 150192 264382 150204
rect 263652 150164 264382 150192
rect 263652 150152 263658 150164
rect 264376 150152 264382 150164
rect 264434 150152 264440 150204
rect 269114 150152 269120 150204
rect 269172 150192 269178 150204
rect 270172 150192 270178 150204
rect 269172 150164 270178 150192
rect 269172 150152 269178 150164
rect 270172 150152 270178 150164
rect 270230 150152 270236 150204
rect 281534 150152 281540 150204
rect 281592 150192 281598 150204
rect 282316 150192 282322 150204
rect 281592 150164 282322 150192
rect 281592 150152 281598 150164
rect 282316 150152 282322 150164
rect 282374 150152 282380 150204
rect 283098 150152 283104 150204
rect 283156 150192 283162 150204
rect 284248 150192 284254 150204
rect 283156 150164 284254 150192
rect 283156 150152 283162 150164
rect 284248 150152 284254 150164
rect 284306 150152 284312 150204
rect 284386 150152 284392 150204
rect 284444 150192 284450 150204
rect 285536 150192 285542 150204
rect 284444 150164 285542 150192
rect 284444 150152 284450 150164
rect 285536 150152 285542 150164
rect 285594 150152 285600 150204
rect 299474 150152 299480 150204
rect 299532 150192 299538 150204
rect 300348 150192 300354 150204
rect 299532 150164 300354 150192
rect 299532 150152 299538 150164
rect 300348 150152 300354 150164
rect 300406 150152 300412 150204
rect 332686 150152 332692 150204
rect 332744 150192 332750 150204
rect 333744 150192 333750 150204
rect 332744 150164 333750 150192
rect 332744 150152 332750 150164
rect 333744 150152 333750 150164
rect 333802 150152 333808 150204
rect 338298 150152 338304 150204
rect 338356 150192 338362 150204
rect 339448 150192 339454 150204
rect 338356 150164 339454 150192
rect 338356 150152 338362 150164
rect 339448 150152 339454 150164
rect 339506 150152 339512 150204
rect 345106 150152 345112 150204
rect 345164 150192 345170 150204
rect 345888 150192 345894 150204
rect 345164 150164 345894 150192
rect 345164 150152 345170 150164
rect 345888 150152 345894 150164
rect 345946 150152 345952 150204
rect 358906 150152 358912 150204
rect 358964 150192 358970 150204
rect 360056 150192 360062 150204
rect 358964 150164 360062 150192
rect 358964 150152 358970 150164
rect 360056 150152 360062 150164
rect 360114 150152 360120 150204
rect 362954 150152 362960 150204
rect 363012 150192 363018 150204
rect 363920 150192 363926 150204
rect 363012 150164 363926 150192
rect 363012 150152 363018 150164
rect 363920 150152 363926 150164
rect 363978 150152 363984 150204
rect 373994 150152 374000 150204
rect 374052 150192 374058 150204
rect 374776 150192 374782 150204
rect 374052 150164 374782 150192
rect 374052 150152 374058 150164
rect 374776 150152 374782 150164
rect 374834 150152 374840 150204
rect 375558 150152 375564 150204
rect 375616 150192 375622 150204
rect 376708 150192 376714 150204
rect 375616 150164 376714 150192
rect 375616 150152 375622 150164
rect 376708 150152 376714 150164
rect 376766 150152 376772 150204
rect 378134 150152 378140 150204
rect 378192 150192 378198 150204
rect 379284 150192 379290 150204
rect 378192 150164 379290 150192
rect 378192 150152 378198 150164
rect 379284 150152 379290 150164
rect 379342 150152 379348 150204
rect 460934 150152 460940 150204
rect 460992 150192 460998 150204
rect 462084 150192 462090 150204
rect 460992 150164 462090 150192
rect 460992 150152 460998 150164
rect 462084 150152 462090 150164
rect 462142 150152 462148 150204
rect 477678 150152 477684 150204
rect 477736 150192 477742 150204
rect 478828 150192 478834 150204
rect 477736 150164 478834 150192
rect 477736 150152 477742 150164
rect 478828 150152 478834 150164
rect 478886 150152 478892 150204
rect 483198 150152 483204 150204
rect 483256 150192 483262 150204
rect 483980 150192 483986 150204
rect 483256 150164 483986 150192
rect 483256 150152 483262 150164
rect 483980 150152 483986 150164
rect 484038 150152 484044 150204
rect 502334 150152 502340 150204
rect 502392 150192 502398 150204
rect 503208 150192 503214 150204
rect 502392 150164 503214 150192
rect 502392 150152 502398 150164
rect 503208 150152 503214 150164
rect 503266 150152 503272 150204
rect 503714 150152 503720 150204
rect 503772 150192 503778 150204
rect 504496 150192 504502 150204
rect 503772 150164 504502 150192
rect 503772 150152 503778 150164
rect 504496 150152 504502 150164
rect 504554 150152 504560 150204
rect 505278 150152 505284 150204
rect 505336 150192 505342 150204
rect 506428 150192 506434 150204
rect 505336 150164 506434 150192
rect 505336 150152 505342 150164
rect 506428 150152 506434 150164
rect 506486 150152 506492 150204
rect 518020 150152 518026 150204
rect 518078 150192 518084 150204
rect 518802 150192 518808 150204
rect 518078 150164 518808 150192
rect 518078 150152 518084 150164
rect 518802 150152 518808 150164
rect 518860 150152 518866 150204
rect 81342 150084 81348 150136
rect 81400 150124 81406 150136
rect 81400 150096 84194 150124
rect 81400 150084 81406 150096
rect 84166 150056 84194 150096
rect 92474 150084 92480 150136
rect 92532 150124 92538 150136
rect 117222 150124 117228 150136
rect 92532 150096 117228 150124
rect 92532 150084 92538 150096
rect 117222 150084 117228 150096
rect 117280 150084 117286 150136
rect 116486 150056 116492 150068
rect 84166 150028 116492 150056
rect 116486 150016 116492 150028
rect 116544 150016 116550 150068
rect 111150 148384 111156 148436
rect 111208 148424 111214 148436
rect 111208 148396 113174 148424
rect 111208 148384 111214 148396
rect 113146 148356 113174 148396
rect 117038 148356 117044 148368
rect 113146 148328 117044 148356
rect 117038 148316 117044 148328
rect 117096 148316 117102 148368
rect 113082 140700 113088 140752
rect 113140 140740 113146 140752
rect 116118 140740 116124 140752
rect 113140 140712 116124 140740
rect 113140 140700 113146 140712
rect 116118 140700 116124 140712
rect 116176 140700 116182 140752
rect 112990 137912 112996 137964
rect 113048 137952 113054 137964
rect 116118 137952 116124 137964
rect 113048 137924 116124 137952
rect 113048 137912 113054 137924
rect 116118 137912 116124 137924
rect 116176 137912 116182 137964
rect 112806 133832 112812 133884
rect 112864 133872 112870 133884
rect 116026 133872 116032 133884
rect 112864 133844 116032 133872
rect 112864 133832 112870 133844
rect 116026 133832 116032 133844
rect 116084 133832 116090 133884
rect 114186 132608 114192 132660
rect 114244 132648 114250 132660
rect 115198 132648 115204 132660
rect 114244 132620 115204 132648
rect 114244 132608 114250 132620
rect 115198 132608 115204 132620
rect 115256 132608 115262 132660
rect 112898 132404 112904 132456
rect 112956 132444 112962 132456
rect 116118 132444 116124 132456
rect 112956 132416 116124 132444
rect 112956 132404 112962 132416
rect 116118 132404 116124 132416
rect 116176 132404 116182 132456
rect 112714 126896 112720 126948
rect 112772 126936 112778 126948
rect 116118 126936 116124 126948
rect 112772 126908 116124 126936
rect 112772 126896 112778 126908
rect 116118 126896 116124 126908
rect 116176 126896 116182 126948
rect 112622 124108 112628 124160
rect 112680 124148 112686 124160
rect 116118 124148 116124 124160
rect 112680 124120 116124 124148
rect 112680 124108 112686 124120
rect 116118 124108 116124 124120
rect 116176 124108 116182 124160
rect 112530 122748 112536 122800
rect 112588 122788 112594 122800
rect 115934 122788 115940 122800
rect 112588 122760 115940 122788
rect 112588 122748 112594 122760
rect 115934 122748 115940 122760
rect 115992 122748 115998 122800
rect 111702 121388 111708 121440
rect 111760 121428 111766 121440
rect 116118 121428 116124 121440
rect 111760 121400 116124 121428
rect 111760 121388 111766 121400
rect 116118 121388 116124 121400
rect 116176 121388 116182 121440
rect 112438 118600 112444 118652
rect 112496 118640 112502 118652
rect 116118 118640 116124 118652
rect 112496 118612 116124 118640
rect 112496 118600 112502 118612
rect 116118 118600 116124 118612
rect 116176 118600 116182 118652
rect 111610 117240 111616 117292
rect 111668 117280 111674 117292
rect 116118 117280 116124 117292
rect 111668 117252 116124 117280
rect 111668 117240 111674 117252
rect 116118 117240 116124 117252
rect 116176 117240 116182 117292
rect 111518 114452 111524 114504
rect 111576 114492 111582 114504
rect 116118 114492 116124 114504
rect 111576 114464 116124 114492
rect 111576 114452 111582 114464
rect 116118 114452 116124 114464
rect 116176 114452 116182 114504
rect 111426 113092 111432 113144
rect 111484 113132 111490 113144
rect 115934 113132 115940 113144
rect 111484 113104 115940 113132
rect 111484 113092 111490 113104
rect 115934 113092 115940 113104
rect 115992 113092 115998 113144
rect 111334 111732 111340 111784
rect 111392 111772 111398 111784
rect 116118 111772 116124 111784
rect 111392 111744 116124 111772
rect 111392 111732 111398 111744
rect 116118 111732 116124 111744
rect 116176 111732 116182 111784
rect 111150 108944 111156 108996
rect 111208 108984 111214 108996
rect 116118 108984 116124 108996
rect 111208 108956 116124 108984
rect 111208 108944 111214 108956
rect 116118 108944 116124 108956
rect 116176 108944 116182 108996
rect 111242 92420 111248 92472
rect 111300 92460 111306 92472
rect 116118 92460 116124 92472
rect 111300 92432 116124 92460
rect 111300 92420 111306 92432
rect 116118 92420 116124 92432
rect 116176 92420 116182 92472
rect 111058 89632 111064 89684
rect 111116 89672 111122 89684
rect 116118 89672 116124 89684
rect 111116 89644 116124 89672
rect 111116 89632 111122 89644
rect 116118 89632 116124 89644
rect 116176 89632 116182 89684
rect 113818 88272 113824 88324
rect 113876 88312 113882 88324
rect 116026 88312 116032 88324
rect 113876 88284 116032 88312
rect 113876 88272 113882 88284
rect 116026 88272 116032 88284
rect 116084 88272 116090 88324
rect 113910 83920 113916 83972
rect 113968 83960 113974 83972
rect 116578 83960 116584 83972
rect 113968 83932 116584 83960
rect 113968 83920 113974 83932
rect 116578 83920 116584 83932
rect 116636 83920 116642 83972
rect 114002 82764 114008 82816
rect 114060 82804 114066 82816
rect 116210 82804 116216 82816
rect 114060 82776 116216 82804
rect 114060 82764 114066 82776
rect 116210 82764 116216 82776
rect 116268 82764 116274 82816
rect 114094 79976 114100 80028
rect 114152 80016 114158 80028
rect 115934 80016 115940 80028
rect 114152 79988 115940 80016
rect 114152 79976 114158 79988
rect 115934 79976 115940 79988
rect 115992 79976 115998 80028
rect 114186 78616 114192 78668
rect 114244 78656 114250 78668
rect 116118 78656 116124 78668
rect 114244 78628 116124 78656
rect 114244 78616 114250 78628
rect 116118 78616 116124 78628
rect 116176 78616 116182 78668
rect 114186 71748 114192 71800
rect 114244 71788 114250 71800
rect 116578 71788 116584 71800
rect 114244 71760 116584 71788
rect 114244 71748 114250 71760
rect 116578 71748 116584 71760
rect 116636 71748 116642 71800
rect 114094 69028 114100 69080
rect 114152 69068 114158 69080
rect 116302 69068 116308 69080
rect 114152 69040 116308 69068
rect 114152 69028 114158 69040
rect 116302 69028 116308 69040
rect 116360 69028 116366 69080
rect 114002 67600 114008 67652
rect 114060 67640 114066 67652
rect 116118 67640 116124 67652
rect 114060 67612 116124 67640
rect 114060 67600 114066 67612
rect 116118 67600 116124 67612
rect 116176 67600 116182 67652
rect 113910 66240 113916 66292
rect 113968 66280 113974 66292
rect 116578 66280 116584 66292
rect 113968 66252 116584 66280
rect 113968 66240 113974 66252
rect 116578 66240 116584 66252
rect 116636 66240 116642 66292
rect 113358 64676 113364 64728
rect 113416 64716 113422 64728
rect 116578 64716 116584 64728
rect 113416 64688 116584 64716
rect 113416 64676 113422 64688
rect 116578 64676 116584 64688
rect 116636 64676 116642 64728
rect 113818 63520 113824 63572
rect 113876 63560 113882 63572
rect 116210 63560 116216 63572
rect 113876 63532 116216 63560
rect 113876 63520 113882 63532
rect 116210 63520 116216 63532
rect 116268 63520 116274 63572
rect 112438 62092 112444 62144
rect 112496 62132 112502 62144
rect 116118 62132 116124 62144
rect 112496 62104 116124 62132
rect 112496 62092 112502 62104
rect 116118 62092 116124 62104
rect 116176 62092 116182 62144
rect 112530 42780 112536 42832
rect 112588 42820 112594 42832
rect 116118 42820 116124 42832
rect 112588 42792 116124 42820
rect 112588 42780 112594 42792
rect 116118 42780 116124 42792
rect 116176 42780 116182 42832
rect 116670 7896 116676 7948
rect 116728 7896 116734 7948
rect 116854 7896 116860 7948
rect 116912 7896 116918 7948
rect 116688 7596 116716 7896
rect 116872 7744 116900 7896
rect 117038 7760 117044 7812
rect 117096 7800 117102 7812
rect 117314 7800 117320 7812
rect 117096 7772 117320 7800
rect 117096 7760 117102 7772
rect 117314 7760 117320 7772
rect 117372 7760 117378 7812
rect 116854 7692 116860 7744
rect 116912 7692 116918 7744
rect 116762 7624 116768 7676
rect 116820 7664 116826 7676
rect 117222 7664 117228 7676
rect 116820 7636 117228 7664
rect 116820 7624 116826 7636
rect 117222 7624 117228 7636
rect 117280 7624 117286 7676
rect 116688 7568 116992 7596
rect 116964 7460 116992 7568
rect 117038 7460 117044 7472
rect 116964 7432 117044 7460
rect 117038 7420 117044 7432
rect 117096 7420 117102 7472
rect 111702 2796 111708 2848
rect 111760 2836 111766 2848
rect 111760 2808 193628 2836
rect 111760 2796 111766 2808
rect 193600 2508 193628 2808
rect 425808 2808 443684 2836
rect 425808 2508 425836 2808
rect 443656 2508 443684 2808
rect 193582 2456 193588 2508
rect 193640 2456 193646 2508
rect 425790 2456 425796 2508
rect 425848 2456 425854 2508
rect 443638 2456 443644 2508
rect 443696 2456 443702 2508
rect 111058 1952 111064 1964
rect 92446 1924 104480 1952
rect 62390 1844 62396 1896
rect 62448 1884 62454 1896
rect 65334 1884 65340 1896
rect 62448 1856 65340 1884
rect 62448 1844 62454 1856
rect 65334 1844 65340 1856
rect 65392 1844 65398 1896
rect 68002 1844 68008 1896
rect 68060 1884 68066 1896
rect 89254 1884 89260 1896
rect 68060 1856 89260 1884
rect 68060 1844 68066 1856
rect 89254 1844 89260 1856
rect 89312 1844 89318 1896
rect 89346 1844 89352 1896
rect 89404 1884 89410 1896
rect 92446 1884 92474 1924
rect 89404 1856 92474 1884
rect 89404 1844 89410 1856
rect 97166 1844 97172 1896
rect 97224 1884 97230 1896
rect 104342 1884 104348 1896
rect 97224 1856 104348 1884
rect 97224 1844 97230 1856
rect 104342 1844 104348 1856
rect 104400 1844 104406 1896
rect 64138 1776 64144 1828
rect 64196 1816 64202 1828
rect 69382 1816 69388 1828
rect 64196 1788 69388 1816
rect 64196 1776 64202 1788
rect 69382 1776 69388 1788
rect 69440 1776 69446 1828
rect 75638 1776 75644 1828
rect 75696 1816 75702 1828
rect 85390 1816 85396 1828
rect 75696 1788 85396 1816
rect 75696 1776 75702 1788
rect 85390 1776 85396 1788
rect 85448 1776 85454 1828
rect 86034 1776 86040 1828
rect 86092 1816 86098 1828
rect 104452 1816 104480 1924
rect 105832 1924 111064 1952
rect 105832 1896 105860 1924
rect 111058 1912 111064 1924
rect 111116 1912 111122 1964
rect 104526 1844 104532 1896
rect 104584 1884 104590 1896
rect 105722 1884 105728 1896
rect 104584 1856 105728 1884
rect 104584 1844 104590 1856
rect 105722 1844 105728 1856
rect 105780 1844 105786 1896
rect 105814 1844 105820 1896
rect 105872 1844 105878 1896
rect 105906 1844 105912 1896
rect 105964 1884 105970 1896
rect 109218 1884 109224 1896
rect 105964 1856 109224 1884
rect 105964 1844 105970 1856
rect 109218 1844 109224 1856
rect 109276 1844 109282 1896
rect 109310 1844 109316 1896
rect 109368 1884 109374 1896
rect 109368 1856 110184 1884
rect 109368 1844 109374 1856
rect 109586 1816 109592 1828
rect 86092 1788 104204 1816
rect 104452 1788 109592 1816
rect 86092 1776 86098 1788
rect 62666 1708 62672 1760
rect 62724 1748 62730 1760
rect 77202 1748 77208 1760
rect 62724 1720 77208 1748
rect 62724 1708 62730 1720
rect 77202 1708 77208 1720
rect 77260 1708 77266 1760
rect 82630 1708 82636 1760
rect 82688 1748 82694 1760
rect 104066 1748 104072 1760
rect 82688 1720 104072 1748
rect 82688 1708 82694 1720
rect 104066 1708 104072 1720
rect 104124 1708 104130 1760
rect 104176 1748 104204 1788
rect 109586 1776 109592 1788
rect 109644 1776 109650 1828
rect 109954 1748 109960 1760
rect 104176 1720 109960 1748
rect 109954 1708 109960 1720
rect 110012 1708 110018 1760
rect 110156 1748 110184 1856
rect 112438 1748 112444 1760
rect 110156 1720 112444 1748
rect 112438 1708 112444 1720
rect 112496 1708 112502 1760
rect 69290 1640 69296 1692
rect 69348 1680 69354 1692
rect 102594 1680 102600 1692
rect 69348 1652 102600 1680
rect 69348 1640 69354 1652
rect 102594 1640 102600 1652
rect 102652 1640 102658 1692
rect 102686 1640 102692 1692
rect 102744 1680 102750 1692
rect 105814 1680 105820 1692
rect 102744 1652 105820 1680
rect 102744 1640 102750 1652
rect 105814 1640 105820 1652
rect 105872 1640 105878 1692
rect 106182 1640 106188 1692
rect 106240 1680 106246 1692
rect 116578 1680 116584 1692
rect 106240 1652 116584 1680
rect 106240 1640 106246 1652
rect 116578 1640 116584 1652
rect 116636 1640 116642 1692
rect 59354 1572 59360 1624
rect 59412 1612 59418 1624
rect 68462 1612 68468 1624
rect 59412 1584 68468 1612
rect 59412 1572 59418 1584
rect 68462 1572 68468 1584
rect 68520 1572 68526 1624
rect 79318 1572 79324 1624
rect 79376 1612 79382 1624
rect 97258 1612 97264 1624
rect 79376 1584 97264 1612
rect 79376 1572 79382 1584
rect 97258 1572 97264 1584
rect 97316 1572 97322 1624
rect 99374 1572 99380 1624
rect 99432 1612 99438 1624
rect 105906 1612 105912 1624
rect 99432 1584 105912 1612
rect 99432 1572 99438 1584
rect 105906 1572 105912 1584
rect 105964 1572 105970 1624
rect 105998 1572 106004 1624
rect 106056 1612 106062 1624
rect 110046 1612 110052 1624
rect 106056 1584 110052 1612
rect 106056 1572 106062 1584
rect 110046 1572 110052 1584
rect 110104 1572 110110 1624
rect 72694 1504 72700 1556
rect 72752 1544 72758 1556
rect 110506 1544 110512 1556
rect 72752 1516 110512 1544
rect 72752 1504 72758 1516
rect 110506 1504 110512 1516
rect 110564 1504 110570 1556
rect 42610 1436 42616 1488
rect 42668 1476 42674 1488
rect 68278 1476 68284 1488
rect 42668 1448 68284 1476
rect 42668 1436 42674 1448
rect 68278 1436 68284 1448
rect 68336 1436 68342 1488
rect 87966 1436 87972 1488
rect 88024 1476 88030 1488
rect 97166 1476 97172 1488
rect 88024 1448 97172 1476
rect 88024 1436 88030 1448
rect 97166 1436 97172 1448
rect 97224 1436 97230 1488
rect 97258 1436 97264 1488
rect 97316 1476 97322 1488
rect 108206 1476 108212 1488
rect 97316 1448 108212 1476
rect 97316 1436 97322 1448
rect 108206 1436 108212 1448
rect 108264 1436 108270 1488
rect 108298 1436 108304 1488
rect 108356 1476 108362 1488
rect 143626 1476 143632 1488
rect 108356 1448 143632 1476
rect 108356 1436 108362 1448
rect 143626 1436 143632 1448
rect 143684 1436 143690 1488
rect 46014 1368 46020 1420
rect 46072 1408 46078 1420
rect 116486 1408 116492 1420
rect 46072 1380 116492 1408
rect 46072 1368 46078 1380
rect 116486 1368 116492 1380
rect 116544 1368 116550 1420
rect 294782 1408 294788 1420
rect 293926 1380 294788 1408
rect 55950 1300 55956 1352
rect 56008 1340 56014 1352
rect 293926 1340 293954 1380
rect 294782 1368 294788 1380
rect 294840 1408 294846 1420
rect 343634 1408 343640 1420
rect 294840 1380 343640 1408
rect 294840 1368 294846 1380
rect 343634 1368 343640 1380
rect 343692 1368 343698 1420
rect 491294 1368 491300 1420
rect 491352 1408 491358 1420
rect 493594 1408 493600 1420
rect 491352 1380 493600 1408
rect 491352 1368 491358 1380
rect 493594 1368 493600 1380
rect 493652 1368 493658 1420
rect 56008 1312 293954 1340
rect 56008 1300 56014 1312
rect 2682 1232 2688 1284
rect 2740 1272 2746 1284
rect 116302 1272 116308 1284
rect 2740 1244 116308 1272
rect 2740 1232 2746 1244
rect 116302 1232 116308 1244
rect 116360 1232 116366 1284
rect 39298 1164 39304 1216
rect 39356 1204 39362 1216
rect 116394 1204 116400 1216
rect 39356 1176 116400 1204
rect 39356 1164 39362 1176
rect 116394 1164 116400 1176
rect 116452 1164 116458 1216
rect 49326 1096 49332 1148
rect 49384 1136 49390 1148
rect 116762 1136 116768 1148
rect 49384 1108 116768 1136
rect 49384 1096 49390 1108
rect 116762 1096 116768 1108
rect 116820 1096 116826 1148
rect 52638 1028 52644 1080
rect 52696 1068 52702 1080
rect 117222 1068 117228 1080
rect 52696 1040 117228 1068
rect 52696 1028 52702 1040
rect 117222 1028 117228 1040
rect 117280 1028 117286 1080
rect 65978 960 65984 1012
rect 66036 1000 66042 1012
rect 116854 1000 116860 1012
rect 66036 972 116860 1000
rect 66036 960 66042 972
rect 116854 960 116860 972
rect 116912 960 116918 1012
rect 76006 892 76012 944
rect 76064 932 76070 944
rect 112530 932 112536 944
rect 76064 904 112536 932
rect 76064 892 76070 904
rect 112530 892 112536 904
rect 112588 892 112594 944
rect 91738 824 91744 876
rect 91796 864 91802 876
rect 99742 864 99748 876
rect 91796 836 99748 864
rect 91796 824 91802 836
rect 99742 824 99748 836
rect 99800 824 99806 876
rect 103882 824 103888 876
rect 103940 864 103946 876
rect 108298 864 108304 876
rect 103940 836 108304 864
rect 103940 824 103946 836
rect 108298 824 108304 836
rect 108356 824 108362 876
rect 95694 756 95700 808
rect 95752 796 95758 808
rect 99558 796 99564 808
rect 95752 768 99564 796
rect 95752 756 95758 768
rect 99558 756 99564 768
rect 99616 756 99622 808
<< via1 >>
rect 129924 160760 129976 160812
rect 134156 160760 134208 160812
rect 63408 160012 63460 160064
rect 143264 160012 143316 160064
rect 143356 160012 143408 160064
rect 156604 160012 156656 160064
rect 156788 160012 156840 160064
rect 191748 160012 191800 160064
rect 197176 160012 197228 160064
rect 207020 160012 207072 160064
rect 211436 160012 211488 160064
rect 280344 160012 280396 160064
rect 281264 160012 281316 160064
rect 332692 160012 332744 160064
rect 334256 160012 334308 160064
rect 374092 160012 374144 160064
rect 378876 160012 378928 160064
rect 398564 160012 398616 160064
rect 25596 159944 25648 159996
rect 109776 159944 109828 159996
rect 117228 159944 117280 159996
rect 191472 159944 191524 159996
rect 198004 159944 198056 159996
rect 269120 159944 269172 159996
rect 271236 159944 271288 159996
rect 271880 159944 271932 159996
rect 275376 159944 275428 159996
rect 329104 159944 329156 159996
rect 329196 159944 329248 159996
rect 369952 159944 370004 159996
rect 374644 159944 374696 159996
rect 388168 159944 388220 159996
rect 389824 159944 389876 159996
rect 413836 159944 413888 159996
rect 76932 159876 76984 159928
rect 162492 159876 162544 159928
rect 166908 159876 166960 159928
rect 186688 159876 186740 159928
rect 191288 159876 191340 159928
rect 264888 159876 264940 159928
rect 268660 159876 268712 159928
rect 324044 159876 324096 159928
rect 328368 159876 328420 159928
rect 369492 159876 369544 159928
rect 372160 159876 372212 159928
rect 396172 159876 396224 159928
rect 403256 159876 403308 159928
rect 416596 159876 416648 159928
rect 476120 159876 476172 159928
rect 480628 159876 480680 159928
rect 485964 159876 486016 159928
rect 56692 159808 56744 159860
rect 132960 159808 133012 159860
rect 133144 159808 133196 159860
rect 143172 159808 143224 159860
rect 143264 159808 143316 159860
rect 146576 159808 146628 159860
rect 146668 159808 146720 159860
rect 176660 159808 176712 159860
rect 184572 159808 184624 159860
rect 259552 159808 259604 159860
rect 261944 159808 261996 159860
rect 318892 159808 318944 159860
rect 320824 159808 320876 159860
rect 362960 159808 363012 159860
rect 376300 159808 376352 159860
rect 406200 159808 406252 159860
rect 409972 159808 410024 159860
rect 417884 159808 417936 159860
rect 424324 159808 424376 159860
rect 442816 159808 442868 159860
rect 446128 159808 446180 159860
rect 456800 159808 456852 159860
rect 458732 159808 458784 159860
rect 465080 159808 465132 159860
rect 470508 159808 470560 159860
rect 471428 159808 471480 159860
rect 477684 159808 477736 159860
rect 70124 159740 70176 159792
rect 156328 159740 156380 159792
rect 156604 159740 156656 159792
rect 160100 159740 160152 159792
rect 177856 159740 177908 159792
rect 253940 159740 253992 159792
rect 255228 159740 255280 159792
rect 313464 159740 313516 159792
rect 314108 159740 314160 159792
rect 357992 159740 358044 159792
rect 365444 159740 365496 159792
rect 395528 159740 395580 159792
rect 396540 159740 396592 159792
rect 413928 159740 413980 159792
rect 420920 159740 420972 159792
rect 440424 159740 440476 159792
rect 450360 159740 450412 159792
rect 462320 159740 462372 159792
rect 473084 159740 473136 159792
rect 480076 159740 480128 159792
rect 18880 159672 18932 159724
rect 109132 159672 109184 159724
rect 113088 159672 113140 159724
rect 126428 159672 126480 159724
rect 126520 159672 126572 159724
rect 156512 159672 156564 159724
rect 49976 159604 50028 159656
rect 132868 159604 132920 159656
rect 43260 159536 43312 159588
rect 136548 159604 136600 159656
rect 136640 159604 136692 159656
rect 139400 159604 139452 159656
rect 139952 159604 140004 159656
rect 163780 159672 163832 159724
rect 167736 159672 167788 159724
rect 246948 159672 247000 159724
rect 248512 159672 248564 159724
rect 161020 159604 161072 159656
rect 240324 159604 240376 159656
rect 244280 159604 244332 159656
rect 305368 159604 305420 159656
rect 308220 159672 308272 159724
rect 342628 159672 342680 159724
rect 342720 159672 342772 159724
rect 343824 159672 343876 159724
rect 347780 159672 347832 159724
rect 378784 159672 378836 159724
rect 379704 159672 379756 159724
rect 405832 159672 405884 159724
rect 417516 159672 417568 159724
rect 437664 159672 437716 159724
rect 449532 159672 449584 159724
rect 460940 159672 460992 159724
rect 463792 159672 463844 159724
rect 471428 159672 471480 159724
rect 478972 159672 479024 159724
rect 484676 159672 484728 159724
rect 308588 159604 308640 159656
rect 309048 159604 309100 159656
rect 341616 159604 341668 159656
rect 134156 159536 134208 159588
rect 154488 159536 154540 159588
rect 157616 159536 157668 159588
rect 239312 159536 239364 159588
rect 250996 159536 251048 159588
rect 310612 159536 310664 159588
rect 315764 159536 315816 159588
rect 342812 159604 342864 159656
rect 354220 159604 354272 159656
rect 357808 159604 357860 159656
rect 369216 159604 369268 159656
rect 369584 159604 369636 159656
rect 401048 159604 401100 159656
rect 407488 159604 407540 159656
rect 429936 159604 429988 159656
rect 453764 159604 453816 159656
rect 465264 159604 465316 159656
rect 468024 159604 468076 159656
rect 476028 159604 476080 159656
rect 479800 159604 479852 159656
rect 485228 159604 485280 159656
rect 358912 159536 358964 159588
rect 362868 159536 362920 159588
rect 394976 159536 395028 159588
rect 399024 159536 399076 159588
rect 408500 159536 408552 159588
rect 410800 159536 410852 159588
rect 432512 159536 432564 159588
rect 452016 159536 452068 159588
rect 463976 159536 464028 159588
rect 467196 159536 467248 159588
rect 473360 159536 473412 159588
rect 32312 159468 32364 159520
rect 36544 159400 36596 159452
rect 126244 159400 126296 159452
rect 126428 159468 126480 159520
rect 127624 159468 127676 159520
rect 133236 159468 133288 159520
rect 144092 159468 144144 159520
rect 144184 159468 144236 159520
rect 225328 159468 225380 159520
rect 230848 159468 230900 159520
rect 293960 159468 294012 159520
rect 294788 159468 294840 159520
rect 126796 159400 126848 159452
rect 6276 159332 6328 159384
rect 122840 159332 122892 159384
rect 123116 159332 123168 159384
rect 147772 159400 147824 159452
rect 150900 159400 150952 159452
rect 233240 159400 233292 159452
rect 234988 159400 235040 159452
rect 298008 159400 298060 159452
rect 301504 159400 301556 159452
rect 341432 159400 341484 159452
rect 341616 159468 341668 159520
rect 354864 159468 354916 159520
rect 356152 159468 356204 159520
rect 390560 159468 390612 159520
rect 400772 159468 400824 159520
rect 424876 159468 424928 159520
rect 459652 159468 459704 159520
rect 466644 159468 466696 159520
rect 468852 159468 468904 159520
rect 474832 159468 474884 159520
rect 477316 159468 477368 159520
rect 483296 159468 483348 159520
rect 342260 159400 342312 159452
rect 342352 159400 342404 159452
rect 349344 159400 349396 159452
rect 358636 159400 358688 159452
rect 392768 159400 392820 159452
rect 404084 159400 404136 159452
rect 427360 159400 427412 159452
rect 427636 159400 427688 159452
rect 445392 159400 445444 159452
rect 451188 159400 451240 159452
rect 462872 159400 462924 159452
rect 518808 159400 518860 159452
rect 522672 159400 522724 159452
rect 132684 159332 132736 159384
rect 137100 159332 137152 159384
rect 137468 159332 137520 159384
rect 223580 159332 223632 159384
rect 231676 159332 231728 159384
rect 295524 159332 295576 159384
rect 295616 159332 295668 159384
rect 342444 159332 342496 159384
rect 346032 159332 346084 159384
rect 382832 159332 382884 159384
rect 383108 159332 383160 159384
rect 411352 159332 411404 159384
rect 414204 159332 414256 159384
rect 435088 159332 435140 159384
rect 448704 159332 448756 159384
rect 461400 159332 461452 159384
rect 469680 159332 469732 159384
rect 477408 159332 477460 159384
rect 478144 159332 478196 159384
rect 483204 159332 483256 159384
rect 518716 159332 518768 159384
rect 523500 159332 523552 159384
rect 73528 159264 73580 159316
rect 80060 159264 80112 159316
rect 83648 159264 83700 159316
rect 167000 159264 167052 159316
rect 170220 159264 170272 159316
rect 195152 159264 195204 159316
rect 195244 159264 195296 159316
rect 201316 159264 201368 159316
rect 201408 159264 201460 159316
rect 212632 159264 212684 159316
rect 214012 159264 214064 159316
rect 281540 159264 281592 159316
rect 282092 159264 282144 159316
rect 334348 159264 334400 159316
rect 335084 159264 335136 159316
rect 374000 159264 374052 159316
rect 374644 159264 374696 159316
rect 382280 159264 382332 159316
rect 388996 159264 389048 159316
rect 404268 159264 404320 159316
rect 457904 159264 457956 159316
rect 464436 159264 464488 159316
rect 80244 159196 80296 159248
rect 91100 159196 91152 159248
rect 100484 159196 100536 159248
rect 184388 159196 184440 159248
rect 187056 159196 187108 159248
rect 214656 159196 214708 159248
rect 218244 159196 218296 159248
rect 284392 159196 284444 159248
rect 287980 159196 288032 159248
rect 338764 159196 338816 159248
rect 339316 159196 339368 159248
rect 377956 159196 378008 159248
rect 86960 159128 87012 159180
rect 93676 159060 93728 159112
rect 162860 159060 162912 159112
rect 163044 159128 163096 159180
rect 172152 159128 172204 159180
rect 173624 159128 173676 159180
rect 193680 159128 193732 159180
rect 193772 159128 193824 159180
rect 218060 159128 218112 159180
rect 224960 159128 225012 159180
rect 290648 159128 290700 159180
rect 293960 159128 294012 159180
rect 295156 159128 295208 159180
rect 302332 159128 302384 159180
rect 169760 159060 169812 159112
rect 171140 159060 171192 159112
rect 173164 159060 173216 159112
rect 180340 159060 180392 159112
rect 204904 159060 204956 159112
rect 220728 159060 220780 159112
rect 283196 159060 283248 159112
rect 284668 159060 284720 159112
rect 285772 159060 285824 159112
rect 107200 158992 107252 159044
rect 183468 158992 183520 159044
rect 183744 158992 183796 159044
rect 195244 158992 195296 159044
rect 203892 158992 203944 159044
rect 213828 158992 213880 159044
rect 214840 158992 214892 159044
rect 222108 158992 222160 159044
rect 224132 158992 224184 159044
rect 288072 159060 288124 159112
rect 288900 159060 288952 159112
rect 338304 159060 338356 159112
rect 338488 159060 338540 159112
rect 339684 159060 339736 159112
rect 341432 159128 341484 159180
rect 345664 159128 345716 159180
rect 345756 159128 345808 159180
rect 351828 159128 351880 159180
rect 351920 159128 351972 159180
rect 385500 159196 385552 159248
rect 385592 159196 385644 159248
rect 398840 159196 398892 159248
rect 457076 159196 457128 159248
rect 464160 159196 464212 159248
rect 349252 159060 349304 159112
rect 349344 159060 349396 159112
rect 298100 158992 298152 159044
rect 300400 158992 300452 159044
rect 307392 158992 307444 159044
rect 345572 158992 345624 159044
rect 345848 158992 345900 159044
rect 349068 158992 349120 159044
rect 351092 158992 351144 159044
rect 374644 158992 374696 159044
rect 378048 159060 378100 159112
rect 388444 159128 388496 159180
rect 392308 159128 392360 159180
rect 404176 159128 404228 159180
rect 461308 159128 461360 159180
rect 468024 159128 468076 159180
rect 395712 159060 395764 159112
rect 405372 159060 405424 159112
rect 405740 159060 405792 159112
rect 409236 159060 409288 159112
rect 460480 159060 460532 159112
rect 466460 159060 466512 159112
rect 472256 159060 472308 159112
rect 479156 159060 479208 159112
rect 378232 158992 378284 159044
rect 447876 158992 447928 159044
rect 460112 158992 460164 159044
rect 462136 158992 462188 159044
rect 467932 158992 467984 159044
rect 473912 158992 473964 159044
rect 480260 158992 480312 159044
rect 96252 158924 96304 158976
rect 121920 158924 121972 158976
rect 124036 158924 124088 158976
rect 193588 158924 193640 158976
rect 193680 158924 193732 158976
rect 197360 158924 197412 158976
rect 200580 158924 200632 158976
rect 224960 158924 225012 158976
rect 237564 158924 237616 158976
rect 299480 158924 299532 158976
rect 314936 158924 314988 158976
rect 357532 158924 357584 158976
rect 361212 158924 361264 158976
rect 102968 158856 103020 158908
rect 125508 158856 125560 158908
rect 126244 158856 126296 158908
rect 129740 158856 129792 158908
rect 130752 158856 130804 158908
rect 195060 158856 195112 158908
rect 195152 158856 195204 158908
rect 198924 158856 198976 158908
rect 208124 158856 208176 158908
rect 212448 158856 212500 158908
rect 109684 158788 109736 158840
rect 132684 158788 132736 158840
rect 133420 158788 133472 158840
rect 158720 158788 158772 158840
rect 163504 158788 163556 158840
rect 195980 158788 196032 158840
rect 207296 158788 207348 158840
rect 230756 158856 230808 158908
rect 241796 158856 241848 158908
rect 303528 158856 303580 158908
rect 305644 158856 305696 158908
rect 307668 158856 307720 158908
rect 310704 158856 310756 158908
rect 312176 158856 312228 158908
rect 312452 158856 312504 158908
rect 313372 158856 313424 158908
rect 322480 158856 322532 158908
rect 365168 158856 365220 158908
rect 217324 158788 217376 158840
rect 220360 158788 220412 158840
rect 238392 158788 238444 158840
rect 242440 158788 242492 158840
rect 261116 158788 261168 158840
rect 317052 158788 317104 158840
rect 319168 158788 319220 158840
rect 321560 158788 321612 158840
rect 327540 158788 327592 158840
rect 330484 158788 330536 158840
rect 90364 158720 90416 158772
rect 92572 158720 92624 158772
rect 92848 158720 92900 158772
rect 114468 158720 114520 158772
rect 119804 158720 119856 158772
rect 147128 158720 147180 158772
rect 147588 158720 147640 158772
rect 149520 158720 149572 158772
rect 153476 158720 153528 158772
rect 179420 158720 179472 158772
rect 194692 158720 194744 158772
rect 203708 158720 203760 158772
rect 210608 158720 210660 158772
rect 215392 158720 215444 158772
rect 221556 158720 221608 158772
rect 224408 158720 224460 158772
rect 240876 158720 240928 158772
rect 243360 158720 243412 158772
rect 254400 158720 254452 158772
rect 255412 158720 255464 158772
rect 258540 158720 258592 158772
rect 260932 158720 260984 158772
rect 264428 158720 264480 158772
rect 266360 158720 266412 158772
rect 267832 158720 267884 158772
rect 320272 158720 320324 158772
rect 321652 158720 321704 158772
rect 81072 158652 81124 158704
rect 180892 158652 180944 158704
rect 181996 158652 182048 158704
rect 256792 158652 256844 158704
rect 363144 158788 363196 158840
rect 369216 158924 369268 158976
rect 384948 158924 385000 158976
rect 416688 158924 416740 158976
rect 419540 158924 419592 158976
rect 456248 158924 456300 158976
rect 463148 158924 463200 158976
rect 466368 158924 466420 158976
rect 472624 158924 472676 158976
rect 475568 158924 475620 158976
rect 481640 158924 481692 158976
rect 374552 158788 374604 158840
rect 374736 158788 374788 158840
rect 386144 158856 386196 158908
rect 391480 158856 391532 158908
rect 394332 158856 394384 158908
rect 412548 158856 412600 158908
rect 412916 158856 412968 158908
rect 420092 158856 420144 158908
rect 423220 158856 423272 158908
rect 454592 158856 454644 158908
rect 461860 158856 461912 158908
rect 465540 158856 465592 158908
rect 472256 158856 472308 158908
rect 474740 158856 474792 158908
rect 481364 158856 481416 158908
rect 482284 158856 482336 158908
rect 487252 158856 487304 158908
rect 508320 158856 508372 158908
rect 510068 158856 510120 158908
rect 384764 158788 384816 158840
rect 389180 158788 389232 158840
rect 455420 158788 455472 158840
rect 462780 158788 462832 158840
rect 464620 158788 464672 158840
rect 471520 158788 471572 158840
rect 476396 158788 476448 158840
rect 482652 158788 482704 158840
rect 505284 158788 505336 158840
rect 507584 158788 507636 158840
rect 330668 158720 330720 158772
rect 367192 158720 367244 158772
rect 367928 158720 367980 158772
rect 386236 158720 386288 158772
rect 388076 158720 388128 158772
rect 390376 158720 390428 158772
rect 409144 158720 409196 158772
rect 410524 158720 410576 158772
rect 413376 158720 413428 158772
rect 419632 158720 419684 158772
rect 452844 158720 452896 158772
rect 459560 158720 459612 158772
rect 462964 158720 463016 158772
rect 469220 158720 469272 158772
rect 481456 158720 481508 158772
rect 486516 158720 486568 158772
rect 505744 158720 505796 158772
rect 506756 158720 506808 158772
rect 507032 158720 507084 158772
rect 508412 158720 508464 158772
rect 509424 158720 509476 158772
rect 511724 158720 511776 158772
rect 514944 158720 514996 158772
rect 518532 158720 518584 158772
rect 67640 158584 67692 158636
rect 170312 158584 170364 158636
rect 171968 158584 172020 158636
rect 250076 158584 250128 158636
rect 74356 158516 74408 158568
rect 71044 158448 71096 158500
rect 173072 158448 173124 158500
rect 175280 158516 175332 158568
rect 252744 158516 252796 158568
rect 175372 158448 175424 158500
rect 178684 158448 178736 158500
rect 255596 158448 255648 158500
rect 60924 158380 60976 158432
rect 164332 158380 164384 158432
rect 165252 158380 165304 158432
rect 245016 158380 245068 158432
rect 64236 158312 64288 158364
rect 167552 158312 167604 158364
rect 168564 158312 168616 158364
rect 247132 158312 247184 158364
rect 54208 158244 54260 158296
rect 160284 158244 160336 158296
rect 161848 158244 161900 158296
rect 242072 158244 242124 158296
rect 47492 158176 47544 158228
rect 155040 158176 155092 158228
rect 155132 158176 155184 158228
rect 237380 158176 237432 158228
rect 256884 158176 256936 158228
rect 315028 158176 315080 158228
rect 50804 158108 50856 158160
rect 157708 158108 157760 158160
rect 158444 158108 158496 158160
rect 238944 158108 238996 158160
rect 246764 158108 246816 158160
rect 306932 158108 306984 158160
rect 37372 158040 37424 158092
rect 146392 158040 146444 158092
rect 148416 158040 148468 158092
rect 231952 158040 232004 158092
rect 243452 158040 243504 158092
rect 304724 158040 304776 158092
rect 388 157972 440 158024
rect 118884 157972 118936 158024
rect 131580 157972 131632 158024
rect 219348 157972 219400 158024
rect 236736 157972 236788 158024
rect 299664 157972 299716 158024
rect 77760 157904 77812 157956
rect 84476 157836 84528 157888
rect 175924 157836 175976 157888
rect 176200 157904 176252 157956
rect 182272 157904 182324 157956
rect 185400 157904 185452 157956
rect 260472 157904 260524 157956
rect 178040 157836 178092 157888
rect 179420 157836 179472 157888
rect 87788 157768 87840 157820
rect 184756 157768 184808 157820
rect 184940 157836 184992 157888
rect 185952 157836 186004 157888
rect 188804 157836 188856 157888
rect 263048 157836 263100 157888
rect 185216 157768 185268 157820
rect 91192 157700 91244 157752
rect 185308 157700 185360 157752
rect 94596 157632 94648 157684
rect 190644 157768 190696 157820
rect 195520 157768 195572 157820
rect 267740 157768 267792 157820
rect 185676 157700 185728 157752
rect 188528 157700 188580 157752
rect 190460 157700 190512 157752
rect 263692 157700 263744 157752
rect 185584 157632 185636 157684
rect 236092 157632 236144 157684
rect 97908 157564 97960 157616
rect 193312 157564 193364 157616
rect 197360 157564 197412 157616
rect 251456 157564 251508 157616
rect 111340 157496 111392 157548
rect 203432 157496 203484 157548
rect 204904 157496 204956 157548
rect 255872 157496 255924 157548
rect 114744 157428 114796 157480
rect 206560 157428 206612 157480
rect 141700 157360 141752 157412
rect 227076 157360 227128 157412
rect 49148 157292 49200 157344
rect 156420 157292 156472 157344
rect 158720 157292 158772 157344
rect 214472 157292 214524 157344
rect 214564 157292 214616 157344
rect 221372 157292 221424 157344
rect 224224 157292 224276 157344
rect 281632 157292 281684 157344
rect 45744 157224 45796 157276
rect 153844 157224 153896 157276
rect 163780 157224 163832 157276
rect 166448 157224 166500 157276
rect 192116 157224 192168 157276
rect 265164 157224 265216 157276
rect 283840 157224 283892 157276
rect 335544 157224 335596 157276
rect 42432 157156 42484 157208
rect 151268 157156 151320 157208
rect 156512 157156 156564 157208
rect 159088 157156 159140 157208
rect 160100 157156 160152 157208
rect 166172 157156 166224 157208
rect 166264 157156 166316 157208
rect 171140 157156 171192 157208
rect 177028 157156 177080 157208
rect 254032 157156 254084 157208
rect 290556 157156 290608 157208
rect 340052 157156 340104 157208
rect 39028 157088 39080 157140
rect 148784 157088 148836 157140
rect 150072 157088 150124 157140
rect 233516 157088 233568 157140
rect 287152 157088 287204 157140
rect 338120 157088 338172 157140
rect 35716 157020 35768 157072
rect 146208 157020 146260 157072
rect 151728 157020 151780 157072
rect 234804 157020 234856 157072
rect 280436 157020 280488 157072
rect 333060 157020 333112 157072
rect 24768 156952 24820 157004
rect 137376 156952 137428 157004
rect 138296 156952 138348 157004
rect 224132 156952 224184 157004
rect 273720 156952 273772 157004
rect 327908 156952 327960 157004
rect 18052 156884 18104 156936
rect 132500 156884 132552 156936
rect 134892 156884 134944 156936
rect 214564 156884 214616 156936
rect 224960 156884 225012 156936
rect 272064 156884 272116 156936
rect 277124 156884 277176 156936
rect 330484 156884 330536 156936
rect 21364 156816 21416 156868
rect 135260 156816 135312 156868
rect 139124 156816 139176 156868
rect 225144 156816 225196 156868
rect 226616 156816 226668 156868
rect 291936 156816 291988 156868
rect 300676 156816 300728 156868
rect 348056 156816 348108 156868
rect 14648 156748 14700 156800
rect 130108 156748 130160 156800
rect 135812 156748 135864 156800
rect 222568 156748 222620 156800
rect 230020 156748 230072 156800
rect 294052 156748 294104 156800
rect 297272 156748 297324 156800
rect 345112 156748 345164 156800
rect 11244 156680 11296 156732
rect 127532 156680 127584 156732
rect 128176 156680 128228 156732
rect 216772 156680 216824 156732
rect 223212 156680 223264 156732
rect 289360 156680 289412 156732
rect 293868 156680 293920 156732
rect 342536 156680 342588 156732
rect 2044 156612 2096 156664
rect 120448 156612 120500 156664
rect 124864 156612 124916 156664
rect 213920 156612 213972 156664
rect 216496 156612 216548 156664
rect 283104 156612 283156 156664
rect 498292 156612 498344 156664
rect 499304 156612 499356 156664
rect 502340 156612 502392 156664
rect 503352 156612 503404 156664
rect 503720 156612 503772 156664
rect 505008 156612 505060 156664
rect 52460 156544 52512 156596
rect 158996 156544 159048 156596
rect 159088 156544 159140 156596
rect 200764 156544 200816 156596
rect 200948 156544 201000 156596
rect 270500 156544 270552 156596
rect 59268 156476 59320 156528
rect 164148 156476 164200 156528
rect 166172 156476 166224 156528
rect 69296 156408 69348 156460
rect 166264 156408 166316 156460
rect 166448 156476 166500 156528
rect 225052 156476 225104 156528
rect 228364 156408 228416 156460
rect 82820 156340 82872 156392
rect 182088 156340 182140 156392
rect 198832 156340 198884 156392
rect 200948 156340 201000 156392
rect 209780 156340 209832 156392
rect 279056 156340 279108 156392
rect 99564 156272 99616 156324
rect 194968 156272 195020 156324
rect 200764 156272 200816 156324
rect 101312 156204 101364 156256
rect 196256 156204 196308 156256
rect 197452 156204 197504 156256
rect 211620 156204 211672 156256
rect 108028 156136 108080 156188
rect 200672 156136 200724 156188
rect 118148 156068 118200 156120
rect 201040 156136 201092 156188
rect 201224 156136 201276 156188
rect 209136 156136 209188 156188
rect 213184 156272 213236 156324
rect 224224 156272 224276 156324
rect 214472 156204 214524 156256
rect 219992 156204 220044 156256
rect 220084 156204 220136 156256
rect 286232 156272 286284 156324
rect 215484 156136 215536 156188
rect 218060 156136 218112 156188
rect 266912 156204 266964 156256
rect 230756 156136 230808 156188
rect 277124 156136 277176 156188
rect 203064 156068 203116 156120
rect 273904 156068 273956 156120
rect 121460 156000 121512 156052
rect 197452 156000 197504 156052
rect 200948 156000 201000 156052
rect 201408 156000 201460 156052
rect 202236 156000 202288 156052
rect 273260 156000 273312 156052
rect 145012 155932 145064 155984
rect 229652 155932 229704 155984
rect 66812 155864 66864 155916
rect 82912 155864 82964 155916
rect 88708 155864 88760 155916
rect 186412 155864 186464 155916
rect 60096 155796 60148 155848
rect 79324 155796 79376 155848
rect 92020 155796 92072 155848
rect 189172 155864 189224 155916
rect 186780 155796 186832 155848
rect 194324 155864 194376 155916
rect 196348 155864 196400 155916
rect 268844 155864 268896 155916
rect 296444 155864 296496 155916
rect 345204 155864 345256 155916
rect 192944 155796 192996 155848
rect 266268 155796 266320 155848
rect 293040 155796 293092 155848
rect 342352 155796 342404 155848
rect 12164 155728 12216 155780
rect 110328 155728 110380 155780
rect 112260 155728 112312 155780
rect 204628 155728 204680 155780
rect 206468 155728 206520 155780
rect 276112 155728 276164 155780
rect 289728 155728 289780 155780
rect 339592 155728 339644 155780
rect 46572 155660 46624 155712
rect 75092 155660 75144 155712
rect 81900 155660 81952 155712
rect 180984 155660 181036 155712
rect 186228 155660 186280 155712
rect 260840 155660 260892 155712
rect 270316 155660 270368 155712
rect 325332 155660 325384 155712
rect 344376 155660 344428 155712
rect 381820 155660 381872 155712
rect 53380 155592 53432 155644
rect 66628 155592 66680 155644
rect 71872 155592 71924 155644
rect 172704 155592 172756 155644
rect 176292 155592 176344 155644
rect 253388 155592 253440 155644
rect 267004 155592 267056 155644
rect 322112 155592 322164 155644
rect 340972 155592 341024 155644
rect 378140 155592 378192 155644
rect 39856 155524 39908 155576
rect 68928 155524 68980 155576
rect 75184 155524 75236 155576
rect 176384 155524 176436 155576
rect 179512 155524 179564 155576
rect 255688 155524 255740 155576
rect 263600 155524 263652 155576
rect 320180 155524 320232 155576
rect 337660 155524 337712 155576
rect 375564 155524 375616 155576
rect 65156 155456 65208 155508
rect 168656 155456 168708 155508
rect 169392 155456 169444 155508
rect 248236 155456 248288 155508
rect 260288 155456 260340 155508
rect 317604 155456 317656 155508
rect 333428 155456 333480 155508
rect 373448 155456 373500 155508
rect 7932 155388 7984 155440
rect 124680 155388 124732 155440
rect 149244 155388 149296 155440
rect 232872 155388 232924 155440
rect 253572 155388 253624 155440
rect 312452 155388 312504 155440
rect 330116 155388 330168 155440
rect 370872 155388 370924 155440
rect 8760 155320 8812 155372
rect 125692 155320 125744 155372
rect 145840 155320 145892 155372
rect 229192 155320 229244 155372
rect 250168 155320 250220 155372
rect 309876 155320 309928 155372
rect 319996 155320 320048 155372
rect 363236 155320 363288 155372
rect 4528 155252 4580 155304
rect 122012 155252 122064 155304
rect 142528 155252 142580 155304
rect 227812 155252 227864 155304
rect 233332 155252 233384 155304
rect 297088 155252 297140 155304
rect 299756 155252 299808 155304
rect 347872 155252 347924 155304
rect 373816 155252 373868 155304
rect 404084 155252 404136 155304
rect 5356 155184 5408 155236
rect 123024 155184 123076 155236
rect 129004 155184 129056 155236
rect 217416 155184 217468 155236
rect 240048 155184 240100 155236
rect 302516 155184 302568 155236
rect 306564 155184 306616 155236
rect 352472 155184 352524 155236
rect 370412 155184 370464 155236
rect 401692 155184 401744 155236
rect 89536 155116 89588 155168
rect 187240 155116 187292 155168
rect 189632 155116 189684 155168
rect 263692 155116 263744 155168
rect 98736 155048 98788 155100
rect 186504 155048 186556 155100
rect 186872 155048 186924 155100
rect 191196 155048 191248 155100
rect 195980 155048 196032 155100
rect 196992 155048 197044 155100
rect 199660 155048 199712 155100
rect 271420 155048 271472 155100
rect 303160 155048 303212 155100
rect 350356 155048 350408 155100
rect 95424 154980 95476 155032
rect 190828 154980 190880 155032
rect 190920 154980 190972 155032
rect 200120 154980 200172 155032
rect 207020 154980 207072 155032
rect 269488 154980 269540 155032
rect 15476 154912 15528 154964
rect 109040 154912 109092 154964
rect 122288 154912 122340 154964
rect 190736 154912 190788 154964
rect 191012 154912 191064 154964
rect 211252 154912 211304 154964
rect 214656 154912 214708 154964
rect 261392 154912 261444 154964
rect 106372 154844 106424 154896
rect 190920 154844 190972 154896
rect 191196 154844 191248 154896
rect 245844 154844 245896 154896
rect 125784 154776 125836 154828
rect 214840 154776 214892 154828
rect 110512 154708 110564 154760
rect 139308 154708 139360 154760
rect 151820 154708 151872 154760
rect 153108 154708 153160 154760
rect 155960 154708 156012 154760
rect 238024 154708 238076 154760
rect 109132 154640 109184 154692
rect 133052 154640 133104 154692
rect 118608 154572 118660 154624
rect 119988 154572 120040 154624
rect 137100 154572 137152 154624
rect 138020 154572 138072 154624
rect 51080 154504 51132 154556
rect 142160 154572 142212 154624
rect 44180 154436 44232 154488
rect 142344 154436 142396 154488
rect 142436 154436 142488 154488
rect 157340 154640 157392 154692
rect 162676 154640 162728 154692
rect 243084 154640 243136 154692
rect 159364 154572 159416 154624
rect 240600 154572 240652 154624
rect 157248 154504 157300 154556
rect 212908 154504 212960 154556
rect 218336 154504 218388 154556
rect 190920 154436 190972 154488
rect 191012 154436 191064 154488
rect 201224 154436 201276 154488
rect 201316 154436 201368 154488
rect 207940 154436 207992 154488
rect 215300 154436 215352 154488
rect 283656 154504 283708 154556
rect 285588 154504 285640 154556
rect 285680 154504 285732 154556
rect 337476 154504 337528 154556
rect 353668 154504 353720 154556
rect 388904 154504 388956 154556
rect 283288 154436 283340 154488
rect 334900 154436 334952 154488
rect 349528 154436 349580 154488
rect 386328 154436 386380 154488
rect 390652 154436 390704 154488
rect 417148 154436 417200 154488
rect 114468 154368 114520 154420
rect 118608 154368 118660 154420
rect 118700 154368 118752 154420
rect 119896 154368 119948 154420
rect 119988 154368 120040 154420
rect 142620 154368 142672 154420
rect 189816 154368 189868 154420
rect 191196 154368 191248 154420
rect 202052 154368 202104 154420
rect 204996 154368 205048 154420
rect 275836 154368 275888 154420
rect 276204 154368 276256 154420
rect 329932 154368 329984 154420
rect 346400 154368 346452 154420
rect 383752 154368 383804 154420
rect 397368 154368 397420 154420
rect 422392 154368 422444 154420
rect 34520 154300 34572 154352
rect 142712 154300 142764 154352
rect 201132 154300 201184 154352
rect 201224 154300 201276 154352
rect 202696 154300 202748 154352
rect 208400 154300 208452 154352
rect 278412 154300 278464 154352
rect 278872 154300 278924 154352
rect 332416 154300 332468 154352
rect 343548 154300 343600 154352
rect 381176 154300 381228 154352
rect 393320 154300 393372 154352
rect 419724 154300 419776 154352
rect 37924 154232 37976 154284
rect 27252 154164 27304 154216
rect 136916 154164 136968 154216
rect 23480 154096 23532 154148
rect 137008 154096 137060 154148
rect 13820 154028 13872 154080
rect 129280 154028 129332 154080
rect 142160 154164 142212 154216
rect 142620 154232 142672 154284
rect 142896 154232 142948 154284
rect 150624 154232 150676 154284
rect 152372 154232 152424 154284
rect 163504 154232 163556 154284
rect 176660 154232 176712 154284
rect 179696 154232 179748 154284
rect 182180 154232 182232 154284
rect 258540 154232 258592 154284
rect 262220 154232 262272 154284
rect 319536 154232 319588 154284
rect 339500 154232 339552 154284
rect 378600 154232 378652 154284
rect 386512 154232 386564 154284
rect 414572 154232 414624 154284
rect 147588 154164 147640 154216
rect 147772 154164 147824 154216
rect 157248 154164 157300 154216
rect 157340 154164 157392 154216
rect 158352 154164 158404 154216
rect 161480 154164 161532 154216
rect 166080 154164 166132 154216
rect 172520 154164 172572 154216
rect 250812 154164 250864 154216
rect 255320 154164 255372 154216
rect 314384 154164 314436 154216
rect 336832 154164 336884 154216
rect 376024 154164 376076 154216
rect 383660 154164 383712 154216
rect 411996 154164 412048 154216
rect 9680 153960 9732 154012
rect 126888 153960 126940 154012
rect 127624 153960 127676 154012
rect 129372 153960 129424 154012
rect 7104 153892 7156 153944
rect 124312 153892 124364 153944
rect 125508 153892 125560 153944
rect 129648 153960 129700 154012
rect 142252 154096 142304 154148
rect 142620 154096 142672 154148
rect 145564 154096 145616 154148
rect 147128 154096 147180 154148
rect 137284 154028 137336 154080
rect 139768 154028 139820 154080
rect 139860 154028 139912 154080
rect 142436 154028 142488 154080
rect 142528 154028 142580 154080
rect 153200 154028 153252 154080
rect 153292 154028 153344 154080
rect 155960 154028 156012 154080
rect 160192 154096 160244 154148
rect 161572 154028 161624 154080
rect 165620 154096 165672 154148
rect 245660 154096 245712 154148
rect 245936 154096 245988 154148
rect 306656 154096 306708 154148
rect 326712 154096 326764 154148
rect 368296 154096 368348 154148
rect 376852 154096 376904 154148
rect 406844 154096 406896 154148
rect 241244 154028 241296 154080
rect 248604 154028 248656 154080
rect 309232 154028 309284 154080
rect 323308 154028 323360 154080
rect 365812 154028 365864 154080
rect 380164 154028 380216 154080
rect 409420 154028 409472 154080
rect 132408 153892 132460 153944
rect 219900 153960 219952 154012
rect 222384 153960 222436 154012
rect 288716 153960 288768 154012
rect 316040 153960 316092 154012
rect 360660 153960 360712 154012
rect 367100 153960 367152 154012
rect 399116 153960 399168 154012
rect 138020 153892 138072 153944
rect 480 153824 532 153876
rect 119804 153824 119856 153876
rect 119896 153824 119948 153876
rect 142804 153824 142856 153876
rect 142988 153892 143040 153944
rect 223212 153892 223264 153944
rect 225236 153892 225288 153944
rect 291292 153892 291344 153944
rect 313280 153892 313332 153944
rect 357900 153892 357952 153944
rect 363052 153892 363104 153944
rect 396540 153892 396592 153944
rect 401600 153892 401652 153944
rect 425520 153892 425572 153944
rect 152464 153824 152516 153876
rect 154488 153824 154540 153876
rect 48320 153756 48372 153808
rect 155776 153756 155828 153808
rect 155960 153824 156012 153876
rect 235448 153824 235500 153876
rect 241888 153824 241940 153876
rect 304080 153824 304132 153876
rect 309140 153824 309192 153876
rect 355508 153824 355560 153876
rect 356244 153824 356296 153876
rect 391480 153824 391532 153876
rect 397460 153824 397512 153876
rect 422944 153824 422996 153876
rect 218060 153756 218112 153808
rect 231860 153756 231912 153808
rect 296444 153756 296496 153808
rect 360384 153756 360436 153808
rect 394056 153756 394108 153808
rect 61108 153688 61160 153740
rect 161480 153688 161532 153740
rect 161572 153688 161624 153740
rect 210424 153688 210476 153740
rect 235080 153688 235132 153740
rect 299020 153688 299072 153740
rect 57980 153620 58032 153672
rect 152372 153620 152424 153672
rect 152464 153620 152516 153672
rect 191012 153620 191064 153672
rect 191748 153620 191800 153672
rect 195888 153620 195940 153672
rect 195980 153620 196032 153672
rect 209780 153620 209832 153672
rect 229100 153620 229152 153672
rect 293868 153620 293920 153672
rect 78680 153552 78732 153604
rect 179604 153552 179656 153604
rect 179696 153552 179748 153604
rect 230940 153552 230992 153604
rect 238852 153552 238904 153604
rect 301596 153552 301648 153604
rect 102140 153484 102192 153536
rect 196900 153484 196952 153536
rect 196992 153484 197044 153536
rect 200856 153484 200908 153536
rect 201132 153484 201184 153536
rect 205272 153484 205324 153536
rect 205364 153484 205416 153536
rect 248880 153484 248932 153536
rect 252652 153484 252704 153536
rect 311808 153484 311860 153536
rect 104900 153416 104952 153468
rect 199476 153416 199528 153468
rect 108304 153348 108356 153400
rect 191196 153348 191248 153400
rect 191288 153348 191340 153400
rect 197544 153348 197596 153400
rect 198924 153348 198976 153400
rect 200580 153348 200632 153400
rect 115940 153280 115992 153332
rect 207848 153416 207900 153468
rect 207940 153416 207992 153468
rect 259184 153416 259236 153468
rect 265440 153416 265492 153468
rect 322020 153416 322072 153468
rect 200764 153348 200816 153400
rect 205364 153348 205416 153400
rect 200856 153280 200908 153332
rect 243728 153348 243780 153400
rect 259460 153348 259512 153400
rect 316960 153348 317012 153400
rect 41604 153212 41656 153264
rect 142712 153212 142764 153264
rect 142804 153212 142856 153264
rect 195980 153212 196032 153264
rect 196072 153212 196124 153264
rect 238668 153280 238720 153332
rect 272892 153280 272944 153332
rect 327264 153280 327316 153332
rect 269212 153212 269264 153264
rect 324688 153212 324740 153264
rect 23296 153144 23348 153196
rect 110972 153144 111024 153196
rect 113180 153144 113232 153196
rect 205916 153144 205968 153196
rect 215392 153144 215444 153196
rect 279700 153144 279752 153196
rect 285496 153144 285548 153196
rect 336832 153144 336884 153196
rect 339684 153144 339736 153196
rect 377312 153144 377364 153196
rect 378232 153144 378284 153196
rect 379888 153144 379940 153196
rect 385500 153144 385552 153196
rect 387616 153144 387668 153196
rect 389180 153144 389232 153196
rect 393504 153144 393556 153196
rect 395528 153144 395580 153196
rect 397828 153144 397880 153196
rect 397920 153144 397972 153196
rect 415216 153144 415268 153196
rect 418160 153144 418212 153196
rect 437572 153144 437624 153196
rect 437848 153144 437900 153196
rect 446404 153144 446456 153196
rect 456800 153144 456852 153196
rect 459468 153144 459520 153196
rect 461860 153144 461912 153196
rect 465908 153144 465960 153196
rect 466460 153144 466512 153196
rect 470416 153144 470468 153196
rect 471520 153144 471572 153196
rect 473636 153144 473688 153196
rect 474832 153144 474884 153196
rect 476948 153144 477000 153196
rect 485688 153144 485740 153196
rect 489644 153144 489696 153196
rect 490748 153144 490800 153196
rect 493508 153144 493560 153196
rect 494060 153144 494112 153196
rect 496084 153144 496136 153196
rect 496636 153144 496688 153196
rect 498016 153144 498068 153196
rect 512276 153144 512328 153196
rect 514852 153144 514904 153196
rect 80060 153076 80112 153128
rect 175096 153076 175148 153128
rect 180800 153076 180852 153128
rect 257252 153076 257304 153128
rect 264980 153076 265032 153128
rect 321468 153076 321520 153128
rect 324320 153076 324372 153128
rect 367008 153076 367060 153128
rect 367192 153076 367244 153128
rect 368940 153076 368992 153128
rect 382188 153076 382240 153128
rect 410708 153076 410760 153128
rect 412916 153076 412968 153128
rect 422208 153076 422260 153128
rect 422300 153076 422352 153128
rect 423128 153076 423180 153128
rect 425152 153076 425204 153128
rect 434628 153076 434680 153128
rect 434720 153076 434772 153128
rect 443920 153076 443972 153128
rect 444012 153076 444064 153128
rect 450544 153076 450596 153128
rect 462780 153076 462832 153128
rect 466552 153076 466604 153128
rect 466644 153076 466696 153128
rect 469772 153076 469824 153128
rect 472256 153076 472308 153128
rect 474280 153076 474332 153128
rect 476120 153076 476172 153128
rect 478144 153076 478196 153128
rect 484032 153076 484084 153128
rect 488448 153076 488500 153128
rect 492404 153076 492456 153128
rect 494796 153076 494848 153128
rect 494980 153076 495032 153128
rect 496728 153076 496780 153128
rect 496820 153076 496872 153128
rect 498660 153076 498712 153128
rect 510988 153076 511040 153128
rect 513472 153076 513524 153128
rect 513564 153076 513616 153128
rect 516140 153076 516192 153128
rect 103520 153008 103572 153060
rect 198188 153008 198240 153060
rect 203708 153008 203760 153060
rect 267556 153008 267608 153060
rect 272156 153008 272208 153060
rect 326620 153008 326672 153060
rect 330944 153008 330996 153060
rect 371516 153008 371568 153060
rect 372620 153008 372672 153060
rect 403624 153008 403676 153060
rect 405832 153008 405884 153060
rect 408776 153008 408828 153060
rect 410524 153008 410576 153060
rect 431132 153008 431184 153060
rect 431960 153008 432012 153060
rect 441988 153008 442040 153060
rect 442080 153008 442132 153060
rect 447416 153008 447468 153060
rect 463148 153008 463200 153060
rect 467196 153008 467248 153060
rect 472624 153008 472676 153060
rect 474924 153008 474976 153060
rect 484492 153008 484544 153060
rect 489000 153008 489052 153060
rect 492680 153008 492732 153060
rect 495440 153008 495492 153060
rect 495532 153008 495584 153060
rect 497372 153008 497424 153060
rect 511632 153008 511684 153060
rect 514300 153008 514352 153060
rect 92572 152940 92624 152992
rect 187884 152940 187936 152992
rect 195060 152940 195112 152992
rect 218704 152940 218756 152992
rect 220360 152940 220412 152992
rect 284852 152940 284904 152992
rect 288072 152940 288124 152992
rect 290004 152940 290056 152992
rect 292212 152940 292264 152992
rect 341984 152940 342036 152992
rect 342260 152940 342312 152992
rect 343916 152940 343968 152992
rect 345296 152940 345348 152992
rect 382464 152940 382516 152992
rect 384948 152940 385000 152992
rect 392124 152940 392176 152992
rect 394884 152940 394936 152992
rect 415308 152940 415360 152992
rect 415400 152940 415452 152992
rect 71412 152872 71464 152924
rect 92480 152872 92532 152924
rect 96620 152872 96672 152924
rect 193036 152872 193088 152924
rect 212448 152872 212500 152924
rect 277768 152872 277820 152924
rect 278780 152872 278832 152924
rect 331772 152872 331824 152924
rect 332600 152872 332652 152924
rect 372804 152872 372856 152924
rect 375472 152872 375524 152924
rect 405556 152872 405608 152924
rect 406660 152872 406712 152924
rect 417608 152872 417660 152924
rect 421012 152940 421064 152992
rect 436376 152872 436428 152924
rect 437572 152940 437624 152992
rect 438308 152940 438360 152992
rect 439044 152940 439096 152992
rect 440332 152940 440384 152992
rect 455696 152940 455748 152992
rect 464160 152940 464212 152992
rect 467840 152940 467892 152992
rect 471428 152940 471480 152992
rect 472992 152940 473044 152992
rect 473360 152940 473412 152992
rect 475568 152940 475620 152992
rect 483112 152940 483164 152992
rect 487804 152940 487856 152992
rect 491576 152940 491628 152992
rect 494152 152940 494204 152992
rect 512920 152940 512972 152992
rect 515956 152940 516008 152992
rect 438860 152872 438912 152924
rect 454408 152872 454460 152924
rect 464436 152872 464488 152924
rect 468392 152872 468444 152924
rect 489920 152872 489972 152924
rect 492864 152872 492916 152924
rect 514208 152872 514260 152924
rect 517428 152872 517480 152924
rect 33140 152804 33192 152856
rect 138020 152804 138072 152856
rect 138112 152804 138164 152856
rect 141700 152804 141752 152856
rect 146576 152804 146628 152856
rect 167368 152804 167420 152856
rect 173900 152804 173952 152856
rect 252100 152804 252152 152856
rect 255412 152804 255464 152856
rect 313096 152804 313148 152856
rect 317052 152804 317104 152856
rect 318248 152804 318300 152856
rect 320272 152804 320324 152856
rect 323124 152804 323176 152856
rect 324228 152804 324280 152856
rect 366364 152804 366416 152856
rect 371332 152804 371384 152856
rect 402336 152804 402388 152856
rect 411260 152804 411312 152856
rect 433156 152804 433208 152856
rect 434352 152804 434404 152856
rect 444012 152804 444064 152856
rect 26424 152736 26476 152788
rect 139124 152736 139176 152788
rect 140780 152736 140832 152788
rect 144276 152736 144328 152788
rect 144368 152736 144420 152788
rect 162216 152736 162268 152788
rect 164424 152736 164476 152788
rect 244372 152736 244424 152788
rect 257712 152736 257764 152788
rect 315672 152736 315724 152788
rect 317420 152736 317472 152788
rect 361304 152736 361356 152788
rect 361580 152736 361632 152788
rect 395344 152736 395396 152788
rect 398840 152736 398892 152788
rect 403808 152736 403860 152788
rect 404360 152736 404412 152788
rect 428004 152736 428056 152788
rect 429292 152736 429344 152788
rect 446680 152804 446732 152856
rect 446772 152804 446824 152856
rect 452476 152804 452528 152856
rect 465080 152804 465132 152856
rect 469128 152804 469180 152856
rect 510344 152804 510396 152856
rect 512000 152804 512052 152856
rect 444472 152736 444524 152788
rect 28172 152668 28224 152720
rect 141056 152668 141108 152720
rect 142804 152668 142856 152720
rect 149428 152668 149480 152720
rect 149520 152668 149572 152720
rect 231584 152668 231636 152720
rect 240324 152668 240376 152720
rect 241888 152668 241940 152720
rect 251180 152668 251232 152720
rect 311164 152668 311216 152720
rect 312176 152668 312228 152720
rect 356152 152668 356204 152720
rect 358820 152668 358872 152720
rect 393412 152668 393464 152720
rect 393504 152668 393556 152720
rect 398104 152668 398156 152720
rect 399208 152668 399260 152720
rect 417332 152668 417384 152720
rect 22192 152600 22244 152652
rect 135904 152600 135956 152652
rect 19340 152532 19392 152584
rect 133972 152532 134024 152584
rect 136640 152532 136692 152584
rect 151912 152600 151964 152652
rect 153568 152600 153620 152652
rect 236736 152600 236788 152652
rect 247040 152600 247092 152652
rect 307944 152600 307996 152652
rect 311532 152600 311584 152652
rect 320824 152600 320876 152652
rect 320916 152600 320968 152652
rect 361948 152600 362000 152652
rect 368480 152600 368532 152652
rect 400404 152600 400456 152652
rect 138112 152532 138164 152584
rect 144276 152532 144328 152584
rect 144368 152532 144420 152584
rect 226432 152532 226484 152584
rect 234160 152532 234212 152584
rect 297732 152532 297784 152584
rect 303620 152532 303672 152584
rect 351000 152532 351052 152584
rect 351920 152532 351972 152584
rect 353484 152532 353536 152584
rect 354496 152532 354548 152584
rect 389548 152532 389600 152584
rect 390376 152532 390428 152584
rect 397920 152532 397972 152584
rect 398012 152532 398064 152584
rect 403348 152532 403400 152584
rect 2872 152464 2924 152516
rect 121092 152464 121144 152516
rect 126980 152464 127032 152516
rect 216128 152464 216180 152516
rect 227720 152464 227772 152516
rect 293224 152464 293276 152516
rect 298652 152464 298704 152516
rect 347136 152464 347188 152516
rect 348148 152464 348200 152516
rect 385040 152464 385092 152516
rect 386420 152464 386472 152516
rect 413928 152600 413980 152652
rect 414020 152600 414072 152652
rect 421656 152668 421708 152720
rect 417608 152600 417660 152652
rect 421748 152600 421800 152652
rect 403532 152532 403584 152584
rect 419080 152532 419132 152584
rect 426348 152668 426400 152720
rect 426440 152668 426492 152720
rect 444748 152668 444800 152720
rect 444932 152736 444984 152788
rect 451188 152736 451240 152788
rect 458180 152668 458232 152720
rect 421932 152600 421984 152652
rect 66628 152396 66680 152448
rect 159640 152396 159692 152448
rect 173164 152396 173216 152448
rect 249524 152396 249576 152448
rect 260932 152396 260984 152448
rect 316316 152396 316368 152448
rect 317512 152396 317564 152448
rect 320640 152396 320692 152448
rect 320732 152396 320784 152448
rect 325976 152396 326028 152448
rect 326068 152396 326120 152448
rect 367652 152396 367704 152448
rect 380992 152396 381044 152448
rect 410064 152464 410116 152516
rect 413836 152464 413888 152516
rect 416504 152464 416556 152516
rect 418620 152464 418672 152516
rect 419540 152464 419592 152516
rect 421932 152464 421984 152516
rect 403716 152396 403768 152448
rect 412640 152396 412692 152448
rect 415308 152396 415360 152448
rect 420368 152396 420420 152448
rect 33600 152328 33652 152380
rect 109684 152328 109736 152380
rect 109776 152328 109828 152380
rect 110512 152328 110564 152380
rect 120080 152328 120132 152380
rect 211068 152328 211120 152380
rect 224408 152328 224460 152380
rect 288072 152328 288124 152380
rect 291384 152328 291436 152380
rect 341340 152328 341392 152380
rect 343824 152328 343876 152380
rect 349804 152328 349856 152380
rect 349896 152328 349948 152380
rect 385684 152328 385736 152380
rect 386236 152328 386288 152380
rect 399760 152328 399812 152380
rect 402428 152328 402480 152380
rect 426072 152532 426124 152584
rect 429200 152600 429252 152652
rect 429384 152600 429436 152652
rect 426532 152532 426584 152584
rect 438952 152532 439004 152584
rect 439044 152532 439096 152584
rect 440884 152532 440936 152584
rect 441988 152600 442040 152652
rect 446128 152600 446180 152652
rect 446404 152600 446456 152652
rect 453764 152600 453816 152652
rect 447324 152532 447376 152584
rect 447416 152532 447468 152584
rect 456984 152532 457036 152584
rect 422852 152464 422904 152516
rect 435732 152464 435784 152516
rect 436928 152464 436980 152516
rect 446772 152464 446824 152516
rect 459560 152464 459612 152516
rect 464620 152464 464672 152516
rect 422208 152396 422260 152448
rect 423036 152396 423088 152448
rect 442172 152396 442224 152448
rect 443000 152396 443052 152448
rect 457628 152396 457680 152448
rect 424416 152328 424468 152380
rect 424508 152328 424560 152380
rect 426900 152328 426952 152380
rect 427820 152328 427872 152380
rect 446036 152328 446088 152380
rect 446128 152328 446180 152380
rect 449256 152328 449308 152380
rect 91100 152260 91152 152312
rect 180248 152260 180300 152312
rect 187976 152260 188028 152312
rect 262404 152260 262456 152312
rect 266360 152260 266412 152312
rect 320916 152260 320968 152312
rect 331220 152260 331272 152312
rect 372160 152260 372212 152312
rect 382280 152260 382332 152312
rect 386972 152260 387024 152312
rect 393136 152260 393188 152312
rect 398012 152260 398064 152312
rect 398104 152260 398156 152312
rect 403716 152260 403768 152312
rect 403808 152260 403860 152312
rect 413284 152260 413336 152312
rect 414296 152260 414348 152312
rect 422852 152260 422904 152312
rect 423128 152260 423180 152312
rect 441528 152260 441580 152312
rect 441620 152260 441672 152312
rect 456340 152260 456392 152312
rect 19800 152192 19852 152244
rect 97908 152192 97960 152244
rect 109040 152192 109092 152244
rect 130752 152192 130804 152244
rect 134064 152192 134116 152244
rect 221280 152192 221332 152244
rect 222108 152192 222160 152244
rect 282920 152192 282972 152244
rect 285772 152192 285824 152244
rect 336188 152192 336240 152244
rect 342444 152192 342496 152244
rect 344560 152192 344612 152244
rect 349160 152192 349212 152244
rect 349896 152192 349948 152244
rect 352012 152192 352064 152244
rect 388260 152192 388312 152244
rect 394332 152192 394384 152244
rect 417792 152192 417844 152244
rect 417884 152192 417936 152244
rect 424324 152192 424376 152244
rect 425980 152192 426032 152244
rect 444104 152192 444156 152244
rect 445300 152192 445352 152244
rect 458824 152192 458876 152244
rect 9496 152124 9548 152176
rect 82820 152124 82872 152176
rect 82912 152124 82964 152176
rect 169944 152124 169996 152176
rect 172152 152124 172204 152176
rect 190460 152124 190512 152176
rect 193588 152124 193640 152176
rect 213552 152124 213604 152176
rect 225328 152124 225380 152176
rect 229008 152124 229060 152176
rect 244464 152124 244516 152176
rect 306012 152124 306064 152176
rect 320824 152124 320876 152176
rect 356796 152124 356848 152176
rect 357532 152124 357584 152176
rect 359372 152124 359424 152176
rect 365720 152124 365772 152176
rect 398472 152124 398524 152176
rect 398564 152124 398616 152176
rect 408132 152124 408184 152176
rect 409236 152124 409288 152176
rect 428648 152124 428700 152176
rect 430672 152124 430724 152176
rect 447968 152124 448020 152176
rect 79324 152056 79376 152108
rect 164792 152056 164844 152108
rect 167000 152056 167052 152108
rect 182732 152056 182784 152108
rect 183468 152056 183520 152108
rect 200764 152056 200816 152108
rect 213828 152056 213880 152108
rect 274548 152056 274600 152108
rect 277400 152056 277452 152108
rect 331128 152056 331180 152108
rect 335360 152056 335412 152108
rect 375380 152056 375432 152108
rect 378784 152056 378836 152108
rect 384396 152056 384448 152108
rect 388444 152056 388496 152108
rect 407488 152056 407540 152108
rect 408500 152056 408552 152108
rect 423588 152056 423640 152108
rect 424416 152056 424468 152108
rect 433800 152056 433852 152108
rect 433892 152056 433944 152108
rect 449900 152056 449952 152108
rect 516692 152056 516744 152108
rect 520280 152056 520332 152108
rect 68928 151988 68980 152040
rect 142804 151988 142856 152040
rect 143172 151988 143224 152040
rect 146944 151988 146996 152040
rect 156328 151988 156380 152040
rect 172520 151988 172572 152040
rect 191472 151988 191524 152040
rect 208492 151988 208544 152040
rect 242440 151988 242492 152040
rect 300952 151988 301004 152040
rect 304172 151988 304224 152040
rect 351644 151988 351696 152040
rect 354680 151988 354732 152040
rect 390192 151988 390244 152040
rect 75092 151920 75144 151972
rect 154488 151920 154540 151972
rect 162492 151920 162544 151972
rect 177672 151920 177724 151972
rect 184388 151920 184440 151972
rect 195612 151920 195664 151972
rect 243360 151920 243412 151972
rect 302884 151920 302936 151972
rect 307668 151920 307720 151972
rect 352288 151920 352340 151972
rect 364616 151920 364668 151972
rect 397184 151988 397236 152040
rect 404912 151988 404964 152040
rect 405372 151988 405424 152040
rect 421012 151988 421064 152040
rect 30196 151852 30248 151904
rect 110328 151852 110380 151904
rect 110512 151852 110564 151904
rect 138480 151852 138532 151904
rect 139308 151852 139360 151904
rect 203340 151852 203392 151904
rect 212632 151852 212684 151904
rect 272708 151852 272760 151904
rect 74816 151784 74868 151836
rect 81348 151784 81400 151836
rect 105820 151784 105872 151836
rect 110236 151784 110288 151836
rect 110420 151784 110472 151836
rect 128176 151784 128228 151836
rect 129740 151784 129792 151836
rect 146852 151784 146904 151836
rect 146944 151784 146996 151836
rect 157064 151784 157116 151836
rect 169760 151784 169812 151836
rect 185308 151784 185360 151836
rect 271880 151784 271932 151836
rect 320732 151852 320784 151904
rect 321560 151852 321612 151904
rect 362592 151852 362644 151904
rect 363144 151852 363196 151904
rect 364524 151852 364576 151904
rect 388168 151852 388220 151904
rect 404176 151920 404228 151972
rect 418436 151920 418488 151972
rect 419632 151920 419684 151972
rect 434444 151988 434496 152040
rect 434628 151988 434680 152040
rect 443460 151988 443512 152040
rect 446312 151988 446364 152040
rect 460020 151988 460072 152040
rect 485780 151988 485832 152040
rect 490288 151988 490340 152040
rect 423220 151920 423272 151972
rect 439596 151920 439648 151972
rect 440240 151920 440292 151972
rect 455052 151920 455104 151972
rect 469220 151920 469272 151972
rect 472348 151920 472400 151972
rect 488540 151920 488592 151972
rect 492220 151920 492272 151972
rect 509056 151920 509108 151972
rect 510896 151920 510948 151972
rect 517428 151920 517480 151972
rect 521568 151920 521620 151972
rect 396172 151852 396224 151904
rect 402980 151852 403032 151904
rect 416596 151852 416648 151904
rect 426808 151852 426860 151904
rect 426900 151852 426952 151904
rect 437020 151852 437072 151904
rect 437480 151852 437532 151904
rect 453120 151852 453172 151904
rect 468024 151852 468076 151904
rect 471060 151852 471112 151904
rect 487344 151852 487396 151904
rect 490932 151852 490984 151904
rect 507768 151852 507820 151904
rect 509516 151852 509568 151904
rect 516048 151852 516100 151904
rect 519912 151852 519964 151904
rect 283196 151784 283248 151836
rect 287428 151784 287480 151836
rect 300400 151784 300452 151836
rect 81716 151716 81768 151768
rect 112812 151716 112864 151768
rect 346492 151784 346544 151836
rect 349804 151784 349856 151836
rect 380532 151784 380584 151836
rect 386144 151784 386196 151836
rect 394700 151784 394752 151836
rect 404268 151784 404320 151836
rect 415860 151784 415912 151836
rect 417332 151784 417384 151836
rect 424232 151784 424284 151836
rect 424324 151784 424376 151836
rect 431868 151784 431920 151836
rect 436100 151784 436152 151836
rect 451832 151784 451884 151836
rect 467932 151784 467984 151836
rect 471704 151784 471756 151836
rect 488172 151784 488224 151836
rect 491576 151784 491628 151836
rect 499120 151784 499172 151836
rect 499948 151784 500000 151836
rect 515496 151784 515548 151836
rect 518992 151784 519044 151836
rect 43904 151648 43956 151700
rect 111432 151648 111484 151700
rect 40500 151580 40552 151632
rect 111340 151580 111392 151632
rect 37004 151512 37056 151564
rect 111064 151512 111116 151564
rect 26700 151444 26752 151496
rect 116952 151444 117004 151496
rect 16396 151376 16448 151428
rect 116768 151376 116820 151428
rect 12992 151308 13044 151360
rect 116676 151308 116728 151360
rect 68008 151240 68060 151292
rect 112720 151240 112772 151292
rect 64512 151172 64564 151224
rect 112628 151172 112680 151224
rect 61108 151104 61160 151156
rect 112536 151104 112588 151156
rect 57704 151036 57756 151088
rect 111708 151036 111760 151088
rect 54208 150968 54260 151020
rect 112444 150968 112496 151020
rect 50804 150900 50856 150952
rect 111616 150900 111668 150952
rect 47308 150832 47360 150884
rect 111524 150832 111576 150884
rect 98920 150764 98972 150816
rect 116032 150764 116084 150816
rect 95516 150696 95568 150748
rect 115296 150696 115348 150748
rect 92020 150628 92072 150680
rect 113088 150628 113140 150680
rect 88616 150560 88668 150612
rect 112996 150560 113048 150612
rect 85212 150492 85264 150544
rect 115204 150492 115256 150544
rect 102324 150424 102376 150476
rect 116124 150424 116176 150476
rect 78312 150288 78364 150340
rect 112904 150288 112956 150340
rect 110328 150220 110380 150272
rect 117136 150220 117188 150272
rect 97908 150152 97960 150204
rect 116860 150152 116912 150204
rect 122840 150152 122892 150204
rect 123714 150152 123766 150204
rect 146392 150152 146444 150204
rect 147542 150152 147594 150204
rect 164332 150152 164384 150204
rect 165482 150152 165534 150204
rect 168380 150152 168432 150204
rect 169346 150152 169398 150204
rect 171140 150152 171192 150204
rect 171922 150152 171974 150204
rect 172704 150152 172756 150204
rect 173854 150152 173906 150204
rect 182272 150152 182324 150204
rect 183422 150152 183474 150204
rect 190828 150152 190880 150204
rect 191794 150152 191846 150204
rect 211252 150152 211304 150204
rect 212310 150152 212362 150204
rect 225052 150152 225104 150204
rect 225834 150152 225886 150204
rect 229192 150152 229244 150204
rect 230342 150152 230394 150204
rect 233240 150152 233292 150204
rect 234206 150152 234258 150204
rect 238944 150152 238996 150204
rect 240002 150152 240054 150204
rect 253940 150152 253992 150204
rect 254722 150152 254774 150204
rect 256792 150152 256844 150204
rect 257942 150152 257994 150204
rect 263600 150152 263652 150204
rect 264382 150152 264434 150204
rect 269120 150152 269172 150204
rect 270178 150152 270230 150204
rect 281540 150152 281592 150204
rect 282322 150152 282374 150204
rect 283104 150152 283156 150204
rect 284254 150152 284306 150204
rect 284392 150152 284444 150204
rect 285542 150152 285594 150204
rect 299480 150152 299532 150204
rect 300354 150152 300406 150204
rect 332692 150152 332744 150204
rect 333750 150152 333802 150204
rect 338304 150152 338356 150204
rect 339454 150152 339506 150204
rect 345112 150152 345164 150204
rect 345894 150152 345946 150204
rect 358912 150152 358964 150204
rect 360062 150152 360114 150204
rect 362960 150152 363012 150204
rect 363926 150152 363978 150204
rect 374000 150152 374052 150204
rect 374782 150152 374834 150204
rect 375564 150152 375616 150204
rect 376714 150152 376766 150204
rect 378140 150152 378192 150204
rect 379290 150152 379342 150204
rect 460940 150152 460992 150204
rect 462090 150152 462142 150204
rect 477684 150152 477736 150204
rect 478834 150152 478886 150204
rect 483204 150152 483256 150204
rect 483986 150152 484038 150204
rect 502340 150152 502392 150204
rect 503214 150152 503266 150204
rect 503720 150152 503772 150204
rect 504502 150152 504554 150204
rect 505284 150152 505336 150204
rect 506434 150152 506486 150204
rect 518026 150152 518078 150204
rect 518808 150152 518860 150204
rect 81348 150084 81400 150136
rect 92480 150084 92532 150136
rect 117228 150084 117280 150136
rect 116492 150016 116544 150068
rect 111156 148384 111208 148436
rect 117044 148316 117096 148368
rect 113088 140700 113140 140752
rect 116124 140700 116176 140752
rect 112996 137912 113048 137964
rect 116124 137912 116176 137964
rect 112812 133832 112864 133884
rect 116032 133832 116084 133884
rect 114192 132608 114244 132660
rect 115204 132608 115256 132660
rect 112904 132404 112956 132456
rect 116124 132404 116176 132456
rect 112720 126896 112772 126948
rect 116124 126896 116176 126948
rect 112628 124108 112680 124160
rect 116124 124108 116176 124160
rect 112536 122748 112588 122800
rect 115940 122748 115992 122800
rect 111708 121388 111760 121440
rect 116124 121388 116176 121440
rect 112444 118600 112496 118652
rect 116124 118600 116176 118652
rect 111616 117240 111668 117292
rect 116124 117240 116176 117292
rect 111524 114452 111576 114504
rect 116124 114452 116176 114504
rect 111432 113092 111484 113144
rect 115940 113092 115992 113144
rect 111340 111732 111392 111784
rect 116124 111732 116176 111784
rect 111156 108944 111208 108996
rect 116124 108944 116176 108996
rect 111248 92420 111300 92472
rect 116124 92420 116176 92472
rect 111064 89632 111116 89684
rect 116124 89632 116176 89684
rect 113824 88272 113876 88324
rect 116032 88272 116084 88324
rect 113916 83920 113968 83972
rect 116584 83920 116636 83972
rect 114008 82764 114060 82816
rect 116216 82764 116268 82816
rect 114100 79976 114152 80028
rect 115940 79976 115992 80028
rect 114192 78616 114244 78668
rect 116124 78616 116176 78668
rect 114192 71748 114244 71800
rect 116584 71748 116636 71800
rect 114100 69028 114152 69080
rect 116308 69028 116360 69080
rect 114008 67600 114060 67652
rect 116124 67600 116176 67652
rect 113916 66240 113968 66292
rect 116584 66240 116636 66292
rect 113364 64676 113416 64728
rect 116584 64676 116636 64728
rect 113824 63520 113876 63572
rect 116216 63520 116268 63572
rect 112444 62092 112496 62144
rect 116124 62092 116176 62144
rect 112536 42780 112588 42832
rect 116124 42780 116176 42832
rect 116676 7896 116728 7948
rect 116860 7896 116912 7948
rect 117044 7760 117096 7812
rect 117320 7760 117372 7812
rect 116860 7692 116912 7744
rect 116768 7624 116820 7676
rect 117228 7624 117280 7676
rect 117044 7420 117096 7472
rect 111708 2796 111760 2848
rect 193588 2456 193640 2508
rect 425796 2456 425848 2508
rect 443644 2456 443696 2508
rect 62396 1844 62448 1896
rect 65340 1844 65392 1896
rect 68008 1844 68060 1896
rect 89260 1844 89312 1896
rect 89352 1844 89404 1896
rect 97172 1844 97224 1896
rect 104348 1844 104400 1896
rect 64144 1776 64196 1828
rect 69388 1776 69440 1828
rect 75644 1776 75696 1828
rect 85396 1776 85448 1828
rect 86040 1776 86092 1828
rect 111064 1912 111116 1964
rect 104532 1844 104584 1896
rect 105728 1844 105780 1896
rect 105820 1844 105872 1896
rect 105912 1844 105964 1896
rect 109224 1844 109276 1896
rect 109316 1844 109368 1896
rect 62672 1708 62724 1760
rect 77208 1708 77260 1760
rect 82636 1708 82688 1760
rect 104072 1708 104124 1760
rect 109592 1776 109644 1828
rect 109960 1708 110012 1760
rect 112444 1708 112496 1760
rect 69296 1640 69348 1692
rect 102600 1640 102652 1692
rect 102692 1640 102744 1692
rect 105820 1640 105872 1692
rect 106188 1640 106240 1692
rect 116584 1640 116636 1692
rect 59360 1572 59412 1624
rect 68468 1572 68520 1624
rect 79324 1572 79376 1624
rect 97264 1572 97316 1624
rect 99380 1572 99432 1624
rect 105912 1572 105964 1624
rect 106004 1572 106056 1624
rect 110052 1572 110104 1624
rect 72700 1504 72752 1556
rect 110512 1504 110564 1556
rect 42616 1436 42668 1488
rect 68284 1436 68336 1488
rect 87972 1436 88024 1488
rect 97172 1436 97224 1488
rect 97264 1436 97316 1488
rect 108212 1436 108264 1488
rect 108304 1436 108356 1488
rect 143632 1436 143684 1488
rect 46020 1368 46072 1420
rect 116492 1368 116544 1420
rect 55956 1300 56008 1352
rect 294788 1368 294840 1420
rect 343640 1368 343692 1420
rect 491300 1368 491352 1420
rect 493600 1368 493652 1420
rect 2688 1232 2740 1284
rect 116308 1232 116360 1284
rect 39304 1164 39356 1216
rect 116400 1164 116452 1216
rect 49332 1096 49384 1148
rect 116768 1096 116820 1148
rect 52644 1028 52696 1080
rect 117228 1028 117280 1080
rect 65984 960 66036 1012
rect 116860 960 116912 1012
rect 76012 892 76064 944
rect 112536 892 112588 944
rect 91744 824 91796 876
rect 99748 824 99800 876
rect 103888 824 103940 876
rect 108304 824 108356 876
rect 95700 756 95752 808
rect 99564 756 99616 808
<< metal2 >>
rect 386 163200 442 164400
rect 492 163254 1164 163282
rect 400 158030 428 163200
rect 388 158024 440 158030
rect 388 157966 440 157972
rect 492 153882 520 163254
rect 1136 163146 1164 163254
rect 1214 163200 1270 164400
rect 2042 163200 2098 164400
rect 2870 163200 2926 164400
rect 2976 163254 3648 163282
rect 1228 163146 1256 163200
rect 1136 163118 1256 163146
rect 2056 156670 2084 163200
rect 2044 156664 2096 156670
rect 2044 156606 2096 156612
rect 480 153876 532 153882
rect 480 153818 532 153824
rect 2884 152522 2912 163200
rect 2976 153785 3004 163254
rect 3620 163146 3648 163254
rect 3698 163200 3754 164400
rect 4526 163200 4582 164400
rect 5354 163200 5410 164400
rect 6274 163200 6330 164400
rect 7102 163200 7158 164400
rect 7930 163200 7986 164400
rect 8758 163200 8814 164400
rect 8864 163254 9536 163282
rect 3712 163146 3740 163200
rect 3620 163118 3740 163146
rect 4540 155310 4568 163200
rect 4528 155304 4580 155310
rect 4528 155246 4580 155252
rect 5368 155242 5396 163200
rect 6288 159390 6316 163200
rect 6276 159384 6328 159390
rect 6276 159326 6328 159332
rect 5356 155236 5408 155242
rect 5356 155178 5408 155184
rect 7116 153950 7144 163200
rect 7944 155446 7972 163200
rect 7932 155440 7984 155446
rect 7932 155382 7984 155388
rect 8772 155378 8800 163200
rect 8760 155372 8812 155378
rect 8760 155314 8812 155320
rect 7104 153944 7156 153950
rect 7104 153886 7156 153892
rect 2962 153776 3018 153785
rect 2962 153711 3018 153720
rect 2872 152516 2924 152522
rect 2872 152458 2924 152464
rect 8864 152425 8892 163254
rect 9508 163146 9536 163254
rect 9586 163200 9642 164400
rect 9692 163254 10364 163282
rect 9600 163146 9628 163200
rect 9508 163118 9628 163146
rect 9692 154018 9720 163254
rect 10336 163146 10364 163254
rect 10414 163200 10470 164400
rect 11242 163200 11298 164400
rect 12162 163200 12218 164400
rect 12452 163254 12940 163282
rect 10428 163146 10456 163200
rect 10336 163118 10456 163146
rect 11256 156738 11284 163200
rect 11244 156732 11296 156738
rect 11244 156674 11296 156680
rect 12176 155786 12204 163200
rect 12164 155780 12216 155786
rect 12164 155722 12216 155728
rect 9680 154012 9732 154018
rect 9680 153954 9732 153960
rect 12452 152561 12480 163254
rect 12912 163146 12940 163254
rect 12990 163200 13046 164400
rect 13818 163200 13874 164400
rect 14646 163200 14702 164400
rect 15474 163200 15530 164400
rect 16302 163200 16358 164400
rect 16592 163254 17080 163282
rect 13004 163146 13032 163200
rect 12912 163118 13032 163146
rect 13832 154086 13860 163200
rect 14660 156806 14688 163200
rect 14648 156800 14700 156806
rect 14648 156742 14700 156748
rect 15488 154970 15516 163200
rect 16316 159361 16344 163200
rect 16302 159352 16358 159361
rect 16302 159287 16358 159296
rect 15476 154964 15528 154970
rect 15476 154906 15528 154912
rect 13820 154080 13872 154086
rect 13820 154022 13872 154028
rect 16592 153921 16620 163254
rect 17052 163146 17080 163254
rect 17130 163200 17186 164400
rect 18050 163200 18106 164400
rect 18878 163200 18934 164400
rect 19352 163254 19656 163282
rect 17144 163146 17172 163200
rect 17052 163118 17172 163146
rect 18064 156942 18092 163200
rect 18892 159730 18920 163200
rect 18880 159724 18932 159730
rect 18880 159666 18932 159672
rect 18052 156936 18104 156942
rect 18052 156878 18104 156884
rect 16578 153912 16634 153921
rect 16578 153847 16634 153856
rect 19352 152590 19380 163254
rect 19628 163146 19656 163254
rect 19706 163200 19762 164400
rect 19904 163254 20484 163282
rect 19720 163146 19748 163200
rect 19628 163118 19748 163146
rect 19904 154057 19932 163254
rect 20456 163146 20484 163254
rect 20534 163200 20590 164400
rect 21362 163200 21418 164400
rect 22190 163200 22246 164400
rect 23018 163200 23074 164400
rect 23492 163254 23888 163282
rect 20548 163146 20576 163200
rect 20456 163118 20576 163146
rect 21376 156874 21404 163200
rect 21364 156868 21416 156874
rect 21364 156810 21416 156816
rect 19890 154048 19946 154057
rect 19890 153983 19946 153992
rect 22204 152658 22232 163200
rect 23032 159497 23060 163200
rect 23018 159488 23074 159497
rect 23018 159423 23074 159432
rect 23492 154154 23520 163254
rect 23860 163146 23888 163254
rect 23938 163200 23994 164400
rect 24766 163200 24822 164400
rect 25594 163200 25650 164400
rect 26422 163200 26478 164400
rect 27250 163200 27306 164400
rect 28078 163200 28134 164400
rect 28184 163254 28856 163282
rect 23952 163146 23980 163200
rect 23860 163118 23980 163146
rect 24780 157010 24808 163200
rect 25608 160002 25636 163200
rect 25596 159996 25648 160002
rect 25596 159938 25648 159944
rect 24768 157004 24820 157010
rect 24768 156946 24820 156952
rect 23480 154148 23532 154154
rect 23480 154090 23532 154096
rect 23296 153196 23348 153202
rect 23296 153138 23348 153144
rect 22192 152652 22244 152658
rect 22192 152594 22244 152600
rect 19340 152584 19392 152590
rect 12438 152552 12494 152561
rect 19340 152526 19392 152532
rect 12438 152487 12494 152496
rect 8850 152416 8906 152425
rect 8850 152351 8906 152360
rect 19800 152244 19852 152250
rect 19800 152186 19852 152192
rect 9496 152176 9548 152182
rect 9496 152118 9548 152124
rect 6090 150648 6146 150657
rect 6090 150583 6146 150592
rect 2686 150512 2742 150521
rect 2686 150447 2742 150456
rect 2700 149940 2728 150447
rect 6104 149940 6132 150583
rect 9508 149940 9536 152118
rect 16396 151428 16448 151434
rect 16396 151370 16448 151376
rect 12992 151360 13044 151366
rect 12992 151302 13044 151308
rect 13004 149940 13032 151302
rect 16408 149940 16436 151370
rect 19812 149940 19840 152186
rect 23308 149940 23336 153138
rect 26436 152794 26464 163200
rect 27264 154222 27292 163200
rect 28092 156641 28120 163200
rect 28078 156632 28134 156641
rect 28078 156567 28134 156576
rect 27252 154216 27304 154222
rect 27252 154158 27304 154164
rect 26424 152788 26476 152794
rect 26424 152730 26476 152736
rect 28184 152726 28212 163254
rect 28828 163146 28856 163254
rect 28906 163200 28962 164400
rect 29826 163200 29882 164400
rect 30392 163254 30604 163282
rect 28920 163146 28948 163200
rect 28828 163118 28948 163146
rect 29840 159633 29868 163200
rect 29826 159624 29882 159633
rect 29826 159559 29882 159568
rect 30392 154193 30420 163254
rect 30576 163146 30604 163254
rect 30654 163200 30710 164400
rect 31482 163200 31538 164400
rect 32310 163200 32366 164400
rect 33138 163200 33194 164400
rect 33966 163200 34022 164400
rect 34532 163254 34744 163282
rect 30668 163146 30696 163200
rect 30576 163118 30696 163146
rect 31496 156777 31524 163200
rect 32324 159526 32352 163200
rect 32312 159520 32364 159526
rect 32312 159462 32364 159468
rect 31482 156768 31538 156777
rect 31482 156703 31538 156712
rect 30378 154184 30434 154193
rect 30378 154119 30434 154128
rect 33152 152862 33180 163200
rect 33980 158001 34008 163200
rect 33966 157992 34022 158001
rect 33966 157927 34022 157936
rect 34532 154358 34560 163254
rect 34716 163146 34744 163254
rect 34794 163200 34850 164400
rect 35714 163200 35770 164400
rect 36542 163200 36598 164400
rect 37370 163200 37426 164400
rect 37936 163254 38148 163282
rect 34808 163146 34836 163200
rect 34716 163118 34836 163146
rect 35728 157078 35756 163200
rect 36556 159458 36584 163200
rect 36544 159452 36596 159458
rect 36544 159394 36596 159400
rect 37384 158098 37412 163200
rect 37372 158092 37424 158098
rect 37372 158034 37424 158040
rect 35716 157072 35768 157078
rect 35716 157014 35768 157020
rect 34520 154352 34572 154358
rect 34520 154294 34572 154300
rect 37936 154290 37964 163254
rect 38120 163146 38148 163254
rect 38198 163200 38254 164400
rect 39026 163200 39082 164400
rect 39854 163200 39910 164400
rect 40682 163200 40738 164400
rect 41602 163200 41658 164400
rect 42430 163200 42486 164400
rect 43258 163200 43314 164400
rect 44086 163200 44142 164400
rect 44192 163254 44864 163282
rect 38212 163146 38240 163200
rect 38120 163118 38240 163146
rect 39040 157146 39068 163200
rect 39028 157140 39080 157146
rect 39028 157082 39080 157088
rect 39868 155582 39896 163200
rect 40696 158273 40724 163200
rect 40682 158264 40738 158273
rect 40682 158199 40738 158208
rect 39856 155576 39908 155582
rect 39856 155518 39908 155524
rect 37924 154284 37976 154290
rect 37924 154226 37976 154232
rect 41616 153270 41644 163200
rect 42444 157214 42472 163200
rect 43272 159594 43300 163200
rect 43260 159588 43312 159594
rect 43260 159530 43312 159536
rect 44100 158137 44128 163200
rect 44086 158128 44142 158137
rect 44086 158063 44142 158072
rect 42432 157208 42484 157214
rect 42432 157150 42484 157156
rect 44192 154494 44220 163254
rect 44836 163146 44864 163254
rect 44914 163200 44970 164400
rect 45742 163200 45798 164400
rect 46570 163200 46626 164400
rect 47490 163200 47546 164400
rect 48318 163200 48374 164400
rect 49146 163200 49202 164400
rect 49974 163200 50030 164400
rect 50802 163200 50858 164400
rect 51092 163254 51580 163282
rect 44928 163146 44956 163200
rect 44836 163118 44956 163146
rect 45756 157282 45784 163200
rect 45744 157276 45796 157282
rect 45744 157218 45796 157224
rect 46584 155718 46612 163200
rect 47504 158234 47532 163200
rect 47492 158228 47544 158234
rect 47492 158170 47544 158176
rect 46572 155712 46624 155718
rect 46572 155654 46624 155660
rect 44180 154488 44232 154494
rect 44180 154430 44232 154436
rect 48332 153814 48360 163200
rect 49160 157350 49188 163200
rect 49988 159662 50016 163200
rect 49976 159656 50028 159662
rect 49976 159598 50028 159604
rect 50816 158166 50844 163200
rect 50804 158160 50856 158166
rect 50804 158102 50856 158108
rect 49148 157344 49200 157350
rect 49148 157286 49200 157292
rect 51092 154562 51120 163254
rect 51552 163146 51580 163254
rect 51630 163200 51686 164400
rect 52458 163200 52514 164400
rect 53378 163200 53434 164400
rect 54206 163200 54262 164400
rect 54312 163254 54984 163282
rect 51644 163146 51672 163200
rect 51552 163118 51672 163146
rect 52472 156602 52500 163200
rect 52460 156596 52512 156602
rect 52460 156538 52512 156544
rect 53392 155650 53420 163200
rect 54220 158302 54248 163200
rect 54208 158296 54260 158302
rect 54208 158238 54260 158244
rect 53380 155644 53432 155650
rect 53380 155586 53432 155592
rect 51080 154556 51132 154562
rect 51080 154498 51132 154504
rect 54312 154329 54340 163254
rect 54956 163146 54984 163254
rect 55034 163200 55090 164400
rect 55862 163200 55918 164400
rect 56690 163200 56746 164400
rect 57518 163200 57574 164400
rect 57992 163254 58296 163282
rect 55048 163146 55076 163200
rect 54956 163118 55076 163146
rect 55876 156913 55904 163200
rect 56704 159866 56732 163200
rect 56692 159860 56744 159866
rect 56692 159802 56744 159808
rect 57532 158409 57560 163200
rect 57518 158400 57574 158409
rect 57518 158335 57574 158344
rect 55862 156904 55918 156913
rect 55862 156839 55918 156848
rect 54298 154320 54354 154329
rect 54298 154255 54354 154264
rect 48320 153808 48372 153814
rect 48320 153750 48372 153756
rect 57992 153678 58020 163254
rect 58268 163146 58296 163254
rect 58346 163200 58402 164400
rect 59266 163200 59322 164400
rect 60094 163200 60150 164400
rect 60922 163200 60978 164400
rect 61120 163254 61700 163282
rect 58360 163146 58388 163200
rect 58268 163118 58388 163146
rect 59280 156534 59308 163200
rect 59268 156528 59320 156534
rect 59268 156470 59320 156476
rect 60108 155854 60136 163200
rect 60936 158438 60964 163200
rect 60924 158432 60976 158438
rect 60924 158374 60976 158380
rect 60096 155848 60148 155854
rect 60096 155790 60148 155796
rect 61120 153746 61148 163254
rect 61672 163146 61700 163254
rect 61750 163200 61806 164400
rect 62578 163200 62634 164400
rect 63406 163200 63462 164400
rect 64234 163200 64290 164400
rect 65154 163200 65210 164400
rect 65982 163200 66038 164400
rect 66810 163200 66866 164400
rect 67638 163200 67694 164400
rect 68466 163200 68522 164400
rect 69294 163200 69350 164400
rect 70122 163200 70178 164400
rect 71042 163200 71098 164400
rect 71870 163200 71926 164400
rect 72698 163200 72754 164400
rect 73526 163200 73582 164400
rect 74354 163200 74410 164400
rect 75182 163200 75238 164400
rect 76010 163200 76066 164400
rect 76930 163200 76986 164400
rect 77758 163200 77814 164400
rect 78586 163200 78642 164400
rect 78692 163254 79364 163282
rect 61764 163146 61792 163200
rect 61672 163118 61792 163146
rect 62592 155553 62620 163200
rect 63420 160070 63448 163200
rect 63408 160064 63460 160070
rect 63408 160006 63460 160012
rect 64248 158370 64276 163200
rect 64236 158364 64288 158370
rect 64236 158306 64288 158312
rect 62578 155544 62634 155553
rect 65168 155514 65196 163200
rect 62578 155479 62634 155488
rect 65156 155508 65208 155514
rect 65156 155450 65208 155456
rect 65996 155281 66024 163200
rect 66824 155922 66852 163200
rect 67652 158642 67680 163200
rect 67640 158636 67692 158642
rect 67640 158578 67692 158584
rect 66812 155916 66864 155922
rect 66812 155858 66864 155864
rect 66628 155644 66680 155650
rect 66628 155586 66680 155592
rect 65982 155272 66038 155281
rect 65982 155207 66038 155216
rect 61108 153740 61160 153746
rect 61108 153682 61160 153688
rect 57980 153672 58032 153678
rect 57980 153614 58032 153620
rect 41604 153264 41656 153270
rect 41604 153206 41656 153212
rect 33140 152856 33192 152862
rect 33140 152798 33192 152804
rect 28172 152720 28224 152726
rect 28172 152662 28224 152668
rect 66640 152454 66668 155586
rect 68480 155417 68508 163200
rect 69308 156466 69336 163200
rect 70136 159798 70164 163200
rect 70124 159792 70176 159798
rect 70124 159734 70176 159740
rect 71056 158506 71084 163200
rect 71044 158500 71096 158506
rect 71044 158442 71096 158448
rect 69296 156460 69348 156466
rect 69296 156402 69348 156408
rect 71884 155650 71912 163200
rect 72712 157049 72740 163200
rect 73540 159322 73568 163200
rect 73528 159316 73580 159322
rect 73528 159258 73580 159264
rect 74368 158574 74396 163200
rect 74356 158568 74408 158574
rect 74356 158510 74408 158516
rect 72698 157040 72754 157049
rect 72698 156975 72754 156984
rect 75092 155712 75144 155718
rect 75092 155654 75144 155660
rect 71872 155644 71924 155650
rect 71872 155586 71924 155592
rect 68928 155576 68980 155582
rect 68928 155518 68980 155524
rect 68466 155408 68522 155417
rect 68466 155343 68522 155352
rect 66628 152448 66680 152454
rect 66628 152390 66680 152396
rect 33600 152380 33652 152386
rect 33600 152322 33652 152328
rect 30196 151904 30248 151910
rect 30196 151846 30248 151852
rect 26700 151496 26752 151502
rect 26700 151438 26752 151444
rect 26712 149940 26740 151438
rect 30208 149940 30236 151846
rect 33612 149940 33640 152322
rect 68940 152046 68968 155518
rect 71412 152924 71464 152930
rect 71412 152866 71464 152872
rect 68928 152040 68980 152046
rect 68928 151982 68980 151988
rect 43904 151700 43956 151706
rect 43904 151642 43956 151648
rect 40500 151632 40552 151638
rect 40500 151574 40552 151580
rect 37004 151564 37056 151570
rect 37004 151506 37056 151512
rect 37016 149940 37044 151506
rect 40512 149940 40540 151574
rect 43916 149940 43944 151642
rect 68008 151292 68060 151298
rect 68008 151234 68060 151240
rect 64512 151224 64564 151230
rect 64512 151166 64564 151172
rect 61108 151156 61160 151162
rect 61108 151098 61160 151104
rect 57704 151088 57756 151094
rect 57704 151030 57756 151036
rect 54208 151020 54260 151026
rect 54208 150962 54260 150968
rect 50804 150952 50856 150958
rect 50804 150894 50856 150900
rect 47308 150884 47360 150890
rect 47308 150826 47360 150832
rect 47320 149940 47348 150826
rect 50816 149940 50844 150894
rect 54220 149940 54248 150962
rect 57716 149940 57744 151030
rect 61120 149940 61148 151098
rect 64524 149940 64552 151166
rect 68020 149940 68048 151234
rect 71424 149940 71452 152866
rect 75104 151978 75132 155654
rect 75196 155582 75224 163200
rect 76024 155825 76052 163200
rect 76944 159934 76972 163200
rect 76932 159928 76984 159934
rect 76932 159870 76984 159876
rect 77772 157962 77800 163200
rect 77760 157956 77812 157962
rect 77760 157898 77812 157904
rect 76010 155816 76066 155825
rect 76010 155751 76066 155760
rect 78600 155689 78628 163200
rect 78586 155680 78642 155689
rect 78586 155615 78642 155624
rect 75184 155576 75236 155582
rect 75184 155518 75236 155524
rect 78692 153610 78720 163254
rect 79336 163146 79364 163254
rect 79414 163200 79470 164400
rect 80242 163200 80298 164400
rect 81070 163200 81126 164400
rect 81898 163200 81954 164400
rect 82818 163200 82874 164400
rect 83646 163200 83702 164400
rect 84474 163200 84530 164400
rect 85302 163200 85358 164400
rect 85592 163254 86080 163282
rect 79428 163146 79456 163200
rect 79336 163118 79456 163146
rect 80060 159316 80112 159322
rect 80060 159258 80112 159264
rect 79324 155848 79376 155854
rect 79324 155790 79376 155796
rect 78680 153604 78732 153610
rect 78680 153546 78732 153552
rect 79336 152114 79364 155790
rect 80072 153134 80100 159258
rect 80256 159254 80284 163200
rect 80244 159248 80296 159254
rect 80244 159190 80296 159196
rect 81084 158710 81112 163200
rect 81072 158704 81124 158710
rect 81072 158646 81124 158652
rect 81912 155718 81940 163200
rect 82832 156398 82860 163200
rect 83660 159322 83688 163200
rect 83648 159316 83700 159322
rect 83648 159258 83700 159264
rect 84488 157894 84516 163200
rect 84476 157888 84528 157894
rect 84476 157830 84528 157836
rect 82820 156392 82872 156398
rect 82820 156334 82872 156340
rect 85316 155961 85344 163200
rect 85302 155952 85358 155961
rect 82912 155916 82964 155922
rect 85302 155887 85358 155896
rect 82912 155858 82964 155864
rect 81900 155712 81952 155718
rect 81900 155654 81952 155660
rect 80060 153128 80112 153134
rect 80060 153070 80112 153076
rect 82924 152182 82952 155858
rect 85592 154465 85620 163254
rect 86052 163146 86080 163254
rect 86130 163200 86186 164400
rect 86958 163200 87014 164400
rect 87786 163200 87842 164400
rect 88706 163200 88762 164400
rect 89534 163200 89590 164400
rect 90362 163200 90418 164400
rect 91190 163200 91246 164400
rect 92018 163200 92074 164400
rect 92846 163200 92902 164400
rect 93674 163200 93730 164400
rect 94594 163200 94650 164400
rect 95422 163200 95478 164400
rect 96250 163200 96306 164400
rect 96632 163254 97028 163282
rect 86144 163146 86172 163200
rect 86052 163118 86172 163146
rect 86972 159186 87000 163200
rect 86960 159180 87012 159186
rect 86960 159122 87012 159128
rect 87800 157826 87828 163200
rect 87788 157820 87840 157826
rect 87788 157762 87840 157768
rect 88720 155922 88748 163200
rect 88708 155916 88760 155922
rect 88708 155858 88760 155864
rect 89548 155174 89576 163200
rect 90376 158778 90404 163200
rect 91100 159248 91152 159254
rect 91100 159190 91152 159196
rect 90364 158772 90416 158778
rect 90364 158714 90416 158720
rect 89536 155168 89588 155174
rect 89536 155110 89588 155116
rect 85578 154456 85634 154465
rect 85578 154391 85634 154400
rect 91112 152318 91140 159190
rect 91204 157758 91232 163200
rect 91192 157752 91244 157758
rect 91192 157694 91244 157700
rect 92032 155854 92060 163200
rect 92860 158778 92888 163200
rect 93688 159118 93716 163200
rect 93676 159112 93728 159118
rect 93676 159054 93728 159060
rect 92572 158772 92624 158778
rect 92572 158714 92624 158720
rect 92848 158772 92900 158778
rect 92848 158714 92900 158720
rect 92020 155848 92072 155854
rect 92020 155790 92072 155796
rect 92584 152998 92612 158714
rect 94608 157690 94636 163200
rect 94596 157684 94648 157690
rect 94596 157626 94648 157632
rect 95436 155038 95464 163200
rect 96264 158982 96292 163200
rect 96252 158976 96304 158982
rect 96252 158918 96304 158924
rect 95424 155032 95476 155038
rect 95424 154974 95476 154980
rect 92572 152992 92624 152998
rect 92572 152934 92624 152940
rect 96632 152930 96660 163254
rect 97000 163146 97028 163254
rect 97078 163200 97134 164400
rect 97906 163200 97962 164400
rect 98734 163200 98790 164400
rect 99562 163200 99618 164400
rect 100482 163200 100538 164400
rect 101310 163200 101366 164400
rect 102138 163200 102194 164400
rect 102966 163200 103022 164400
rect 103532 163254 103744 163282
rect 97092 163146 97120 163200
rect 97000 163118 97120 163146
rect 97920 157622 97948 163200
rect 97908 157616 97960 157622
rect 97908 157558 97960 157564
rect 98748 155106 98776 163200
rect 99576 156330 99604 163200
rect 100496 159254 100524 163200
rect 100484 159248 100536 159254
rect 100484 159190 100536 159196
rect 99564 156324 99616 156330
rect 99564 156266 99616 156272
rect 101324 156262 101352 163200
rect 101312 156256 101364 156262
rect 101312 156198 101364 156204
rect 98736 155100 98788 155106
rect 98736 155042 98788 155048
rect 102152 153542 102180 163200
rect 102980 158914 103008 163200
rect 102968 158908 103020 158914
rect 102968 158850 103020 158856
rect 102140 153536 102192 153542
rect 102140 153478 102192 153484
rect 103532 153066 103560 163254
rect 103716 163146 103744 163254
rect 103794 163200 103850 164400
rect 104622 163200 104678 164400
rect 104912 163254 105400 163282
rect 103808 163146 103836 163200
rect 103716 163118 103836 163146
rect 104636 158545 104664 163200
rect 104622 158536 104678 158545
rect 104622 158471 104678 158480
rect 104912 153474 104940 163254
rect 105372 163146 105400 163254
rect 105450 163200 105506 164400
rect 106370 163200 106426 164400
rect 107198 163200 107254 164400
rect 108026 163200 108082 164400
rect 108316 163254 108804 163282
rect 105464 163146 105492 163200
rect 105372 163118 105492 163146
rect 106384 154902 106412 163200
rect 107212 159050 107240 163200
rect 107200 159044 107252 159050
rect 107200 158986 107252 158992
rect 108040 156194 108068 163200
rect 108028 156188 108080 156194
rect 108028 156130 108080 156136
rect 106372 154896 106424 154902
rect 106372 154838 106424 154844
rect 104900 153468 104952 153474
rect 104900 153410 104952 153416
rect 108316 153406 108344 163254
rect 108776 163146 108804 163254
rect 108854 163200 108910 164400
rect 109682 163200 109738 164400
rect 110510 163200 110566 164400
rect 111338 163200 111394 164400
rect 112258 163200 112314 164400
rect 113086 163200 113142 164400
rect 113192 163254 113864 163282
rect 108868 163146 108896 163200
rect 108776 163118 108896 163146
rect 109132 159724 109184 159730
rect 109132 159666 109184 159672
rect 109040 154964 109092 154970
rect 109040 154906 109092 154912
rect 108304 153400 108356 153406
rect 108304 153342 108356 153348
rect 103520 153060 103572 153066
rect 103520 153002 103572 153008
rect 92480 152924 92532 152930
rect 92480 152866 92532 152872
rect 96620 152924 96672 152930
rect 96620 152866 96672 152872
rect 91100 152312 91152 152318
rect 91100 152254 91152 152260
rect 82820 152176 82872 152182
rect 82820 152118 82872 152124
rect 82912 152176 82964 152182
rect 82912 152118 82964 152124
rect 79324 152108 79376 152114
rect 79324 152050 79376 152056
rect 75092 151972 75144 151978
rect 75092 151914 75144 151920
rect 74816 151836 74868 151842
rect 81348 151836 81400 151842
rect 74868 151786 74948 151814
rect 74816 151778 74868 151784
rect 74920 149954 74948 151786
rect 81348 151778 81400 151784
rect 78312 150340 78364 150346
rect 78312 150282 78364 150288
rect 74842 149926 74948 149954
rect 78324 149940 78352 150282
rect 81360 150142 81388 151778
rect 81716 151768 81768 151774
rect 81716 151710 81768 151716
rect 81348 150136 81400 150142
rect 81348 150078 81400 150084
rect 81728 149940 81756 151710
rect 82832 149705 82860 152118
rect 92020 150680 92072 150686
rect 92020 150622 92072 150628
rect 88616 150612 88668 150618
rect 88616 150554 88668 150560
rect 85212 150544 85264 150550
rect 85212 150486 85264 150492
rect 85224 149940 85252 150486
rect 88628 149940 88656 150554
rect 92032 149940 92060 150622
rect 92492 150142 92520 152866
rect 109052 152250 109080 154906
rect 109144 154698 109172 159666
rect 109696 158846 109724 163200
rect 109776 159996 109828 160002
rect 109776 159938 109828 159944
rect 109684 158840 109736 158846
rect 109684 158782 109736 158788
rect 109132 154692 109184 154698
rect 109132 154634 109184 154640
rect 109788 152386 109816 159938
rect 110328 155780 110380 155786
rect 110328 155722 110380 155728
rect 109684 152380 109736 152386
rect 109684 152322 109736 152328
rect 109776 152380 109828 152386
rect 109776 152322 109828 152328
rect 97908 152244 97960 152250
rect 97908 152186 97960 152192
rect 109040 152244 109092 152250
rect 109040 152186 109092 152192
rect 95516 150748 95568 150754
rect 95516 150690 95568 150696
rect 92480 150136 92532 150142
rect 92480 150078 92532 150084
rect 95528 149940 95556 150690
rect 97920 150210 97948 152186
rect 105820 151836 105872 151842
rect 105740 151786 105820 151814
rect 98920 150816 98972 150822
rect 98920 150758 98972 150764
rect 97908 150204 97960 150210
rect 97908 150146 97960 150152
rect 98932 149940 98960 150758
rect 102324 150476 102376 150482
rect 102324 150418 102376 150424
rect 102336 149940 102364 150418
rect 105740 149954 105768 151786
rect 105820 151778 105872 151784
rect 105740 149926 105846 149954
rect 82818 149696 82874 149705
rect 82818 149631 82874 149640
rect 109250 149382 109632 149410
rect 109604 148073 109632 149382
rect 109590 148064 109646 148073
rect 109590 147999 109646 148008
rect 109696 132494 109724 152322
rect 110340 151994 110368 155722
rect 110524 154766 110552 163200
rect 111352 157554 111380 163200
rect 111340 157548 111392 157554
rect 111340 157490 111392 157496
rect 112272 155786 112300 163200
rect 113100 159730 113128 163200
rect 113088 159724 113140 159730
rect 113088 159666 113140 159672
rect 112260 155780 112312 155786
rect 112260 155722 112312 155728
rect 110512 154760 110564 154766
rect 110512 154702 110564 154708
rect 113192 153202 113220 163254
rect 113836 163146 113864 163254
rect 113914 163200 113970 164400
rect 114742 163200 114798 164400
rect 115570 163200 115626 164400
rect 115952 163254 116348 163282
rect 113928 163146 113956 163200
rect 113836 163118 113956 163146
rect 114468 158772 114520 158778
rect 114468 158714 114520 158720
rect 114480 154426 114508 158714
rect 114756 157486 114784 163200
rect 114744 157480 114796 157486
rect 114744 157422 114796 157428
rect 115584 157185 115612 163200
rect 115570 157176 115626 157185
rect 115570 157111 115626 157120
rect 114468 154420 114520 154426
rect 114468 154362 114520 154368
rect 115952 153338 115980 163254
rect 116320 163146 116348 163254
rect 116398 163200 116454 164400
rect 117226 163200 117282 164400
rect 118146 163200 118202 164400
rect 118712 163254 118924 163282
rect 116412 163146 116440 163200
rect 116320 163118 116440 163146
rect 117240 160002 117268 163200
rect 117228 159996 117280 160002
rect 117228 159938 117280 159944
rect 118160 156126 118188 163200
rect 118148 156120 118200 156126
rect 118148 156062 118200 156068
rect 118608 154624 118660 154630
rect 118608 154566 118660 154572
rect 118620 154426 118648 154566
rect 118712 154426 118740 163254
rect 118896 163146 118924 163254
rect 118974 163200 119030 164400
rect 119802 163200 119858 164400
rect 120092 163254 120580 163282
rect 118988 163146 119016 163200
rect 118896 163118 119016 163146
rect 119816 158778 119844 163200
rect 119804 158772 119856 158778
rect 119804 158714 119856 158720
rect 118884 158024 118936 158030
rect 118884 157966 118936 157972
rect 118608 154420 118660 154426
rect 118608 154362 118660 154368
rect 118700 154420 118752 154426
rect 118700 154362 118752 154368
rect 115940 153332 115992 153338
rect 115940 153274 115992 153280
rect 110972 153196 111024 153202
rect 110972 153138 111024 153144
rect 113180 153196 113232 153202
rect 113180 153138 113232 153144
rect 110512 152380 110564 152386
rect 110512 152322 110564 152328
rect 110340 151966 110460 151994
rect 110328 151904 110380 151910
rect 110328 151846 110380 151852
rect 110236 151836 110288 151842
rect 110236 151778 110288 151784
rect 110248 146418 110276 151778
rect 110340 150278 110368 151846
rect 110432 151842 110460 151966
rect 110524 151910 110552 152322
rect 110512 151904 110564 151910
rect 110512 151846 110564 151852
rect 110420 151836 110472 151842
rect 110984 151814 111012 153138
rect 110984 151786 111196 151814
rect 110420 151778 110472 151784
rect 111064 151564 111116 151570
rect 111064 151506 111116 151512
rect 110878 150512 110934 150521
rect 110878 150447 110934 150456
rect 110328 150272 110380 150278
rect 110328 150214 110380 150220
rect 110892 148050 110920 150447
rect 111076 148322 111104 151506
rect 111168 148442 111196 151786
rect 112812 151768 112864 151774
rect 112812 151710 112864 151716
rect 111432 151700 111484 151706
rect 111432 151642 111484 151648
rect 111340 151632 111392 151638
rect 111340 151574 111392 151580
rect 111246 150648 111302 150657
rect 111246 150583 111302 150592
rect 111156 148436 111208 148442
rect 111156 148378 111208 148384
rect 111076 148294 111196 148322
rect 110892 148022 111104 148050
rect 110326 146432 110382 146441
rect 110248 146390 110326 146418
rect 110326 146367 110382 146376
rect 109696 132466 110368 132494
rect 110340 106321 110368 132466
rect 110326 106312 110382 106321
rect 110326 106247 110382 106256
rect 111076 89690 111104 148022
rect 111168 109002 111196 148294
rect 111156 108996 111208 109002
rect 111156 108938 111208 108944
rect 111260 92478 111288 150583
rect 111352 111790 111380 151574
rect 111444 113150 111472 151642
rect 112720 151292 112772 151298
rect 112720 151234 112772 151240
rect 112628 151224 112680 151230
rect 112628 151166 112680 151172
rect 112536 151156 112588 151162
rect 112536 151098 112588 151104
rect 111708 151088 111760 151094
rect 111708 151030 111760 151036
rect 111616 150952 111668 150958
rect 111616 150894 111668 150900
rect 111524 150884 111576 150890
rect 111524 150826 111576 150832
rect 111536 114510 111564 150826
rect 111628 117298 111656 150894
rect 111720 121446 111748 151030
rect 112444 151020 112496 151026
rect 112444 150962 112496 150968
rect 111708 121440 111760 121446
rect 111708 121382 111760 121388
rect 112456 118658 112484 150962
rect 112548 122806 112576 151098
rect 112640 124166 112668 151166
rect 112732 126954 112760 151234
rect 112824 133890 112852 151710
rect 116952 151496 117004 151502
rect 116952 151438 117004 151444
rect 116768 151428 116820 151434
rect 116768 151370 116820 151376
rect 116676 151360 116728 151366
rect 116676 151302 116728 151308
rect 116032 150816 116084 150822
rect 116032 150758 116084 150764
rect 115296 150748 115348 150754
rect 115296 150690 115348 150696
rect 113088 150680 113140 150686
rect 113088 150622 113140 150628
rect 112996 150612 113048 150618
rect 112996 150554 113048 150560
rect 112904 150340 112956 150346
rect 112904 150282 112956 150288
rect 112812 133884 112864 133890
rect 112812 133826 112864 133832
rect 112916 132462 112944 150282
rect 113008 137970 113036 150554
rect 113100 140758 113128 150622
rect 115204 150544 115256 150550
rect 115204 150486 115256 150492
rect 113822 144256 113878 144265
rect 113822 144191 113878 144200
rect 113088 140752 113140 140758
rect 113088 140694 113140 140700
rect 112996 137964 113048 137970
rect 112996 137906 113048 137912
rect 112904 132456 112956 132462
rect 112904 132398 112956 132404
rect 112720 126948 112772 126954
rect 112720 126890 112772 126896
rect 112628 124160 112680 124166
rect 112628 124102 112680 124108
rect 112536 122800 112588 122806
rect 112536 122742 112588 122748
rect 112444 118652 112496 118658
rect 112444 118594 112496 118600
rect 111616 117292 111668 117298
rect 111616 117234 111668 117240
rect 111524 114504 111576 114510
rect 111524 114446 111576 114452
rect 111432 113144 111484 113150
rect 111432 113086 111484 113092
rect 111340 111784 111392 111790
rect 111340 111726 111392 111732
rect 111248 92472 111300 92478
rect 111248 92414 111300 92420
rect 111064 89684 111116 89690
rect 111064 89626 111116 89632
rect 113836 88330 113864 144191
rect 115216 135561 115244 150486
rect 115308 141409 115336 150690
rect 116044 143313 116072 150758
rect 116124 150476 116176 150482
rect 116124 150418 116176 150424
rect 116136 145217 116164 150418
rect 116492 150068 116544 150074
rect 116492 150010 116544 150016
rect 116122 145208 116178 145217
rect 116122 145143 116178 145152
rect 116030 143304 116086 143313
rect 116030 143239 116086 143248
rect 115294 141400 115350 141409
rect 115294 141335 115350 141344
rect 116124 140752 116176 140758
rect 116124 140694 116176 140700
rect 116136 139505 116164 140694
rect 116122 139496 116178 139505
rect 116122 139431 116178 139440
rect 116124 137964 116176 137970
rect 116124 137906 116176 137912
rect 116136 137601 116164 137906
rect 116122 137592 116178 137601
rect 116122 137527 116178 137536
rect 115202 135552 115258 135561
rect 115202 135487 115258 135496
rect 116032 133884 116084 133890
rect 116032 133826 116084 133832
rect 116044 133657 116072 133826
rect 116030 133648 116086 133657
rect 116030 133583 116086 133592
rect 114190 132832 114246 132841
rect 114190 132767 114246 132776
rect 114204 132666 114232 132767
rect 114192 132660 114244 132666
rect 114192 132602 114244 132608
rect 115204 132660 115256 132666
rect 115204 132602 115256 132608
rect 113914 121408 113970 121417
rect 113914 121343 113970 121352
rect 113824 88324 113876 88330
rect 113824 88266 113876 88272
rect 113928 83978 113956 121343
rect 114006 110120 114062 110129
rect 114006 110055 114062 110064
rect 113916 83972 113968 83978
rect 113916 83914 113968 83920
rect 114020 82822 114048 110055
rect 114098 98696 114154 98705
rect 114098 98631 114154 98640
rect 114008 82816 114060 82822
rect 114008 82758 114060 82764
rect 114112 80034 114140 98631
rect 114190 87272 114246 87281
rect 114190 87207 114246 87216
rect 114100 80028 114152 80034
rect 114100 79970 114152 79976
rect 114204 78674 114232 87207
rect 115216 85649 115244 132602
rect 116124 132456 116176 132462
rect 116124 132398 116176 132404
rect 116136 131753 116164 132398
rect 116122 131744 116178 131753
rect 116122 131679 116178 131688
rect 116504 129849 116532 150010
rect 116582 149696 116638 149705
rect 116582 149631 116638 149640
rect 116490 129840 116546 129849
rect 116490 129775 116546 129784
rect 116124 126948 116176 126954
rect 116124 126890 116176 126896
rect 116136 126041 116164 126890
rect 116122 126032 116178 126041
rect 116122 125967 116178 125976
rect 116124 124160 116176 124166
rect 116122 124128 116124 124137
rect 116176 124128 116178 124137
rect 116122 124063 116178 124072
rect 115940 122800 115992 122806
rect 115940 122742 115992 122748
rect 115952 122233 115980 122742
rect 115938 122224 115994 122233
rect 115938 122159 115994 122168
rect 116124 121440 116176 121446
rect 116124 121382 116176 121388
rect 116136 120193 116164 121382
rect 116122 120184 116178 120193
rect 116122 120119 116178 120128
rect 116124 118652 116176 118658
rect 116124 118594 116176 118600
rect 116136 118289 116164 118594
rect 116122 118280 116178 118289
rect 116122 118215 116178 118224
rect 116124 117292 116176 117298
rect 116124 117234 116176 117240
rect 116136 116385 116164 117234
rect 116122 116376 116178 116385
rect 116122 116311 116178 116320
rect 116124 114504 116176 114510
rect 116122 114472 116124 114481
rect 116176 114472 116178 114481
rect 116122 114407 116178 114416
rect 115940 113144 115992 113150
rect 115940 113086 115992 113092
rect 115952 112577 115980 113086
rect 115938 112568 115994 112577
rect 115938 112503 115994 112512
rect 116124 111784 116176 111790
rect 116124 111726 116176 111732
rect 116136 110673 116164 111726
rect 116122 110664 116178 110673
rect 116122 110599 116178 110608
rect 116124 108996 116176 109002
rect 116124 108938 116176 108944
rect 116136 108769 116164 108938
rect 116122 108760 116178 108769
rect 116122 108695 116178 108704
rect 116596 93401 116624 149631
rect 116688 95305 116716 151302
rect 116780 97209 116808 151370
rect 116860 150204 116912 150210
rect 116860 150146 116912 150152
rect 116872 99113 116900 150146
rect 116964 102921 116992 151438
rect 117136 150272 117188 150278
rect 117136 150214 117188 150220
rect 117044 148368 117096 148374
rect 117044 148310 117096 148316
rect 116950 102912 117006 102921
rect 116950 102847 117006 102856
rect 117056 101017 117084 148310
rect 117148 104825 117176 150214
rect 117228 150136 117280 150142
rect 117228 150078 117280 150084
rect 117240 132546 117268 150078
rect 118896 149954 118924 157966
rect 119988 154624 120040 154630
rect 119988 154566 120040 154572
rect 120000 154426 120028 154566
rect 119896 154420 119948 154426
rect 119896 154362 119948 154368
rect 119988 154420 120040 154426
rect 119988 154362 120040 154368
rect 119908 153882 119936 154362
rect 119804 153876 119856 153882
rect 119804 153818 119856 153824
rect 119896 153876 119948 153882
rect 119896 153818 119948 153824
rect 119816 150226 119844 153818
rect 120092 152386 120120 163254
rect 120552 163146 120580 163254
rect 120630 163200 120686 164400
rect 121458 163200 121514 164400
rect 122286 163200 122342 164400
rect 123114 163200 123170 164400
rect 124034 163200 124090 164400
rect 124862 163200 124918 164400
rect 125690 163200 125746 164400
rect 126518 163200 126574 164400
rect 126992 163254 127296 163282
rect 120644 163146 120672 163200
rect 120552 163118 120672 163146
rect 120448 156664 120500 156670
rect 120448 156606 120500 156612
rect 120080 152380 120132 152386
rect 120080 152322 120132 152328
rect 120460 150226 120488 156606
rect 121472 156058 121500 163200
rect 121920 158976 121972 158982
rect 121920 158918 121972 158924
rect 121460 156052 121512 156058
rect 121460 155994 121512 156000
rect 121932 153785 121960 158918
rect 122012 155304 122064 155310
rect 122012 155246 122064 155252
rect 121734 153776 121790 153785
rect 121734 153711 121790 153720
rect 121918 153776 121974 153785
rect 121918 153711 121974 153720
rect 121092 152516 121144 152522
rect 121092 152458 121144 152464
rect 121104 150226 121132 152458
rect 121748 150226 121776 153711
rect 122024 151814 122052 155246
rect 122300 154970 122328 163200
rect 123128 159390 123156 163200
rect 122840 159384 122892 159390
rect 122840 159326 122892 159332
rect 123116 159384 123168 159390
rect 123116 159326 123168 159332
rect 122288 154964 122340 154970
rect 122288 154906 122340 154912
rect 122024 151786 122420 151814
rect 122392 150226 122420 151786
rect 119816 150198 119890 150226
rect 120460 150198 120534 150226
rect 121104 150198 121178 150226
rect 121748 150198 121822 150226
rect 122392 150198 122466 150226
rect 122852 150210 122880 159326
rect 124048 158982 124076 163200
rect 124036 158976 124088 158982
rect 124036 158918 124088 158924
rect 124876 156670 124904 163200
rect 125704 161474 125732 163200
rect 125704 161446 125824 161474
rect 125508 158908 125560 158914
rect 125508 158850 125560 158856
rect 124864 156664 124916 156670
rect 124864 156606 124916 156612
rect 124680 155440 124732 155446
rect 124680 155382 124732 155388
rect 123024 155236 123076 155242
rect 123024 155178 123076 155184
rect 123036 150226 123064 155178
rect 124312 153944 124364 153950
rect 124312 153886 124364 153892
rect 124324 150226 124352 153886
rect 124692 151814 124720 155382
rect 125520 153950 125548 158850
rect 125692 155372 125744 155378
rect 125692 155314 125744 155320
rect 125508 153944 125560 153950
rect 125508 153886 125560 153892
rect 124692 151786 124996 151814
rect 124968 150226 124996 151786
rect 125704 150226 125732 155314
rect 125796 154834 125824 161446
rect 126532 159730 126560 163200
rect 126428 159724 126480 159730
rect 126428 159666 126480 159672
rect 126520 159724 126572 159730
rect 126520 159666 126572 159672
rect 126440 159526 126468 159666
rect 126428 159520 126480 159526
rect 126428 159462 126480 159468
rect 126244 159452 126296 159458
rect 126244 159394 126296 159400
rect 126796 159452 126848 159458
rect 126796 159394 126848 159400
rect 126256 158914 126284 159394
rect 126244 158908 126296 158914
rect 126244 158850 126296 158856
rect 125784 154828 125836 154834
rect 125784 154770 125836 154776
rect 126808 152425 126836 159394
rect 126888 154012 126940 154018
rect 126888 153954 126940 153960
rect 126242 152416 126298 152425
rect 126242 152351 126298 152360
rect 126794 152416 126850 152425
rect 126794 152351 126850 152360
rect 118896 149926 119324 149954
rect 119862 149940 119890 150198
rect 120506 149940 120534 150198
rect 121150 149940 121178 150198
rect 121794 149940 121822 150198
rect 122438 149940 122466 150198
rect 122840 150204 122892 150210
rect 123036 150198 123110 150226
rect 122840 150146 122892 150152
rect 123082 149940 123110 150198
rect 123714 150204 123766 150210
rect 124324 150198 124398 150226
rect 124968 150198 125042 150226
rect 123714 150146 123766 150152
rect 123726 149940 123754 150146
rect 124370 149940 124398 150198
rect 125014 149940 125042 150198
rect 125658 150198 125732 150226
rect 126256 150226 126284 152351
rect 126900 150226 126928 153954
rect 126992 152522 127020 163254
rect 127268 163146 127296 163254
rect 127346 163200 127402 164400
rect 128174 163200 128230 164400
rect 129002 163200 129058 164400
rect 129922 163200 129978 164400
rect 130750 163200 130806 164400
rect 131578 163200 131634 164400
rect 132406 163200 132462 164400
rect 133234 163200 133290 164400
rect 134062 163200 134118 164400
rect 134890 163200 134946 164400
rect 135810 163200 135866 164400
rect 136638 163200 136694 164400
rect 137466 163200 137522 164400
rect 138294 163200 138350 164400
rect 139122 163200 139178 164400
rect 139950 163200 140006 164400
rect 140778 163200 140834 164400
rect 141698 163200 141754 164400
rect 142526 163200 142582 164400
rect 143354 163200 143410 164400
rect 144182 163200 144238 164400
rect 145010 163200 145066 164400
rect 145838 163200 145894 164400
rect 146666 163200 146722 164400
rect 147586 163200 147642 164400
rect 148414 163200 148470 164400
rect 149242 163200 149298 164400
rect 150070 163200 150126 164400
rect 150898 163200 150954 164400
rect 151726 163200 151782 164400
rect 151832 163254 152504 163282
rect 127360 163146 127388 163200
rect 127268 163118 127388 163146
rect 127624 159520 127676 159526
rect 127624 159462 127676 159468
rect 127532 156732 127584 156738
rect 127532 156674 127584 156680
rect 126980 152516 127032 152522
rect 126980 152458 127032 152464
rect 127544 150226 127572 156674
rect 127636 154018 127664 159462
rect 128188 156738 128216 163200
rect 128176 156732 128228 156738
rect 128176 156674 128228 156680
rect 129016 155242 129044 163200
rect 129936 160818 129964 163200
rect 129924 160812 129976 160818
rect 129924 160754 129976 160760
rect 130764 158914 130792 163200
rect 131026 159352 131082 159361
rect 131026 159287 131082 159296
rect 129740 158908 129792 158914
rect 129740 158850 129792 158856
rect 130752 158908 130804 158914
rect 130752 158850 130804 158856
rect 129004 155236 129056 155242
rect 129004 155178 129056 155184
rect 129384 154142 129688 154170
rect 129280 154080 129332 154086
rect 129280 154022 129332 154028
rect 127624 154012 127676 154018
rect 127624 153954 127676 153960
rect 128818 152552 128874 152561
rect 128818 152487 128874 152496
rect 128176 151836 128228 151842
rect 128176 151778 128228 151784
rect 128188 150226 128216 151778
rect 128832 150226 128860 152487
rect 129292 151814 129320 154022
rect 129384 154018 129412 154142
rect 129660 154018 129688 154142
rect 129372 154012 129424 154018
rect 129372 153954 129424 153960
rect 129648 154012 129700 154018
rect 129648 153954 129700 153960
rect 129752 151842 129780 158850
rect 130108 156800 130160 156806
rect 130108 156742 130160 156748
rect 129740 151836 129792 151842
rect 129292 151786 129504 151814
rect 129476 150226 129504 151786
rect 129740 151778 129792 151784
rect 130120 150226 130148 156742
rect 130752 152244 130804 152250
rect 130752 152186 130804 152192
rect 130764 150226 130792 152186
rect 131040 151814 131068 159287
rect 131592 158030 131620 163200
rect 131580 158024 131632 158030
rect 131580 157966 131632 157972
rect 132420 153950 132448 163200
rect 132880 159990 133184 160018
rect 132880 159662 132908 159990
rect 133156 159866 133184 159990
rect 132960 159860 133012 159866
rect 132960 159802 133012 159808
rect 133144 159860 133196 159866
rect 133144 159802 133196 159808
rect 132868 159656 132920 159662
rect 132868 159598 132920 159604
rect 132972 159474 133000 159802
rect 133248 159610 133276 163200
rect 133248 159582 133460 159610
rect 133236 159520 133288 159526
rect 132972 159468 133236 159474
rect 132972 159462 133288 159468
rect 132972 159446 133276 159462
rect 132684 159384 132736 159390
rect 132684 159326 132736 159332
rect 132696 158846 132724 159326
rect 133432 158846 133460 159582
rect 133602 159488 133658 159497
rect 133602 159423 133658 159432
rect 132684 158840 132736 158846
rect 132684 158782 132736 158788
rect 133420 158840 133472 158846
rect 133420 158782 133472 158788
rect 132500 156936 132552 156942
rect 132500 156878 132552 156884
rect 132408 153944 132460 153950
rect 132038 153912 132094 153921
rect 132408 153886 132460 153892
rect 132038 153847 132094 153856
rect 131040 151786 131436 151814
rect 131408 150226 131436 151786
rect 132052 150226 132080 153847
rect 132512 151814 132540 156878
rect 133052 154692 133104 154698
rect 133052 154634 133104 154640
rect 133064 151814 133092 154634
rect 133616 153105 133644 159423
rect 133602 153096 133658 153105
rect 133602 153031 133658 153040
rect 133972 152584 134024 152590
rect 133972 152526 134024 152532
rect 132512 151786 132724 151814
rect 133064 151786 133368 151814
rect 132696 150226 132724 151786
rect 133340 150226 133368 151786
rect 133984 150226 134012 152526
rect 134076 152250 134104 163200
rect 134156 160812 134208 160818
rect 134156 160754 134208 160760
rect 134168 159594 134196 160754
rect 134156 159588 134208 159594
rect 134156 159530 134208 159536
rect 134904 156942 134932 163200
rect 134892 156936 134944 156942
rect 134892 156878 134944 156884
rect 135260 156868 135312 156874
rect 135260 156810 135312 156816
rect 134614 154048 134670 154057
rect 134614 153983 134670 153992
rect 134064 152244 134116 152250
rect 134064 152186 134116 152192
rect 134628 150226 134656 153983
rect 135272 150226 135300 156810
rect 135824 156806 135852 163200
rect 136652 159662 136680 163200
rect 136548 159656 136600 159662
rect 136548 159598 136600 159604
rect 136640 159656 136692 159662
rect 136640 159598 136692 159604
rect 136560 159474 136588 159598
rect 136560 159446 136680 159474
rect 135812 156800 135864 156806
rect 135812 156742 135864 156748
rect 136546 153096 136602 153105
rect 136546 153031 136602 153040
rect 135904 152652 135956 152658
rect 135904 152594 135956 152600
rect 135916 150226 135944 152594
rect 136560 150226 136588 153031
rect 136652 152590 136680 159446
rect 137480 159390 137508 163200
rect 138018 159624 138074 159633
rect 138018 159559 138074 159568
rect 137100 159384 137152 159390
rect 137100 159326 137152 159332
rect 137468 159384 137520 159390
rect 137468 159326 137520 159332
rect 137112 154630 137140 159326
rect 138032 157334 138060 159559
rect 138032 157306 138152 157334
rect 137376 157004 137428 157010
rect 137376 156946 137428 156952
rect 137100 154624 137152 154630
rect 137100 154566 137152 154572
rect 136928 154278 137140 154306
rect 136928 154222 136956 154278
rect 136916 154216 136968 154222
rect 136916 154158 136968 154164
rect 137112 154170 137140 154278
rect 137008 154148 137060 154154
rect 137112 154142 137324 154170
rect 137008 154090 137060 154096
rect 136640 152584 136692 152590
rect 136640 152526 136692 152532
rect 137020 151814 137048 154090
rect 137296 154086 137324 154142
rect 137284 154080 137336 154086
rect 137284 154022 137336 154028
rect 137388 151814 137416 156946
rect 138020 154624 138072 154630
rect 138020 154566 138072 154572
rect 138032 153950 138060 154566
rect 138020 153944 138072 153950
rect 138020 153886 138072 153892
rect 138124 152862 138152 157306
rect 138308 157010 138336 163200
rect 138296 157004 138348 157010
rect 138296 156946 138348 156952
rect 139136 156874 139164 163200
rect 139964 159662 139992 163200
rect 139400 159656 139452 159662
rect 139400 159598 139452 159604
rect 139952 159656 140004 159662
rect 139952 159598 140004 159604
rect 139412 157334 139440 159598
rect 139412 157306 139900 157334
rect 139124 156868 139176 156874
rect 139124 156810 139176 156816
rect 139308 154760 139360 154766
rect 139308 154702 139360 154708
rect 138020 152856 138072 152862
rect 138020 152798 138072 152804
rect 138112 152856 138164 152862
rect 138112 152798 138164 152804
rect 138032 152674 138060 152798
rect 139124 152788 139176 152794
rect 139124 152730 139176 152736
rect 138032 152646 138152 152674
rect 138124 152590 138152 152646
rect 138112 152584 138164 152590
rect 138112 152526 138164 152532
rect 138480 151904 138532 151910
rect 138480 151846 138532 151852
rect 137020 151786 137232 151814
rect 137388 151786 137876 151814
rect 137204 150226 137232 151786
rect 137848 150226 137876 151786
rect 126256 150198 126330 150226
rect 126900 150198 126974 150226
rect 127544 150198 127618 150226
rect 128188 150198 128262 150226
rect 128832 150198 128906 150226
rect 129476 150198 129550 150226
rect 130120 150198 130194 150226
rect 130764 150198 130838 150226
rect 131408 150198 131482 150226
rect 132052 150198 132126 150226
rect 132696 150198 132770 150226
rect 133340 150198 133414 150226
rect 133984 150198 134058 150226
rect 134628 150198 134702 150226
rect 135272 150198 135346 150226
rect 135916 150198 135990 150226
rect 136560 150198 136634 150226
rect 137204 150198 137278 150226
rect 137848 150198 137922 150226
rect 125658 149940 125686 150198
rect 126302 149940 126330 150198
rect 126946 149940 126974 150198
rect 127590 149940 127618 150198
rect 128234 149940 128262 150198
rect 128878 149940 128906 150198
rect 129522 149940 129550 150198
rect 130166 149940 130194 150198
rect 130810 149940 130838 150198
rect 131454 149940 131482 150198
rect 132098 149940 132126 150198
rect 132742 149940 132770 150198
rect 133386 149940 133414 150198
rect 134030 149940 134058 150198
rect 134674 149940 134702 150198
rect 135318 149940 135346 150198
rect 135962 149940 135990 150198
rect 136606 149940 136634 150198
rect 137250 149940 137278 150198
rect 137894 149940 137922 150198
rect 138492 150090 138520 151846
rect 139136 150090 139164 152730
rect 139320 151910 139348 154702
rect 139872 154086 139900 157306
rect 140410 156632 140466 156641
rect 140410 156567 140466 156576
rect 139768 154080 139820 154086
rect 139768 154022 139820 154028
rect 139860 154080 139912 154086
rect 139860 154022 139912 154028
rect 139308 151904 139360 151910
rect 139308 151846 139360 151852
rect 139780 150090 139808 154022
rect 140424 150090 140452 156567
rect 140792 152794 140820 163200
rect 141712 157418 141740 163200
rect 141700 157412 141752 157418
rect 141700 157354 141752 157360
rect 142540 155310 142568 163200
rect 143368 160070 143396 163200
rect 143264 160064 143316 160070
rect 143264 160006 143316 160012
rect 143356 160064 143408 160070
rect 143356 160006 143408 160012
rect 143276 159866 143304 160006
rect 143172 159860 143224 159866
rect 143172 159802 143224 159808
rect 143264 159860 143316 159866
rect 143264 159802 143316 159808
rect 143078 156768 143134 156777
rect 143078 156703 143134 156712
rect 142528 155304 142580 155310
rect 142528 155246 142580 155252
rect 142160 154624 142212 154630
rect 142160 154566 142212 154572
rect 142172 154222 142200 154566
rect 142264 154550 142752 154578
rect 142160 154216 142212 154222
rect 142160 154158 142212 154164
rect 142264 154154 142292 154550
rect 142344 154488 142396 154494
rect 142344 154430 142396 154436
rect 142436 154488 142488 154494
rect 142488 154436 142660 154442
rect 142436 154430 142660 154436
rect 142356 154204 142384 154430
rect 142448 154426 142660 154430
rect 142448 154420 142672 154426
rect 142448 154414 142620 154420
rect 142620 154362 142672 154368
rect 142724 154358 142752 154550
rect 142712 154352 142764 154358
rect 142712 154294 142764 154300
rect 142620 154284 142672 154290
rect 142620 154226 142672 154232
rect 142896 154284 142948 154290
rect 142896 154226 142948 154232
rect 142356 154176 142568 154204
rect 142252 154148 142304 154154
rect 142252 154090 142304 154096
rect 142540 154086 142568 154176
rect 142632 154154 142660 154226
rect 142908 154170 142936 154226
rect 142620 154148 142672 154154
rect 142620 154090 142672 154096
rect 142724 154142 142936 154170
rect 142436 154080 142488 154086
rect 142250 154048 142306 154057
rect 142434 154048 142436 154057
rect 142528 154080 142580 154086
rect 142488 154048 142490 154057
rect 142306 154006 142384 154034
rect 142250 153983 142306 153992
rect 141700 152856 141752 152862
rect 141700 152798 141752 152804
rect 140780 152788 140832 152794
rect 140780 152730 140832 152736
rect 141056 152720 141108 152726
rect 141056 152662 141108 152668
rect 141068 150090 141096 152662
rect 141712 150090 141740 152798
rect 142356 150226 142384 154006
rect 142528 154022 142580 154028
rect 142434 153983 142490 153992
rect 142724 153270 142752 154142
rect 142986 154048 143042 154057
rect 142986 153983 143042 153992
rect 143000 153950 143028 153983
rect 142988 153944 143040 153950
rect 142988 153886 143040 153892
rect 142804 153876 142856 153882
rect 142804 153818 142856 153824
rect 142816 153270 142844 153818
rect 142712 153264 142764 153270
rect 142712 153206 142764 153212
rect 142804 153264 142856 153270
rect 142804 153206 142856 153212
rect 142804 152720 142856 152726
rect 142804 152662 142856 152668
rect 142816 152046 142844 152662
rect 142804 152040 142856 152046
rect 142804 151982 142856 151988
rect 142356 150198 142430 150226
rect 138492 150062 138566 150090
rect 139136 150062 139210 150090
rect 139780 150062 139854 150090
rect 140424 150062 140498 150090
rect 141068 150062 141142 150090
rect 141712 150062 141786 150090
rect 138538 149940 138566 150062
rect 139182 149940 139210 150062
rect 139826 149940 139854 150062
rect 140470 149940 140498 150062
rect 141114 149940 141142 150062
rect 141758 149940 141786 150062
rect 142402 149940 142430 150198
rect 143092 150090 143120 156703
rect 143184 152046 143212 159802
rect 144196 159526 144224 163200
rect 144092 159520 144144 159526
rect 144092 159462 144144 159468
rect 144184 159520 144236 159526
rect 144184 159462 144236 159468
rect 144104 159338 144132 159462
rect 144104 159310 144408 159338
rect 144380 152794 144408 159310
rect 145024 155990 145052 163200
rect 145102 157992 145158 158001
rect 145102 157927 145158 157936
rect 145012 155984 145064 155990
rect 145012 155926 145064 155932
rect 144276 152788 144328 152794
rect 144276 152730 144328 152736
rect 144368 152788 144420 152794
rect 144368 152730 144420 152736
rect 144288 152674 144316 152730
rect 144288 152646 144408 152674
rect 144380 152590 144408 152646
rect 144276 152584 144328 152590
rect 144276 152526 144328 152532
rect 144368 152584 144420 152590
rect 144368 152526 144420 152532
rect 143630 152416 143686 152425
rect 143630 152351 143686 152360
rect 143172 152040 143224 152046
rect 143172 151982 143224 151988
rect 143046 150062 143120 150090
rect 143644 150090 143672 152351
rect 144288 150090 144316 152526
rect 145116 150226 145144 157927
rect 145852 155378 145880 163200
rect 146680 159866 146708 163200
rect 146576 159860 146628 159866
rect 146576 159802 146628 159808
rect 146668 159860 146720 159866
rect 146668 159802 146720 159808
rect 146392 158092 146444 158098
rect 146392 158034 146444 158040
rect 146208 157072 146260 157078
rect 146208 157014 146260 157020
rect 145840 155372 145892 155378
rect 145840 155314 145892 155320
rect 145564 154148 145616 154154
rect 145564 154090 145616 154096
rect 144978 150198 145144 150226
rect 143644 150062 143718 150090
rect 144288 150062 144362 150090
rect 143046 149940 143074 150062
rect 143690 149940 143718 150062
rect 144334 149940 144362 150062
rect 144978 149940 145006 150198
rect 145576 150090 145604 154090
rect 146220 150090 146248 157014
rect 146404 150210 146432 158034
rect 146588 152862 146616 159802
rect 147600 158778 147628 163200
rect 147772 159452 147824 159458
rect 147772 159394 147824 159400
rect 147128 158772 147180 158778
rect 147128 158714 147180 158720
rect 147588 158772 147640 158778
rect 147588 158714 147640 158720
rect 147140 154154 147168 158714
rect 147784 154222 147812 159394
rect 148428 158098 148456 163200
rect 148416 158092 148468 158098
rect 148416 158034 148468 158040
rect 148784 157140 148836 157146
rect 148784 157082 148836 157088
rect 147588 154216 147640 154222
rect 147586 154184 147588 154193
rect 147772 154216 147824 154222
rect 147640 154184 147642 154193
rect 147128 154148 147180 154154
rect 147772 154158 147824 154164
rect 148138 154184 148194 154193
rect 147586 154119 147642 154128
rect 148138 154119 148194 154128
rect 147128 154090 147180 154096
rect 146576 152856 146628 152862
rect 146576 152798 146628 152804
rect 146944 152040 146996 152046
rect 146944 151982 146996 151988
rect 146956 151842 146984 151982
rect 146852 151836 146904 151842
rect 146852 151778 146904 151784
rect 146944 151836 146996 151842
rect 146944 151778 146996 151784
rect 146392 150204 146444 150210
rect 146392 150146 146444 150152
rect 146864 150090 146892 151778
rect 147542 150204 147594 150210
rect 147542 150146 147594 150152
rect 145576 150062 145650 150090
rect 146220 150062 146294 150090
rect 146864 150062 146938 150090
rect 145622 149940 145650 150062
rect 146266 149940 146294 150062
rect 146910 149940 146938 150062
rect 147554 149940 147582 150146
rect 148152 150090 148180 154119
rect 148796 150090 148824 157082
rect 149256 155446 149284 163200
rect 149520 158772 149572 158778
rect 149520 158714 149572 158720
rect 149244 155440 149296 155446
rect 149244 155382 149296 155388
rect 149532 152726 149560 158714
rect 149610 158264 149666 158273
rect 149610 158199 149666 158208
rect 149624 157334 149652 158199
rect 149624 157306 150020 157334
rect 149428 152720 149480 152726
rect 149428 152662 149480 152668
rect 149520 152720 149572 152726
rect 149520 152662 149572 152668
rect 149440 150090 149468 152662
rect 149992 150226 150020 157306
rect 150084 157146 150112 163200
rect 150912 159458 150940 163200
rect 150900 159452 150952 159458
rect 150900 159394 150952 159400
rect 151268 157208 151320 157214
rect 151268 157150 151320 157156
rect 150072 157140 150124 157146
rect 150072 157082 150124 157088
rect 150624 154284 150676 154290
rect 150624 154226 150676 154232
rect 149992 150198 150066 150226
rect 148152 150062 148226 150090
rect 148796 150062 148870 150090
rect 149440 150062 149514 150090
rect 148198 149940 148226 150062
rect 148842 149940 148870 150062
rect 149486 149940 149514 150062
rect 150038 149940 150066 150198
rect 150636 150090 150664 154226
rect 151280 150226 151308 157150
rect 151740 157078 151768 163200
rect 151728 157072 151780 157078
rect 151728 157014 151780 157020
rect 151832 154766 151860 163254
rect 152476 163146 152504 163254
rect 152554 163200 152610 164400
rect 153474 163200 153530 164400
rect 153580 163254 154252 163282
rect 152568 163146 152596 163200
rect 152476 163118 152596 163146
rect 153488 158778 153516 163200
rect 153476 158772 153528 158778
rect 153476 158714 153528 158720
rect 152554 158128 152610 158137
rect 152554 158063 152610 158072
rect 151820 154760 151872 154766
rect 151820 154702 151872 154708
rect 152372 154284 152424 154290
rect 152372 154226 152424 154232
rect 152384 153678 152412 154226
rect 152464 153876 152516 153882
rect 152464 153818 152516 153824
rect 152476 153678 152504 153818
rect 152372 153672 152424 153678
rect 152372 153614 152424 153620
rect 152464 153672 152516 153678
rect 152464 153614 152516 153620
rect 151912 152652 151964 152658
rect 151912 152594 151964 152600
rect 151280 150198 151354 150226
rect 150636 150062 150710 150090
rect 150682 149940 150710 150062
rect 151326 149940 151354 150198
rect 151924 150090 151952 152594
rect 152568 150226 152596 158063
rect 153108 154760 153160 154766
rect 153108 154702 153160 154708
rect 153120 154170 153148 154702
rect 153120 154142 153332 154170
rect 153304 154086 153332 154142
rect 153200 154080 153252 154086
rect 153200 154022 153252 154028
rect 153292 154080 153344 154086
rect 153292 154022 153344 154028
rect 152568 150198 152642 150226
rect 151924 150062 151998 150090
rect 151970 149940 151998 150062
rect 152614 149940 152642 150198
rect 153212 150090 153240 154022
rect 153580 152658 153608 163254
rect 154224 163146 154252 163254
rect 154302 163200 154358 164400
rect 155130 163200 155186 164400
rect 155958 163200 156014 164400
rect 156786 163200 156842 164400
rect 157614 163200 157670 164400
rect 158442 163200 158498 164400
rect 159362 163200 159418 164400
rect 160190 163200 160246 164400
rect 161018 163200 161074 164400
rect 161846 163200 161902 164400
rect 162674 163200 162730 164400
rect 163502 163200 163558 164400
rect 164330 163200 164386 164400
rect 165250 163200 165306 164400
rect 165632 163254 166028 163282
rect 154316 163146 154344 163200
rect 154224 163118 154344 163146
rect 154488 159588 154540 159594
rect 154488 159530 154540 159536
rect 153844 157276 153896 157282
rect 153844 157218 153896 157224
rect 153568 152652 153620 152658
rect 153568 152594 153620 152600
rect 153856 150090 153884 157218
rect 154500 153882 154528 159530
rect 155144 158234 155172 163200
rect 155040 158228 155092 158234
rect 155040 158170 155092 158176
rect 155132 158228 155184 158234
rect 155132 158170 155184 158176
rect 155052 157334 155080 158170
rect 155052 157306 155172 157334
rect 154488 153876 154540 153882
rect 154488 153818 154540 153824
rect 154488 151972 154540 151978
rect 154488 151914 154540 151920
rect 154500 150090 154528 151914
rect 155144 150226 155172 157306
rect 155972 154766 156000 163200
rect 156800 160070 156828 163200
rect 156604 160064 156656 160070
rect 156604 160006 156656 160012
rect 156788 160064 156840 160070
rect 156788 160006 156840 160012
rect 156616 159798 156644 160006
rect 156328 159792 156380 159798
rect 156328 159734 156380 159740
rect 156604 159792 156656 159798
rect 156604 159734 156656 159740
rect 155960 154760 156012 154766
rect 155960 154702 156012 154708
rect 155960 154080 156012 154086
rect 155960 154022 156012 154028
rect 155972 153882 156000 154022
rect 155960 153876 156012 153882
rect 155960 153818 156012 153824
rect 155776 153808 155828 153814
rect 155776 153750 155828 153756
rect 155144 150198 155218 150226
rect 153212 150062 153286 150090
rect 153856 150062 153930 150090
rect 154500 150062 154574 150090
rect 153258 149940 153286 150062
rect 153902 149940 153930 150062
rect 154546 149940 154574 150062
rect 155190 149940 155218 150198
rect 155788 150090 155816 153750
rect 156340 152046 156368 159734
rect 156512 159724 156564 159730
rect 156512 159666 156564 159672
rect 156420 157344 156472 157350
rect 156420 157286 156472 157292
rect 156328 152040 156380 152046
rect 156328 151982 156380 151988
rect 156432 150090 156460 157286
rect 156524 157214 156552 159666
rect 157628 159594 157656 163200
rect 157616 159588 157668 159594
rect 157616 159530 157668 159536
rect 158456 158166 158484 163200
rect 158720 158840 158772 158846
rect 158720 158782 158772 158788
rect 157708 158160 157760 158166
rect 157708 158102 157760 158108
rect 158444 158160 158496 158166
rect 158444 158102 158496 158108
rect 156512 157208 156564 157214
rect 156512 157150 156564 157156
rect 157340 154692 157392 154698
rect 157340 154634 157392 154640
rect 157248 154556 157300 154562
rect 157248 154498 157300 154504
rect 157260 154222 157288 154498
rect 157352 154222 157380 154634
rect 157248 154216 157300 154222
rect 157248 154158 157300 154164
rect 157340 154216 157392 154222
rect 157340 154158 157392 154164
rect 157064 151836 157116 151842
rect 157064 151778 157116 151784
rect 157076 150090 157104 151778
rect 157720 150226 157748 158102
rect 158732 157350 158760 158782
rect 158720 157344 158772 157350
rect 158720 157286 158772 157292
rect 159088 157208 159140 157214
rect 159088 157150 159140 157156
rect 159100 156602 159128 157150
rect 158996 156596 159048 156602
rect 158996 156538 159048 156544
rect 159088 156596 159140 156602
rect 159088 156538 159140 156544
rect 158352 154216 158404 154222
rect 158352 154158 158404 154164
rect 158364 150226 158392 154158
rect 159008 150226 159036 156538
rect 159376 154630 159404 163200
rect 160100 159792 160152 159798
rect 160100 159734 160152 159740
rect 160112 157214 160140 159734
rect 160100 157208 160152 157214
rect 160100 157150 160152 157156
rect 159364 154624 159416 154630
rect 159364 154566 159416 154572
rect 160204 154154 160232 163200
rect 161032 159662 161060 163200
rect 161020 159656 161072 159662
rect 161020 159598 161072 159604
rect 161860 158302 161888 163200
rect 162492 159928 162544 159934
rect 162492 159870 162544 159876
rect 160284 158296 160336 158302
rect 160284 158238 160336 158244
rect 161848 158296 161900 158302
rect 161848 158238 161900 158244
rect 160192 154148 160244 154154
rect 160192 154090 160244 154096
rect 159640 152448 159692 152454
rect 159640 152390 159692 152396
rect 159652 150226 159680 152390
rect 160296 150226 160324 158238
rect 161662 156904 161718 156913
rect 161662 156839 161718 156848
rect 160926 154320 160982 154329
rect 160926 154255 160982 154264
rect 160940 150226 160968 154255
rect 161480 154216 161532 154222
rect 161480 154158 161532 154164
rect 161492 153746 161520 154158
rect 161572 154080 161624 154086
rect 161572 154022 161624 154028
rect 161584 153746 161612 154022
rect 161480 153740 161532 153746
rect 161480 153682 161532 153688
rect 161572 153740 161624 153746
rect 161572 153682 161624 153688
rect 161676 150226 161704 156839
rect 162216 152788 162268 152794
rect 162216 152730 162268 152736
rect 157720 150198 157794 150226
rect 158364 150198 158438 150226
rect 159008 150198 159082 150226
rect 159652 150198 159726 150226
rect 160296 150198 160370 150226
rect 160940 150198 161014 150226
rect 155788 150062 155862 150090
rect 156432 150062 156506 150090
rect 157076 150062 157150 150090
rect 155834 149940 155862 150062
rect 156478 149940 156506 150062
rect 157122 149940 157150 150062
rect 157766 149940 157794 150198
rect 158410 149940 158438 150198
rect 159054 149940 159082 150198
rect 159698 149940 159726 150198
rect 160342 149940 160370 150198
rect 160986 149940 161014 150198
rect 161630 150198 161704 150226
rect 162228 150226 162256 152730
rect 162504 151978 162532 159870
rect 162688 154698 162716 163200
rect 162872 159186 163084 159202
rect 162872 159180 163096 159186
rect 162872 159174 163044 159180
rect 162872 159118 162900 159174
rect 163044 159122 163096 159128
rect 162860 159112 162912 159118
rect 162860 159054 162912 159060
rect 163516 158846 163544 163200
rect 164344 161474 164372 163200
rect 164344 161446 164464 161474
rect 163780 159724 163832 159730
rect 163780 159666 163832 159672
rect 163504 158840 163556 158846
rect 163504 158782 163556 158788
rect 162858 158400 162914 158409
rect 162858 158335 162914 158344
rect 162676 154692 162728 154698
rect 162676 154634 162728 154640
rect 162492 151972 162544 151978
rect 162492 151914 162544 151920
rect 162872 150226 162900 158335
rect 163792 157282 163820 159666
rect 164332 158432 164384 158438
rect 164332 158374 164384 158380
rect 163780 157276 163832 157282
rect 163780 157218 163832 157224
rect 164148 156528 164200 156534
rect 164148 156470 164200 156476
rect 163504 154284 163556 154290
rect 163504 154226 163556 154232
rect 163516 150226 163544 154226
rect 164160 150226 164188 156470
rect 162228 150198 162302 150226
rect 162872 150198 162946 150226
rect 163516 150198 163590 150226
rect 164160 150198 164234 150226
rect 164344 150210 164372 158374
rect 164436 152794 164464 161446
rect 165264 158438 165292 163200
rect 165252 158432 165304 158438
rect 165252 158374 165304 158380
rect 165632 154154 165660 163254
rect 166000 163146 166028 163254
rect 166078 163200 166134 164400
rect 166906 163200 166962 164400
rect 167734 163200 167790 164400
rect 168562 163200 168618 164400
rect 169390 163200 169446 164400
rect 170218 163200 170274 164400
rect 171138 163200 171194 164400
rect 171966 163200 172022 164400
rect 172532 163254 172744 163282
rect 166092 163146 166120 163200
rect 166000 163118 166120 163146
rect 166920 159934 166948 163200
rect 166908 159928 166960 159934
rect 166908 159870 166960 159876
rect 167748 159730 167776 163200
rect 167736 159724 167788 159730
rect 167736 159666 167788 159672
rect 167000 159316 167052 159322
rect 167000 159258 167052 159264
rect 166448 157276 166500 157282
rect 166448 157218 166500 157224
rect 166172 157208 166224 157214
rect 166172 157150 166224 157156
rect 166264 157208 166316 157214
rect 166264 157150 166316 157156
rect 166184 156534 166212 157150
rect 166172 156528 166224 156534
rect 166172 156470 166224 156476
rect 166276 156466 166304 157150
rect 166460 156534 166488 157218
rect 166448 156528 166500 156534
rect 166448 156470 166500 156476
rect 166264 156460 166316 156466
rect 166264 156402 166316 156408
rect 166722 155544 166778 155553
rect 166722 155479 166778 155488
rect 166080 154216 166132 154222
rect 166080 154158 166132 154164
rect 165620 154148 165672 154154
rect 165620 154090 165672 154096
rect 164424 152788 164476 152794
rect 164424 152730 164476 152736
rect 164792 152108 164844 152114
rect 164792 152050 164844 152056
rect 164804 150226 164832 152050
rect 166092 150226 166120 154158
rect 166736 150226 166764 155479
rect 167012 152114 167040 159258
rect 168576 158370 168604 163200
rect 167552 158364 167604 158370
rect 167552 158306 167604 158312
rect 168564 158364 168616 158370
rect 168564 158306 168616 158312
rect 167368 152856 167420 152862
rect 167368 152798 167420 152804
rect 167000 152108 167052 152114
rect 167000 152050 167052 152056
rect 167380 150226 167408 152798
rect 167564 151814 167592 158306
rect 169404 155514 169432 163200
rect 170232 159322 170260 163200
rect 170220 159316 170272 159322
rect 170220 159258 170272 159264
rect 171152 159118 171180 163200
rect 169760 159112 169812 159118
rect 169760 159054 169812 159060
rect 171140 159112 171192 159118
rect 171140 159054 171192 159060
rect 168656 155508 168708 155514
rect 168656 155450 168708 155456
rect 169392 155508 169444 155514
rect 169392 155450 169444 155456
rect 168378 155272 168434 155281
rect 168378 155207 168434 155216
rect 167564 151786 168052 151814
rect 168024 150226 168052 151786
rect 161630 149940 161658 150198
rect 162274 149940 162302 150198
rect 162918 149940 162946 150198
rect 163562 149940 163590 150198
rect 164206 149940 164234 150198
rect 164332 150204 164384 150210
rect 164804 150198 164878 150226
rect 164332 150146 164384 150152
rect 164850 149940 164878 150198
rect 165482 150204 165534 150210
rect 166092 150198 166166 150226
rect 166736 150198 166810 150226
rect 167380 150198 167454 150226
rect 168024 150198 168098 150226
rect 168392 150210 168420 155207
rect 168668 150226 168696 155450
rect 169772 151842 169800 159054
rect 171980 158642 172008 163200
rect 172152 159180 172204 159186
rect 172152 159122 172204 159128
rect 170312 158636 170364 158642
rect 170312 158578 170364 158584
rect 171968 158636 172020 158642
rect 171968 158578 172020 158584
rect 169944 152176 169996 152182
rect 169944 152118 169996 152124
rect 169760 151836 169812 151842
rect 169760 151778 169812 151784
rect 169956 150226 169984 152118
rect 170324 151814 170352 158578
rect 171140 157208 171192 157214
rect 171140 157150 171192 157156
rect 170324 151786 170628 151814
rect 170600 150226 170628 151786
rect 165482 150146 165534 150152
rect 165494 149940 165522 150146
rect 166138 149940 166166 150198
rect 166782 149940 166810 150198
rect 167426 149940 167454 150198
rect 168070 149940 168098 150198
rect 168380 150204 168432 150210
rect 168668 150198 168742 150226
rect 168380 150146 168432 150152
rect 168714 149940 168742 150198
rect 169346 150204 169398 150210
rect 169956 150198 170030 150226
rect 170600 150198 170674 150226
rect 171152 150210 171180 157150
rect 171230 155408 171286 155417
rect 171230 155343 171286 155352
rect 171244 150226 171272 155343
rect 172164 152182 172192 159122
rect 172532 154222 172560 163254
rect 172716 163146 172744 163254
rect 172794 163200 172850 164400
rect 173622 163200 173678 164400
rect 173912 163254 174400 163282
rect 172808 163146 172836 163200
rect 172716 163118 172836 163146
rect 173636 159186 173664 163200
rect 173624 159180 173676 159186
rect 173624 159122 173676 159128
rect 173164 159112 173216 159118
rect 173164 159054 173216 159060
rect 173072 158500 173124 158506
rect 173072 158442 173124 158448
rect 172704 155644 172756 155650
rect 172704 155586 172756 155592
rect 172520 154216 172572 154222
rect 172520 154158 172572 154164
rect 172152 152176 172204 152182
rect 172152 152118 172204 152124
rect 172520 152040 172572 152046
rect 172520 151982 172572 151988
rect 172532 150226 172560 151982
rect 169346 150146 169398 150152
rect 169358 149940 169386 150146
rect 170002 149940 170030 150198
rect 170646 149940 170674 150198
rect 171140 150204 171192 150210
rect 171244 150198 171318 150226
rect 171140 150146 171192 150152
rect 171290 149940 171318 150198
rect 171922 150204 171974 150210
rect 172532 150198 172606 150226
rect 172716 150210 172744 155586
rect 173084 151814 173112 158442
rect 173176 152454 173204 159054
rect 173912 152862 173940 163254
rect 174372 163146 174400 163254
rect 174450 163200 174506 164400
rect 175278 163200 175334 164400
rect 176106 163200 176162 164400
rect 177026 163200 177082 164400
rect 177854 163200 177910 164400
rect 178682 163200 178738 164400
rect 179510 163200 179566 164400
rect 180338 163200 180394 164400
rect 180812 163254 181116 163282
rect 174464 163146 174492 163200
rect 174372 163118 174492 163146
rect 175292 158574 175320 163200
rect 176120 161474 176148 163200
rect 176120 161446 176332 161474
rect 175280 158568 175332 158574
rect 175280 158510 175332 158516
rect 175372 158500 175424 158506
rect 175372 158442 175424 158448
rect 174450 157040 174506 157049
rect 174450 156975 174506 156984
rect 173900 152856 173952 152862
rect 173900 152798 173952 152804
rect 173164 152448 173216 152454
rect 173164 152390 173216 152396
rect 173084 151786 173204 151814
rect 173176 150226 173204 151786
rect 174464 150226 174492 156975
rect 175096 153128 175148 153134
rect 175096 153070 175148 153076
rect 175108 150226 175136 153070
rect 175384 151814 175412 158442
rect 176200 157956 176252 157962
rect 176200 157898 176252 157904
rect 175924 157888 175976 157894
rect 176212 157842 176240 157898
rect 175976 157836 176240 157842
rect 175924 157830 176240 157836
rect 175936 157814 176240 157830
rect 176304 155650 176332 161446
rect 176660 159860 176712 159866
rect 176660 159802 176712 159808
rect 176292 155644 176344 155650
rect 176292 155586 176344 155592
rect 176384 155576 176436 155582
rect 176384 155518 176436 155524
rect 175384 151786 175780 151814
rect 175752 150226 175780 151786
rect 176396 150226 176424 155518
rect 176672 154290 176700 159802
rect 177040 157214 177068 163200
rect 177868 159798 177896 163200
rect 177856 159792 177908 159798
rect 177856 159734 177908 159740
rect 178696 158506 178724 163200
rect 179420 158772 179472 158778
rect 179420 158714 179472 158720
rect 178684 158500 178736 158506
rect 178684 158442 178736 158448
rect 179432 157894 179460 158714
rect 178040 157888 178092 157894
rect 178040 157830 178092 157836
rect 179420 157888 179472 157894
rect 179420 157830 179472 157836
rect 177028 157208 177080 157214
rect 177028 157150 177080 157156
rect 177026 155816 177082 155825
rect 177026 155751 177082 155760
rect 176660 154284 176712 154290
rect 176660 154226 176712 154232
rect 177040 150226 177068 155751
rect 177672 151972 177724 151978
rect 177672 151914 177724 151920
rect 177684 150226 177712 151914
rect 178052 151814 178080 157830
rect 178958 155680 179014 155689
rect 178958 155615 179014 155624
rect 178052 151786 178356 151814
rect 178328 150226 178356 151786
rect 178972 150226 179000 155615
rect 179524 155582 179552 163200
rect 180352 159118 180380 163200
rect 180340 159112 180392 159118
rect 180340 159054 180392 159060
rect 179512 155576 179564 155582
rect 179512 155518 179564 155524
rect 179696 154284 179748 154290
rect 179696 154226 179748 154232
rect 179708 153610 179736 154226
rect 179604 153604 179656 153610
rect 179604 153546 179656 153552
rect 179696 153604 179748 153610
rect 179696 153546 179748 153552
rect 179616 150226 179644 153546
rect 180812 153134 180840 163254
rect 181088 163146 181116 163254
rect 181166 163200 181222 164400
rect 181994 163200 182050 164400
rect 182192 163254 182864 163282
rect 181180 163146 181208 163200
rect 181088 163118 181208 163146
rect 182008 158710 182036 163200
rect 180892 158704 180944 158710
rect 180892 158646 180944 158652
rect 181996 158704 182048 158710
rect 181996 158646 182048 158652
rect 180800 153128 180852 153134
rect 180800 153070 180852 153076
rect 180248 152312 180300 152318
rect 180248 152254 180300 152260
rect 180260 150226 180288 152254
rect 180904 150226 180932 158646
rect 182088 156392 182140 156398
rect 182088 156334 182140 156340
rect 180984 155712 181036 155718
rect 180984 155654 181036 155660
rect 180996 151814 181024 155654
rect 180996 151786 181484 151814
rect 171922 150146 171974 150152
rect 171934 149940 171962 150146
rect 172578 149940 172606 150198
rect 172704 150204 172756 150210
rect 173176 150198 173250 150226
rect 172704 150146 172756 150152
rect 173222 149940 173250 150198
rect 173854 150204 173906 150210
rect 174464 150198 174538 150226
rect 175108 150198 175182 150226
rect 175752 150198 175826 150226
rect 176396 150198 176470 150226
rect 177040 150198 177114 150226
rect 177684 150198 177758 150226
rect 178328 150198 178402 150226
rect 178972 150198 179046 150226
rect 179616 150198 179690 150226
rect 180260 150198 180334 150226
rect 173854 150146 173906 150152
rect 173866 149940 173894 150146
rect 174510 149940 174538 150198
rect 175154 149940 175182 150198
rect 175798 149940 175826 150198
rect 176442 149940 176470 150198
rect 177086 149940 177114 150198
rect 177730 149940 177758 150198
rect 178374 149940 178402 150198
rect 179018 149940 179046 150198
rect 179662 149940 179690 150198
rect 180306 149940 180334 150198
rect 180858 150198 180932 150226
rect 181456 150226 181484 151786
rect 182100 150226 182128 156334
rect 182192 154290 182220 163254
rect 182836 163146 182864 163254
rect 182914 163200 182970 164400
rect 183742 163200 183798 164400
rect 184570 163200 184626 164400
rect 185398 163200 185454 164400
rect 186226 163200 186282 164400
rect 187054 163200 187110 164400
rect 187882 163200 187938 164400
rect 188802 163200 188858 164400
rect 189630 163200 189686 164400
rect 190458 163200 190514 164400
rect 191286 163200 191342 164400
rect 192114 163200 192170 164400
rect 192942 163200 192998 164400
rect 193770 163200 193826 164400
rect 194690 163200 194746 164400
rect 195518 163200 195574 164400
rect 196346 163200 196402 164400
rect 197174 163200 197230 164400
rect 198002 163200 198058 164400
rect 198830 163200 198886 164400
rect 199658 163200 199714 164400
rect 200578 163200 200634 164400
rect 201406 163200 201462 164400
rect 202234 163200 202290 164400
rect 203062 163200 203118 164400
rect 203890 163200 203946 164400
rect 204718 163200 204774 164400
rect 205008 163254 205496 163282
rect 182928 163146 182956 163200
rect 182836 163118 182956 163146
rect 183756 159050 183784 163200
rect 184584 159866 184612 163200
rect 184572 159860 184624 159866
rect 184572 159802 184624 159808
rect 184388 159248 184440 159254
rect 184388 159190 184440 159196
rect 183468 159044 183520 159050
rect 183468 158986 183520 158992
rect 183744 159044 183796 159050
rect 183744 158986 183796 158992
rect 182272 157956 182324 157962
rect 182272 157898 182324 157904
rect 182180 154284 182232 154290
rect 182180 154226 182232 154232
rect 181456 150198 181530 150226
rect 182100 150198 182174 150226
rect 182284 150210 182312 157898
rect 183480 152114 183508 158986
rect 184018 155952 184074 155961
rect 184018 155887 184074 155896
rect 182732 152108 182784 152114
rect 182732 152050 182784 152056
rect 183468 152108 183520 152114
rect 183468 152050 183520 152056
rect 182744 150226 182772 152050
rect 184032 150226 184060 155887
rect 184400 151978 184428 159190
rect 185412 157962 185440 163200
rect 185400 157956 185452 157962
rect 185400 157898 185452 157904
rect 184940 157888 184992 157894
rect 184768 157836 184940 157842
rect 185952 157888 186004 157894
rect 184768 157830 184992 157836
rect 184768 157826 184980 157830
rect 184756 157820 184980 157826
rect 184808 157814 184980 157820
rect 185216 157820 185268 157826
rect 184756 157762 184808 157768
rect 185216 157762 185268 157768
rect 185320 157814 185716 157842
rect 185952 157830 186004 157836
rect 185228 157570 185256 157762
rect 185320 157758 185348 157814
rect 185688 157758 185716 157814
rect 185308 157752 185360 157758
rect 185308 157694 185360 157700
rect 185676 157752 185728 157758
rect 185676 157694 185728 157700
rect 185584 157684 185636 157690
rect 185584 157626 185636 157632
rect 185596 157570 185624 157626
rect 185228 157542 185624 157570
rect 184662 154456 184718 154465
rect 184662 154391 184718 154400
rect 184388 151972 184440 151978
rect 184388 151914 184440 151920
rect 184676 150226 184704 154391
rect 185308 151836 185360 151842
rect 185308 151778 185360 151784
rect 185320 150226 185348 151778
rect 185964 150226 185992 157830
rect 186240 155718 186268 163200
rect 186688 159928 186740 159934
rect 186688 159870 186740 159876
rect 186700 157334 186728 159870
rect 187068 159254 187096 163200
rect 187896 161474 187924 163200
rect 187896 161446 188016 161474
rect 187056 159248 187108 159254
rect 187056 159190 187108 159196
rect 186700 157306 186912 157334
rect 186412 155916 186464 155922
rect 186412 155858 186464 155864
rect 186228 155712 186280 155718
rect 186228 155654 186280 155660
rect 186424 150226 186452 155858
rect 186780 155848 186832 155854
rect 186780 155790 186832 155796
rect 186792 155700 186820 155790
rect 186516 155672 186820 155700
rect 186516 155106 186544 155672
rect 186884 155106 186912 157306
rect 187240 155168 187292 155174
rect 187240 155110 187292 155116
rect 186504 155100 186556 155106
rect 186504 155042 186556 155048
rect 186872 155100 186924 155106
rect 186872 155042 186924 155048
rect 180858 149940 180886 150198
rect 181502 149940 181530 150198
rect 182146 149940 182174 150198
rect 182272 150204 182324 150210
rect 182744 150198 182818 150226
rect 182272 150146 182324 150152
rect 182790 149940 182818 150198
rect 183422 150204 183474 150210
rect 184032 150198 184106 150226
rect 184676 150198 184750 150226
rect 185320 150198 185394 150226
rect 185964 150198 186038 150226
rect 186424 150198 186682 150226
rect 183422 150146 183474 150152
rect 183434 149940 183462 150146
rect 184078 149940 184106 150198
rect 184722 149940 184750 150198
rect 185366 149940 185394 150198
rect 186010 149940 186038 150198
rect 186654 149940 186682 150198
rect 187252 150090 187280 155110
rect 187884 152992 187936 152998
rect 187884 152934 187936 152940
rect 187896 150090 187924 152934
rect 187988 152318 188016 161446
rect 188816 157894 188844 163200
rect 188804 157888 188856 157894
rect 188804 157830 188856 157836
rect 188528 157752 188580 157758
rect 188528 157694 188580 157700
rect 187976 152312 188028 152318
rect 187976 152254 188028 152260
rect 188540 150226 188568 157694
rect 189172 155916 189224 155922
rect 189172 155858 189224 155864
rect 188540 150198 188614 150226
rect 187252 150062 187326 150090
rect 187896 150062 187970 150090
rect 187298 149940 187326 150062
rect 187942 149940 187970 150062
rect 188586 149940 188614 150198
rect 189184 150090 189212 155858
rect 189644 155174 189672 163200
rect 190472 157758 190500 163200
rect 191300 159934 191328 163200
rect 191748 160064 191800 160070
rect 191748 160006 191800 160012
rect 191472 159996 191524 160002
rect 191472 159938 191524 159944
rect 191288 159928 191340 159934
rect 191288 159870 191340 159876
rect 190644 157820 190696 157826
rect 190644 157762 190696 157768
rect 190460 157752 190512 157758
rect 190460 157694 190512 157700
rect 190656 157334 190684 157762
rect 190656 157306 191144 157334
rect 189632 155168 189684 155174
rect 189632 155110 189684 155116
rect 190748 155094 191052 155122
rect 190748 154970 190776 155094
rect 190828 155032 190880 155038
rect 190828 154974 190880 154980
rect 190920 155032 190972 155038
rect 190920 154974 190972 154980
rect 190736 154964 190788 154970
rect 190736 154906 190788 154912
rect 189816 154420 189868 154426
rect 189816 154362 189868 154368
rect 189828 150090 189856 154362
rect 190460 152176 190512 152182
rect 190460 152118 190512 152124
rect 190472 150090 190500 152118
rect 190840 150210 190868 154974
rect 190932 154902 190960 154974
rect 191024 154970 191052 155094
rect 191012 154964 191064 154970
rect 191012 154906 191064 154912
rect 190920 154896 190972 154902
rect 190920 154838 190972 154844
rect 190920 154488 190972 154494
rect 190918 154456 190920 154465
rect 191012 154488 191064 154494
rect 190972 154456 190974 154465
rect 191012 154430 191064 154436
rect 190918 154391 190974 154400
rect 191024 153678 191052 154430
rect 191012 153672 191064 153678
rect 191012 153614 191064 153620
rect 191116 150226 191144 157306
rect 191196 155100 191248 155106
rect 191196 155042 191248 155048
rect 191208 154902 191236 155042
rect 191196 154896 191248 154902
rect 191196 154838 191248 154844
rect 191286 154456 191342 154465
rect 191196 154420 191248 154426
rect 191286 154391 191342 154400
rect 191196 154362 191248 154368
rect 191208 153406 191236 154362
rect 191300 153406 191328 154391
rect 191196 153400 191248 153406
rect 191196 153342 191248 153348
rect 191288 153400 191340 153406
rect 191288 153342 191340 153348
rect 191484 152046 191512 159938
rect 191760 153678 191788 160006
rect 192128 157282 192156 163200
rect 192116 157276 192168 157282
rect 192116 157218 192168 157224
rect 192956 155854 192984 163200
rect 193784 159186 193812 163200
rect 193680 159180 193732 159186
rect 193680 159122 193732 159128
rect 193772 159180 193824 159186
rect 193772 159122 193824 159128
rect 193692 158982 193720 159122
rect 193588 158976 193640 158982
rect 193588 158918 193640 158924
rect 193680 158976 193732 158982
rect 193680 158918 193732 158924
rect 193312 157616 193364 157622
rect 193312 157558 193364 157564
rect 193324 157334 193352 157558
rect 193324 157306 193536 157334
rect 192944 155848 192996 155854
rect 192944 155790 192996 155796
rect 192390 153776 192446 153785
rect 192390 153711 192446 153720
rect 191748 153672 191800 153678
rect 191748 153614 191800 153620
rect 191472 152040 191524 152046
rect 191472 151982 191524 151988
rect 190828 150204 190880 150210
rect 191116 150198 191190 150226
rect 190828 150146 190880 150152
rect 189184 150062 189258 150090
rect 189828 150062 189902 150090
rect 190472 150062 190546 150090
rect 189230 149940 189258 150062
rect 189874 149940 189902 150062
rect 190518 149940 190546 150062
rect 191162 149940 191190 150198
rect 191794 150204 191846 150210
rect 191794 150146 191846 150152
rect 191806 149940 191834 150146
rect 192404 150090 192432 153711
rect 193036 152924 193088 152930
rect 193036 152866 193088 152872
rect 193048 150090 193076 152866
rect 193508 150226 193536 157306
rect 193600 152182 193628 158918
rect 194704 158778 194732 163200
rect 195152 159316 195204 159322
rect 195152 159258 195204 159264
rect 195244 159316 195296 159322
rect 195244 159258 195296 159264
rect 195164 158914 195192 159258
rect 195256 159050 195284 159258
rect 195244 159044 195296 159050
rect 195244 158986 195296 158992
rect 195060 158908 195112 158914
rect 195060 158850 195112 158856
rect 195152 158908 195204 158914
rect 195152 158850 195204 158856
rect 194692 158772 194744 158778
rect 194692 158714 194744 158720
rect 194968 156324 195020 156330
rect 194968 156266 195020 156272
rect 194324 155916 194376 155922
rect 194324 155858 194376 155864
rect 193588 152176 193640 152182
rect 193588 152118 193640 152124
rect 193508 150198 193766 150226
rect 192404 150062 192478 150090
rect 193048 150062 193122 150090
rect 192450 149940 192478 150062
rect 193094 149940 193122 150062
rect 193738 149940 193766 150198
rect 194336 150090 194364 155858
rect 194980 150090 195008 156266
rect 195072 152998 195100 158850
rect 195532 157826 195560 163200
rect 195980 158840 196032 158846
rect 195980 158782 196032 158788
rect 195520 157820 195572 157826
rect 195520 157762 195572 157768
rect 195992 155106 196020 158782
rect 196256 156256 196308 156262
rect 196256 156198 196308 156204
rect 195980 155100 196032 155106
rect 195980 155042 196032 155048
rect 195888 153672 195940 153678
rect 195888 153614 195940 153620
rect 195980 153672 196032 153678
rect 195980 153614 196032 153620
rect 195900 153513 195928 153614
rect 195886 153504 195942 153513
rect 195886 153439 195942 153448
rect 195992 153270 196020 153614
rect 196070 153504 196126 153513
rect 196070 153439 196126 153448
rect 196084 153270 196112 153439
rect 195980 153264 196032 153270
rect 195980 153206 196032 153212
rect 196072 153264 196124 153270
rect 196072 153206 196124 153212
rect 195060 152992 195112 152998
rect 195060 152934 195112 152940
rect 195612 151972 195664 151978
rect 195612 151914 195664 151920
rect 195624 150090 195652 151914
rect 196268 150090 196296 156198
rect 196360 155922 196388 163200
rect 197188 160070 197216 163200
rect 197176 160064 197228 160070
rect 197176 160006 197228 160012
rect 198016 160002 198044 163200
rect 198004 159996 198056 160002
rect 198004 159938 198056 159944
rect 197360 158976 197412 158982
rect 197360 158918 197412 158924
rect 197372 157622 197400 158918
rect 198738 158536 198794 158545
rect 198738 158471 198794 158480
rect 197360 157616 197412 157622
rect 197360 157558 197412 157564
rect 197452 156256 197504 156262
rect 197452 156198 197504 156204
rect 197464 156058 197492 156198
rect 197452 156052 197504 156058
rect 197452 155994 197504 156000
rect 196348 155916 196400 155922
rect 196348 155858 196400 155864
rect 196992 155100 197044 155106
rect 196992 155042 197044 155048
rect 197004 153542 197032 155042
rect 196900 153536 196952 153542
rect 196900 153478 196952 153484
rect 196992 153536 197044 153542
rect 196992 153478 197044 153484
rect 196912 150090 196940 153478
rect 197544 153400 197596 153406
rect 197544 153342 197596 153348
rect 197556 150090 197584 153342
rect 198188 153060 198240 153066
rect 198188 153002 198240 153008
rect 198200 150090 198228 153002
rect 198752 150226 198780 158471
rect 198844 156398 198872 163200
rect 198924 158908 198976 158914
rect 198924 158850 198976 158856
rect 198832 156392 198884 156398
rect 198832 156334 198884 156340
rect 198936 153406 198964 158850
rect 199672 155106 199700 163200
rect 200592 158982 200620 163200
rect 201420 159322 201448 163200
rect 201316 159316 201368 159322
rect 201316 159258 201368 159264
rect 201408 159316 201460 159322
rect 201408 159258 201460 159264
rect 200580 158976 200632 158982
rect 200580 158918 200632 158924
rect 200764 156596 200816 156602
rect 200764 156538 200816 156544
rect 200948 156596 201000 156602
rect 200948 156538 201000 156544
rect 200776 156330 200804 156538
rect 200960 156398 200988 156538
rect 200948 156392 201000 156398
rect 200948 156334 201000 156340
rect 200764 156324 200816 156330
rect 200764 156266 200816 156272
rect 200672 156188 200724 156194
rect 200672 156130 200724 156136
rect 201040 156188 201092 156194
rect 201224 156188 201276 156194
rect 201092 156148 201224 156176
rect 201040 156130 201092 156136
rect 201224 156130 201276 156136
rect 200684 156074 200712 156130
rect 200684 156058 200988 156074
rect 200684 156052 201000 156058
rect 200684 156046 200948 156052
rect 200948 155994 201000 156000
rect 199660 155100 199712 155106
rect 199660 155042 199712 155048
rect 200120 155032 200172 155038
rect 200120 154974 200172 154980
rect 199476 153468 199528 153474
rect 199476 153410 199528 153416
rect 198924 153400 198976 153406
rect 198924 153342 198976 153348
rect 198752 150198 198918 150226
rect 194336 150062 194410 150090
rect 194980 150062 195054 150090
rect 195624 150062 195698 150090
rect 196268 150062 196342 150090
rect 196912 150062 196986 150090
rect 197556 150062 197630 150090
rect 198200 150062 198274 150090
rect 194382 149940 194410 150062
rect 195026 149940 195054 150062
rect 195670 149940 195698 150062
rect 196314 149940 196342 150062
rect 196958 149940 196986 150062
rect 197602 149940 197630 150062
rect 198246 149940 198274 150062
rect 198890 149940 198918 150198
rect 199488 150090 199516 153410
rect 200132 150090 200160 154974
rect 201328 154494 201356 159258
rect 202248 156058 202276 163200
rect 203076 156126 203104 163200
rect 203904 159050 203932 163200
rect 204732 159361 204760 163200
rect 204718 159352 204774 159361
rect 204718 159287 204774 159296
rect 204904 159112 204956 159118
rect 204904 159054 204956 159060
rect 203892 159044 203944 159050
rect 203892 158986 203944 158992
rect 203708 158772 203760 158778
rect 203708 158714 203760 158720
rect 203432 157548 203484 157554
rect 203432 157490 203484 157496
rect 203444 157334 203472 157490
rect 203444 157306 203656 157334
rect 203064 156120 203116 156126
rect 203064 156062 203116 156068
rect 201408 156052 201460 156058
rect 201408 155994 201460 156000
rect 202236 156052 202288 156058
rect 202236 155994 202288 156000
rect 201224 154488 201276 154494
rect 201224 154430 201276 154436
rect 201316 154488 201368 154494
rect 201316 154430 201368 154436
rect 201236 154358 201264 154430
rect 201132 154352 201184 154358
rect 201132 154294 201184 154300
rect 201224 154352 201276 154358
rect 201224 154294 201276 154300
rect 201144 153542 201172 154294
rect 200856 153536 200908 153542
rect 200856 153478 200908 153484
rect 201132 153536 201184 153542
rect 201132 153478 201184 153484
rect 200580 153400 200632 153406
rect 200764 153400 200816 153406
rect 200632 153348 200764 153354
rect 200580 153342 200816 153348
rect 200592 153326 200804 153342
rect 200868 153338 200896 153478
rect 200856 153332 200908 153338
rect 200856 153274 200908 153280
rect 200764 152108 200816 152114
rect 200764 152050 200816 152056
rect 200776 150090 200804 152050
rect 201420 150090 201448 155994
rect 202052 154420 202104 154426
rect 202052 154362 202104 154368
rect 202064 150090 202092 154362
rect 202696 154352 202748 154358
rect 202696 154294 202748 154300
rect 202708 150090 202736 154294
rect 203340 151904 203392 151910
rect 203340 151846 203392 151852
rect 203352 150090 203380 151846
rect 203628 150226 203656 157306
rect 203720 153066 203748 158714
rect 204916 157554 204944 159054
rect 204904 157548 204956 157554
rect 204904 157490 204956 157496
rect 204628 155780 204680 155786
rect 204628 155722 204680 155728
rect 203708 153060 203760 153066
rect 203708 153002 203760 153008
rect 203628 150198 204070 150226
rect 199488 150062 199562 150090
rect 200132 150062 200206 150090
rect 200776 150062 200850 150090
rect 201420 150062 201494 150090
rect 202064 150062 202138 150090
rect 202708 150062 202782 150090
rect 203352 150062 203426 150090
rect 199534 149940 199562 150062
rect 200178 149940 200206 150062
rect 200822 149940 200850 150062
rect 201466 149940 201494 150062
rect 202110 149940 202138 150062
rect 202754 149940 202782 150062
rect 203398 149940 203426 150062
rect 204042 149940 204070 150198
rect 204640 150090 204668 155722
rect 205008 154426 205036 163254
rect 205468 163146 205496 163254
rect 205546 163200 205602 164400
rect 206466 163200 206522 164400
rect 207294 163200 207350 164400
rect 208122 163200 208178 164400
rect 208412 163254 208900 163282
rect 205560 163146 205588 163200
rect 205468 163118 205588 163146
rect 206480 155786 206508 163200
rect 207020 160064 207072 160070
rect 207020 160006 207072 160012
rect 206560 157480 206612 157486
rect 206560 157422 206612 157428
rect 206468 155780 206520 155786
rect 206468 155722 206520 155728
rect 204996 154420 205048 154426
rect 204996 154362 205048 154368
rect 205272 153536 205324 153542
rect 205272 153478 205324 153484
rect 205364 153536 205416 153542
rect 205364 153478 205416 153484
rect 205284 150090 205312 153478
rect 205376 153406 205404 153478
rect 205364 153400 205416 153406
rect 205364 153342 205416 153348
rect 205916 153196 205968 153202
rect 205916 153138 205968 153144
rect 205928 150226 205956 153138
rect 206572 150226 206600 157422
rect 207032 155038 207060 160006
rect 207308 158846 207336 163200
rect 208136 158914 208164 163200
rect 208124 158908 208176 158914
rect 208124 158850 208176 158856
rect 207296 158840 207348 158846
rect 207296 158782 207348 158788
rect 207202 157176 207258 157185
rect 207202 157111 207258 157120
rect 207020 155032 207072 155038
rect 207020 154974 207072 154980
rect 207216 150226 207244 157111
rect 207940 154488 207992 154494
rect 207940 154430 207992 154436
rect 207952 153474 207980 154430
rect 208412 154358 208440 163254
rect 208872 163146 208900 163254
rect 208950 163200 209006 164400
rect 209778 163200 209834 164400
rect 210606 163200 210662 164400
rect 211434 163200 211490 164400
rect 211540 163254 212304 163282
rect 208964 163146 208992 163200
rect 208872 163118 208992 163146
rect 209792 156398 209820 163200
rect 210620 158778 210648 163200
rect 211448 160070 211476 163200
rect 211436 160064 211488 160070
rect 211436 160006 211488 160012
rect 210608 158772 210660 158778
rect 210608 158714 210660 158720
rect 209780 156392 209832 156398
rect 209780 156334 209832 156340
rect 209136 156188 209188 156194
rect 209136 156130 209188 156136
rect 208400 154352 208452 154358
rect 208400 154294 208452 154300
rect 207848 153468 207900 153474
rect 207848 153410 207900 153416
rect 207940 153468 207992 153474
rect 207940 153410 207992 153416
rect 207860 150226 207888 153410
rect 208492 152040 208544 152046
rect 208492 151982 208544 151988
rect 208504 150226 208532 151982
rect 209148 150226 209176 156130
rect 211252 154964 211304 154970
rect 211252 154906 211304 154912
rect 210424 153740 210476 153746
rect 210424 153682 210476 153688
rect 209780 153672 209832 153678
rect 209780 153614 209832 153620
rect 209792 150226 209820 153614
rect 210436 150226 210464 153682
rect 211068 152380 211120 152386
rect 211068 152322 211120 152328
rect 211080 150226 211108 152322
rect 205928 150198 206002 150226
rect 206572 150198 206646 150226
rect 207216 150198 207290 150226
rect 207860 150198 207934 150226
rect 208504 150198 208578 150226
rect 209148 150198 209222 150226
rect 209792 150198 209866 150226
rect 210436 150198 210510 150226
rect 211080 150198 211154 150226
rect 211264 150210 211292 154906
rect 211540 153785 211568 163254
rect 212276 163146 212304 163254
rect 212354 163200 212410 164400
rect 213182 163200 213238 164400
rect 214010 163200 214066 164400
rect 214838 163200 214894 164400
rect 215312 163254 215616 163282
rect 212368 163146 212396 163200
rect 212276 163118 212396 163146
rect 212632 159316 212684 159322
rect 212632 159258 212684 159264
rect 212448 158908 212500 158914
rect 212448 158850 212500 158856
rect 211620 156256 211672 156262
rect 211620 156198 211672 156204
rect 211526 153776 211582 153785
rect 211526 153711 211582 153720
rect 211632 150226 211660 156198
rect 212460 152930 212488 158850
rect 212448 152924 212500 152930
rect 212448 152866 212500 152872
rect 212644 151910 212672 159258
rect 213196 156330 213224 163200
rect 214024 159322 214052 163200
rect 214012 159316 214064 159322
rect 214012 159258 214064 159264
rect 214656 159248 214708 159254
rect 214656 159190 214708 159196
rect 213828 159044 213880 159050
rect 213828 158986 213880 158992
rect 213184 156324 213236 156330
rect 213184 156266 213236 156272
rect 212908 154556 212960 154562
rect 212908 154498 212960 154504
rect 212632 151904 212684 151910
rect 212632 151846 212684 151852
rect 212920 150226 212948 154498
rect 213552 152176 213604 152182
rect 213552 152118 213604 152124
rect 213564 150226 213592 152118
rect 213840 152114 213868 158986
rect 214472 157344 214524 157350
rect 214472 157286 214524 157292
rect 214564 157344 214616 157350
rect 214564 157286 214616 157292
rect 213920 156664 213972 156670
rect 213920 156606 213972 156612
rect 213828 152108 213880 152114
rect 213828 152050 213880 152056
rect 213932 151814 213960 156606
rect 214484 156262 214512 157286
rect 214576 156942 214604 157286
rect 214564 156936 214616 156942
rect 214564 156878 214616 156884
rect 214472 156256 214524 156262
rect 214472 156198 214524 156204
rect 214668 154970 214696 159190
rect 214852 159050 214880 163200
rect 214840 159044 214892 159050
rect 214840 158986 214892 158992
rect 214656 154964 214708 154970
rect 214656 154906 214708 154912
rect 214840 154828 214892 154834
rect 214840 154770 214892 154776
rect 213932 151786 214236 151814
rect 214208 150226 214236 151786
rect 214852 150226 214880 154770
rect 215312 154494 215340 163254
rect 215588 163146 215616 163254
rect 215666 163200 215722 164400
rect 216494 163200 216550 164400
rect 217322 163200 217378 164400
rect 218242 163200 218298 164400
rect 218348 163254 219020 163282
rect 215680 163146 215708 163200
rect 215588 163118 215708 163146
rect 215392 158772 215444 158778
rect 215392 158714 215444 158720
rect 215300 154488 215352 154494
rect 215300 154430 215352 154436
rect 215404 153202 215432 158714
rect 216508 156670 216536 163200
rect 217336 158846 217364 163200
rect 218256 159254 218284 163200
rect 218244 159248 218296 159254
rect 218244 159190 218296 159196
rect 218060 159180 218112 159186
rect 218060 159122 218112 159128
rect 217324 158840 217376 158846
rect 217324 158782 217376 158788
rect 216772 156732 216824 156738
rect 216772 156674 216824 156680
rect 216496 156664 216548 156670
rect 216496 156606 216548 156612
rect 215484 156188 215536 156194
rect 215484 156130 215536 156136
rect 215392 153196 215444 153202
rect 215392 153138 215444 153144
rect 215496 150226 215524 156130
rect 216128 152516 216180 152522
rect 216128 152458 216180 152464
rect 216140 150226 216168 152458
rect 216784 150226 216812 156674
rect 218072 156194 218100 159122
rect 218060 156188 218112 156194
rect 218060 156130 218112 156136
rect 217416 155236 217468 155242
rect 217416 155178 217468 155184
rect 217428 150226 217456 155178
rect 218348 154562 218376 163254
rect 218992 163146 219020 163254
rect 219070 163200 219126 164400
rect 219898 163200 219954 164400
rect 220726 163200 220782 164400
rect 221554 163200 221610 164400
rect 222382 163200 222438 164400
rect 223210 163200 223266 164400
rect 224130 163200 224186 164400
rect 224958 163200 225014 164400
rect 225248 163254 225736 163282
rect 219084 163146 219112 163200
rect 218992 163118 219112 163146
rect 219912 161474 219940 163200
rect 219912 161446 220124 161474
rect 219348 158024 219400 158030
rect 219348 157966 219400 157972
rect 218336 154556 218388 154562
rect 218336 154498 218388 154504
rect 218060 153808 218112 153814
rect 218060 153750 218112 153756
rect 218072 150226 218100 153750
rect 218704 152992 218756 152998
rect 218704 152934 218756 152940
rect 218716 150226 218744 152934
rect 219360 150226 219388 157966
rect 220096 156262 220124 161446
rect 220740 159118 220768 163200
rect 220728 159112 220780 159118
rect 220728 159054 220780 159060
rect 220360 158840 220412 158846
rect 220360 158782 220412 158788
rect 219992 156256 220044 156262
rect 219992 156198 220044 156204
rect 220084 156256 220136 156262
rect 220084 156198 220136 156204
rect 219900 154012 219952 154018
rect 219900 153954 219952 153960
rect 204640 150062 204714 150090
rect 205284 150062 205358 150090
rect 204686 149940 204714 150062
rect 205330 149940 205358 150062
rect 205974 149940 206002 150198
rect 206618 149940 206646 150198
rect 207262 149940 207290 150198
rect 207906 149940 207934 150198
rect 208550 149940 208578 150198
rect 209194 149940 209222 150198
rect 209838 149940 209866 150198
rect 210482 149940 210510 150198
rect 211126 149940 211154 150198
rect 211252 150204 211304 150210
rect 211632 150198 211706 150226
rect 211252 150146 211304 150152
rect 211678 149940 211706 150198
rect 212310 150204 212362 150210
rect 212920 150198 212994 150226
rect 213564 150198 213638 150226
rect 214208 150198 214282 150226
rect 214852 150198 214926 150226
rect 215496 150198 215570 150226
rect 216140 150198 216214 150226
rect 216784 150198 216858 150226
rect 217428 150198 217502 150226
rect 218072 150198 218146 150226
rect 218716 150198 218790 150226
rect 219360 150198 219434 150226
rect 212310 150146 212362 150152
rect 212322 149940 212350 150146
rect 212966 149940 212994 150198
rect 213610 149940 213638 150198
rect 214254 149940 214282 150198
rect 214898 149940 214926 150198
rect 215542 149940 215570 150198
rect 216186 149940 216214 150198
rect 216830 149940 216858 150198
rect 217474 149940 217502 150198
rect 218118 149940 218146 150198
rect 218762 149940 218790 150198
rect 219406 149940 219434 150198
rect 219912 150192 219940 153954
rect 220004 151814 220032 156198
rect 220372 152998 220400 158782
rect 221568 158778 221596 163200
rect 222108 159044 222160 159050
rect 222108 158986 222160 158992
rect 221556 158772 221608 158778
rect 221556 158714 221608 158720
rect 221372 157344 221424 157350
rect 221372 157286 221424 157292
rect 220360 152992 220412 152998
rect 220360 152934 220412 152940
rect 221280 152244 221332 152250
rect 221280 152186 221332 152192
rect 220004 151786 220676 151814
rect 220648 150226 220676 151786
rect 221292 150226 221320 152186
rect 221384 151814 221412 157286
rect 222120 152250 222148 158986
rect 222396 154018 222424 163200
rect 222568 156800 222620 156806
rect 222568 156742 222620 156748
rect 222384 154012 222436 154018
rect 222384 153954 222436 153960
rect 222108 152244 222160 152250
rect 222108 152186 222160 152192
rect 221384 151786 221964 151814
rect 221936 150226 221964 151786
rect 222580 150226 222608 156742
rect 223224 156738 223252 163200
rect 223580 159384 223632 159390
rect 223580 159326 223632 159332
rect 223212 156732 223264 156738
rect 223212 156674 223264 156680
rect 223212 153944 223264 153950
rect 223212 153886 223264 153892
rect 223224 150226 223252 153886
rect 223592 151814 223620 159326
rect 224144 159050 224172 163200
rect 224972 159186 225000 163200
rect 224960 159180 225012 159186
rect 224960 159122 225012 159128
rect 224132 159044 224184 159050
rect 224132 158986 224184 158992
rect 224960 158976 225012 158982
rect 224960 158918 225012 158924
rect 224408 158772 224460 158778
rect 224408 158714 224460 158720
rect 224224 157344 224276 157350
rect 224224 157286 224276 157292
rect 224132 157004 224184 157010
rect 224132 156946 224184 156952
rect 224144 151814 224172 156946
rect 224236 156330 224264 157286
rect 224224 156324 224276 156330
rect 224224 156266 224276 156272
rect 224420 152386 224448 158714
rect 224972 156942 225000 158918
rect 224960 156936 225012 156942
rect 224960 156878 225012 156884
rect 225144 156868 225196 156874
rect 225144 156810 225196 156816
rect 225052 156528 225104 156534
rect 225052 156470 225104 156476
rect 224408 152380 224460 152386
rect 224408 152322 224460 152328
rect 223592 151786 223896 151814
rect 224144 151786 224540 151814
rect 223868 150226 223896 151786
rect 224512 150226 224540 151786
rect 220648 150198 220722 150226
rect 221292 150198 221366 150226
rect 221936 150198 222010 150226
rect 222580 150198 222654 150226
rect 223224 150198 223298 150226
rect 223868 150198 223942 150226
rect 224512 150198 224586 150226
rect 225064 150210 225092 156470
rect 225156 150226 225184 156810
rect 225248 153950 225276 163254
rect 225708 163146 225736 163254
rect 225786 163200 225842 164400
rect 226614 163200 226670 164400
rect 227442 163200 227498 164400
rect 227732 163254 228220 163282
rect 225800 163146 225828 163200
rect 225708 163118 225828 163146
rect 225328 159520 225380 159526
rect 225328 159462 225380 159468
rect 225236 153944 225288 153950
rect 225236 153886 225288 153892
rect 225340 152182 225368 159462
rect 226628 156874 226656 163200
rect 227076 157412 227128 157418
rect 227076 157354 227128 157360
rect 226616 156868 226668 156874
rect 226616 156810 226668 156816
rect 226432 152584 226484 152590
rect 226432 152526 226484 152532
rect 225328 152176 225380 152182
rect 225328 152118 225380 152124
rect 226444 150226 226472 152526
rect 227088 150226 227116 157354
rect 227456 152425 227484 163200
rect 227732 152522 227760 163254
rect 228192 163146 228220 163254
rect 228270 163200 228326 164400
rect 229098 163200 229154 164400
rect 230018 163200 230074 164400
rect 230846 163200 230902 164400
rect 231674 163200 231730 164400
rect 231872 163254 232452 163282
rect 228284 163146 228312 163200
rect 228192 163118 228312 163146
rect 228364 156460 228416 156466
rect 228364 156402 228416 156408
rect 227812 155304 227864 155310
rect 227812 155246 227864 155252
rect 227720 152516 227772 152522
rect 227720 152458 227772 152464
rect 227442 152416 227498 152425
rect 227442 152351 227498 152360
rect 227824 150226 227852 155246
rect 219912 150164 220078 150192
rect 220050 149940 220078 150164
rect 220694 149940 220722 150198
rect 221338 149940 221366 150198
rect 221982 149940 222010 150198
rect 222626 149940 222654 150198
rect 223270 149940 223298 150198
rect 223914 149940 223942 150198
rect 224558 149940 224586 150198
rect 225052 150204 225104 150210
rect 225156 150198 225230 150226
rect 225052 150146 225104 150152
rect 225202 149940 225230 150198
rect 225834 150204 225886 150210
rect 226444 150198 226518 150226
rect 227088 150198 227162 150226
rect 225834 150146 225886 150152
rect 225846 149940 225874 150146
rect 226490 149940 226518 150198
rect 227134 149940 227162 150198
rect 227778 150198 227852 150226
rect 228376 150226 228404 156402
rect 229112 153678 229140 163200
rect 230032 156806 230060 163200
rect 230860 159526 230888 163200
rect 230848 159520 230900 159526
rect 230848 159462 230900 159468
rect 231688 159390 231716 163200
rect 231676 159384 231728 159390
rect 231676 159326 231728 159332
rect 230756 158908 230808 158914
rect 230756 158850 230808 158856
rect 230020 156800 230072 156806
rect 230020 156742 230072 156748
rect 230768 156194 230796 158850
rect 230756 156188 230808 156194
rect 230756 156130 230808 156136
rect 229652 155984 229704 155990
rect 229652 155926 229704 155932
rect 229192 155372 229244 155378
rect 229192 155314 229244 155320
rect 229100 153672 229152 153678
rect 229100 153614 229152 153620
rect 229008 152176 229060 152182
rect 229008 152118 229060 152124
rect 229020 150226 229048 152118
rect 228376 150198 228450 150226
rect 229020 150198 229094 150226
rect 229204 150210 229232 155314
rect 229664 150226 229692 155926
rect 231872 153814 231900 163254
rect 232424 163146 232452 163254
rect 232502 163200 232558 164400
rect 233330 163200 233386 164400
rect 234158 163200 234214 164400
rect 234986 163200 235042 164400
rect 235092 163254 235856 163282
rect 232516 163146 232544 163200
rect 232424 163118 232544 163146
rect 233240 159452 233292 159458
rect 233240 159394 233292 159400
rect 231952 158092 232004 158098
rect 231952 158034 232004 158040
rect 231860 153808 231912 153814
rect 231860 153750 231912 153756
rect 230940 153604 230992 153610
rect 230940 153546 230992 153552
rect 230952 150226 230980 153546
rect 231584 152720 231636 152726
rect 231584 152662 231636 152668
rect 231596 150226 231624 152662
rect 231964 151814 231992 158034
rect 232872 155440 232924 155446
rect 232872 155382 232924 155388
rect 231964 151786 232268 151814
rect 232240 150226 232268 151786
rect 232884 150226 232912 155382
rect 227778 149940 227806 150198
rect 228422 149940 228450 150198
rect 229066 149940 229094 150198
rect 229192 150204 229244 150210
rect 229664 150198 229738 150226
rect 229192 150146 229244 150152
rect 229710 149940 229738 150198
rect 230342 150204 230394 150210
rect 230952 150198 231026 150226
rect 231596 150198 231670 150226
rect 232240 150198 232314 150226
rect 232884 150198 232958 150226
rect 233252 150210 233280 159394
rect 233344 155310 233372 163200
rect 233516 157140 233568 157146
rect 233516 157082 233568 157088
rect 233332 155304 233384 155310
rect 233332 155246 233384 155252
rect 233528 150226 233556 157082
rect 234172 152590 234200 163200
rect 235000 159458 235028 163200
rect 234988 159452 235040 159458
rect 234988 159394 235040 159400
rect 234804 157072 234856 157078
rect 234804 157014 234856 157020
rect 234160 152584 234212 152590
rect 234160 152526 234212 152532
rect 234816 150226 234844 157014
rect 235092 153746 235120 163254
rect 235828 163146 235856 163254
rect 235906 163200 235962 164400
rect 236734 163200 236790 164400
rect 237562 163200 237618 164400
rect 238390 163200 238446 164400
rect 238864 163254 239168 163282
rect 235920 163146 235948 163200
rect 235828 163118 235948 163146
rect 236748 158030 236776 163200
rect 237576 158982 237604 163200
rect 237564 158976 237616 158982
rect 237564 158918 237616 158924
rect 238404 158846 238432 163200
rect 238392 158840 238444 158846
rect 238392 158782 238444 158788
rect 237380 158228 237432 158234
rect 237380 158170 237432 158176
rect 236736 158024 236788 158030
rect 236736 157966 236788 157972
rect 236092 157684 236144 157690
rect 236092 157626 236144 157632
rect 235448 153876 235500 153882
rect 235448 153818 235500 153824
rect 235080 153740 235132 153746
rect 235080 153682 235132 153688
rect 235460 150226 235488 153818
rect 236104 150226 236132 157626
rect 236736 152652 236788 152658
rect 236736 152594 236788 152600
rect 236748 150226 236776 152594
rect 237392 150226 237420 158170
rect 238024 154760 238076 154766
rect 238024 154702 238076 154708
rect 238036 150226 238064 154702
rect 238864 153610 238892 163254
rect 239140 163146 239168 163254
rect 239218 163200 239274 164400
rect 240046 163200 240102 164400
rect 240874 163200 240930 164400
rect 241794 163200 241850 164400
rect 241900 163254 242572 163282
rect 239232 163146 239260 163200
rect 239140 163118 239260 163146
rect 239312 159588 239364 159594
rect 239312 159530 239364 159536
rect 238944 158160 238996 158166
rect 238944 158102 238996 158108
rect 238852 153604 238904 153610
rect 238852 153546 238904 153552
rect 238668 153332 238720 153338
rect 238668 153274 238720 153280
rect 238680 150226 238708 153274
rect 230342 150146 230394 150152
rect 230354 149940 230382 150146
rect 230998 149940 231026 150198
rect 231642 149940 231670 150198
rect 232286 149940 232314 150198
rect 232930 149940 232958 150198
rect 233240 150204 233292 150210
rect 233528 150198 233602 150226
rect 233240 150146 233292 150152
rect 233574 149940 233602 150198
rect 234206 150204 234258 150210
rect 234816 150198 234890 150226
rect 235460 150198 235534 150226
rect 236104 150198 236178 150226
rect 236748 150198 236822 150226
rect 237392 150198 237466 150226
rect 238036 150198 238110 150226
rect 238680 150198 238754 150226
rect 238956 150210 238984 158102
rect 239324 150226 239352 159530
rect 240060 155242 240088 163200
rect 240324 159656 240376 159662
rect 240324 159598 240376 159604
rect 240048 155236 240100 155242
rect 240048 155178 240100 155184
rect 240336 152726 240364 159598
rect 240888 158778 240916 163200
rect 241808 158914 241836 163200
rect 241796 158908 241848 158914
rect 241796 158850 241848 158856
rect 240876 158772 240928 158778
rect 240876 158714 240928 158720
rect 240600 154624 240652 154630
rect 240600 154566 240652 154572
rect 240324 152720 240376 152726
rect 240324 152662 240376 152668
rect 240612 150226 240640 154566
rect 241244 154080 241296 154086
rect 241244 154022 241296 154028
rect 241256 150226 241284 154022
rect 241900 153882 241928 163254
rect 242544 163146 242572 163254
rect 242622 163200 242678 164400
rect 243450 163200 243506 164400
rect 244278 163200 244334 164400
rect 244476 163254 245056 163282
rect 242636 163146 242664 163200
rect 242544 163118 242664 163146
rect 242440 158840 242492 158846
rect 242440 158782 242492 158788
rect 242072 158296 242124 158302
rect 242072 158238 242124 158244
rect 241888 153876 241940 153882
rect 241888 153818 241940 153824
rect 241888 152720 241940 152726
rect 241888 152662 241940 152668
rect 241900 150226 241928 152662
rect 242084 151814 242112 158238
rect 242452 152046 242480 158782
rect 243360 158772 243412 158778
rect 243360 158714 243412 158720
rect 243084 154692 243136 154698
rect 243084 154634 243136 154640
rect 242440 152040 242492 152046
rect 242440 151982 242492 151988
rect 242084 151786 242480 151814
rect 242452 150226 242480 151786
rect 243096 150226 243124 154634
rect 243372 151978 243400 158714
rect 243464 158098 243492 163200
rect 244292 159662 244320 163200
rect 244280 159656 244332 159662
rect 244280 159598 244332 159604
rect 243452 158092 243504 158098
rect 243452 158034 243504 158040
rect 243728 153400 243780 153406
rect 243728 153342 243780 153348
rect 243360 151972 243412 151978
rect 243360 151914 243412 151920
rect 243740 150226 243768 153342
rect 244372 152788 244424 152794
rect 244372 152730 244424 152736
rect 244384 150226 244412 152730
rect 244476 152182 244504 163254
rect 245028 163146 245056 163254
rect 245106 163200 245162 164400
rect 245934 163200 245990 164400
rect 246762 163200 246818 164400
rect 247052 163254 247632 163282
rect 245120 163146 245148 163200
rect 245028 163118 245148 163146
rect 245016 158432 245068 158438
rect 245016 158374 245068 158380
rect 244464 152176 244516 152182
rect 244464 152118 244516 152124
rect 245028 150226 245056 158374
rect 245844 154896 245896 154902
rect 245844 154838 245896 154844
rect 245660 154148 245712 154154
rect 245660 154090 245712 154096
rect 245672 150226 245700 154090
rect 245856 151814 245884 154838
rect 245948 154154 245976 163200
rect 246776 158166 246804 163200
rect 246948 159724 247000 159730
rect 246948 159666 247000 159672
rect 246764 158160 246816 158166
rect 246764 158102 246816 158108
rect 245936 154148 245988 154154
rect 245936 154090 245988 154096
rect 245856 151786 246344 151814
rect 246316 150226 246344 151786
rect 246960 150226 246988 159666
rect 247052 152658 247080 163254
rect 247604 163146 247632 163254
rect 247682 163200 247738 164400
rect 248510 163200 248566 164400
rect 248616 163254 249288 163282
rect 247696 163146 247724 163200
rect 247604 163118 247724 163146
rect 248524 159730 248552 163200
rect 248512 159724 248564 159730
rect 248512 159666 248564 159672
rect 247132 158364 247184 158370
rect 247132 158306 247184 158312
rect 247040 152652 247092 152658
rect 247040 152594 247092 152600
rect 247144 151814 247172 158306
rect 248236 155508 248288 155514
rect 248236 155450 248288 155456
rect 247144 151786 247632 151814
rect 247604 150226 247632 151786
rect 248248 150226 248276 155450
rect 248616 154086 248644 163254
rect 249260 163146 249288 163254
rect 249338 163200 249394 164400
rect 250166 163200 250222 164400
rect 250994 163200 251050 164400
rect 251192 163254 251772 163282
rect 249352 163146 249380 163200
rect 249260 163118 249380 163146
rect 250076 158636 250128 158642
rect 250076 158578 250128 158584
rect 248604 154080 248656 154086
rect 248604 154022 248656 154028
rect 248880 153536 248932 153542
rect 248880 153478 248932 153484
rect 248892 150226 248920 153478
rect 249524 152448 249576 152454
rect 249524 152390 249576 152396
rect 249536 150226 249564 152390
rect 250088 151814 250116 158578
rect 250180 155378 250208 163200
rect 251008 159594 251036 163200
rect 250996 159588 251048 159594
rect 250996 159530 251048 159536
rect 250168 155372 250220 155378
rect 250168 155314 250220 155320
rect 250812 154216 250864 154222
rect 250812 154158 250864 154164
rect 250088 151786 250208 151814
rect 250180 150226 250208 151786
rect 250824 150226 250852 154158
rect 251192 152726 251220 163254
rect 251744 163146 251772 163254
rect 251822 163200 251878 164400
rect 252650 163200 252706 164400
rect 253570 163200 253626 164400
rect 254398 163200 254454 164400
rect 255226 163200 255282 164400
rect 255332 163254 256004 163282
rect 251836 163146 251864 163200
rect 251744 163118 251864 163146
rect 251456 157616 251508 157622
rect 251456 157558 251508 157564
rect 251180 152720 251232 152726
rect 251180 152662 251232 152668
rect 251468 150226 251496 157558
rect 252664 153542 252692 163200
rect 252744 158568 252796 158574
rect 252744 158510 252796 158516
rect 252652 153536 252704 153542
rect 252652 153478 252704 153484
rect 252100 152856 252152 152862
rect 252100 152798 252152 152804
rect 252112 150226 252140 152798
rect 252756 150226 252784 158510
rect 253388 155644 253440 155650
rect 253388 155586 253440 155592
rect 253400 150226 253428 155586
rect 253584 155446 253612 163200
rect 253940 159792 253992 159798
rect 253940 159734 253992 159740
rect 253572 155440 253624 155446
rect 253572 155382 253624 155388
rect 234206 150146 234258 150152
rect 234218 149940 234246 150146
rect 234862 149940 234890 150198
rect 235506 149940 235534 150198
rect 236150 149940 236178 150198
rect 236794 149940 236822 150198
rect 237438 149940 237466 150198
rect 238082 149940 238110 150198
rect 238726 149940 238754 150198
rect 238944 150204 238996 150210
rect 239324 150198 239398 150226
rect 238944 150146 238996 150152
rect 239370 149940 239398 150198
rect 240002 150204 240054 150210
rect 240612 150198 240686 150226
rect 241256 150198 241330 150226
rect 241900 150198 241974 150226
rect 242452 150198 242526 150226
rect 243096 150198 243170 150226
rect 243740 150198 243814 150226
rect 244384 150198 244458 150226
rect 245028 150198 245102 150226
rect 245672 150198 245746 150226
rect 246316 150198 246390 150226
rect 246960 150198 247034 150226
rect 247604 150198 247678 150226
rect 248248 150198 248322 150226
rect 248892 150198 248966 150226
rect 249536 150198 249610 150226
rect 250180 150198 250254 150226
rect 250824 150198 250898 150226
rect 251468 150198 251542 150226
rect 252112 150198 252186 150226
rect 252756 150198 252830 150226
rect 253400 150198 253474 150226
rect 253952 150210 253980 159734
rect 254412 158778 254440 163200
rect 255240 159798 255268 163200
rect 255228 159792 255280 159798
rect 255228 159734 255280 159740
rect 254400 158772 254452 158778
rect 254400 158714 254452 158720
rect 254032 157208 254084 157214
rect 254032 157150 254084 157156
rect 254044 150226 254072 157150
rect 255332 154222 255360 163254
rect 255976 163146 256004 163254
rect 256054 163200 256110 164400
rect 256882 163200 256938 164400
rect 257710 163200 257766 164400
rect 258538 163200 258594 164400
rect 259458 163200 259514 164400
rect 260286 163200 260342 164400
rect 261114 163200 261170 164400
rect 261942 163200 261998 164400
rect 262232 163254 262720 163282
rect 256068 163146 256096 163200
rect 255976 163118 256096 163146
rect 255412 158772 255464 158778
rect 255412 158714 255464 158720
rect 255320 154216 255372 154222
rect 255320 154158 255372 154164
rect 255424 152862 255452 158714
rect 256792 158704 256844 158710
rect 256792 158646 256844 158652
rect 255596 158500 255648 158506
rect 255596 158442 255648 158448
rect 255412 152856 255464 152862
rect 255412 152798 255464 152804
rect 255608 152538 255636 158442
rect 255872 157548 255924 157554
rect 255872 157490 255924 157496
rect 255688 155576 255740 155582
rect 255688 155518 255740 155524
rect 255424 152510 255636 152538
rect 255424 150226 255452 152510
rect 255700 151814 255728 155518
rect 255884 151814 255912 157490
rect 255700 151786 255820 151814
rect 255884 151786 256648 151814
rect 240002 150146 240054 150152
rect 240014 149940 240042 150146
rect 240658 149940 240686 150198
rect 241302 149940 241330 150198
rect 241946 149940 241974 150198
rect 242498 149940 242526 150198
rect 243142 149940 243170 150198
rect 243786 149940 243814 150198
rect 244430 149940 244458 150198
rect 245074 149940 245102 150198
rect 245718 149940 245746 150198
rect 246362 149940 246390 150198
rect 247006 149940 247034 150198
rect 247650 149940 247678 150198
rect 248294 149940 248322 150198
rect 248938 149940 248966 150198
rect 249582 149940 249610 150198
rect 250226 149940 250254 150198
rect 250870 149940 250898 150198
rect 251514 149940 251542 150198
rect 252158 149940 252186 150198
rect 252802 149940 252830 150198
rect 253446 149940 253474 150198
rect 253940 150204 253992 150210
rect 254044 150198 254118 150226
rect 253940 150146 253992 150152
rect 254090 149940 254118 150198
rect 254722 150204 254774 150210
rect 254722 150146 254774 150152
rect 255378 150198 255452 150226
rect 255792 150226 255820 151786
rect 256620 150226 256648 151786
rect 255792 150198 256050 150226
rect 256620 150198 256694 150226
rect 256804 150210 256832 158646
rect 256896 158234 256924 163200
rect 256884 158228 256936 158234
rect 256884 158170 256936 158176
rect 257252 153128 257304 153134
rect 257252 153070 257304 153076
rect 257264 150226 257292 153070
rect 257724 152794 257752 163200
rect 258552 158778 258580 163200
rect 258540 158772 258592 158778
rect 258540 158714 258592 158720
rect 258540 154284 258592 154290
rect 258540 154226 258592 154232
rect 257712 152788 257764 152794
rect 257712 152730 257764 152736
rect 258552 150226 258580 154226
rect 259184 153468 259236 153474
rect 259184 153410 259236 153416
rect 259196 150226 259224 153410
rect 259472 153406 259500 163200
rect 259552 159860 259604 159866
rect 259552 159802 259604 159808
rect 259460 153400 259512 153406
rect 259460 153342 259512 153348
rect 259564 151814 259592 159802
rect 260300 155514 260328 163200
rect 261128 158846 261156 163200
rect 261956 159866 261984 163200
rect 261944 159860 261996 159866
rect 261944 159802 261996 159808
rect 261116 158840 261168 158846
rect 261116 158782 261168 158788
rect 260932 158772 260984 158778
rect 260932 158714 260984 158720
rect 260472 157956 260524 157962
rect 260472 157898 260524 157904
rect 260288 155508 260340 155514
rect 260288 155450 260340 155456
rect 259564 151786 259868 151814
rect 259840 150226 259868 151786
rect 260484 150226 260512 157898
rect 260840 155712 260892 155718
rect 260840 155654 260892 155660
rect 260852 151814 260880 155654
rect 260944 152454 260972 158714
rect 261392 154964 261444 154970
rect 261392 154906 261444 154912
rect 260932 152448 260984 152454
rect 260932 152390 260984 152396
rect 261404 151814 261432 154906
rect 262232 154290 262260 163254
rect 262692 163146 262720 163254
rect 262770 163200 262826 164400
rect 263598 163200 263654 164400
rect 264426 163200 264482 164400
rect 264992 163254 265296 163282
rect 262784 163146 262812 163200
rect 262692 163118 262812 163146
rect 263048 157888 263100 157894
rect 263048 157830 263100 157836
rect 262220 154284 262272 154290
rect 262220 154226 262272 154232
rect 262404 152312 262456 152318
rect 262404 152254 262456 152260
rect 260852 151786 261156 151814
rect 261404 151786 261800 151814
rect 261128 150226 261156 151786
rect 261772 150226 261800 151786
rect 262416 150226 262444 152254
rect 263060 150226 263088 157830
rect 263612 155582 263640 163200
rect 264440 158778 264468 163200
rect 264888 159928 264940 159934
rect 264888 159870 264940 159876
rect 264428 158772 264480 158778
rect 264428 158714 264480 158720
rect 263692 157752 263744 157758
rect 263692 157694 263744 157700
rect 263600 155576 263652 155582
rect 263600 155518 263652 155524
rect 263704 155394 263732 157694
rect 263612 155366 263732 155394
rect 254734 149940 254762 150146
rect 255378 149940 255406 150198
rect 256022 149940 256050 150198
rect 256666 149940 256694 150198
rect 256792 150204 256844 150210
rect 257264 150198 257338 150226
rect 256792 150146 256844 150152
rect 257310 149940 257338 150198
rect 257942 150204 257994 150210
rect 258552 150198 258626 150226
rect 259196 150198 259270 150226
rect 259840 150198 259914 150226
rect 260484 150198 260558 150226
rect 261128 150198 261202 150226
rect 261772 150198 261846 150226
rect 262416 150198 262490 150226
rect 263060 150198 263134 150226
rect 263612 150210 263640 155366
rect 263692 155168 263744 155174
rect 263692 155110 263744 155116
rect 263704 150226 263732 155110
rect 264900 151814 264928 159870
rect 264992 153134 265020 163254
rect 265268 163146 265296 163254
rect 265346 163200 265402 164400
rect 265452 163254 266124 163282
rect 265360 163146 265388 163200
rect 265268 163118 265388 163146
rect 265164 157276 265216 157282
rect 265164 157218 265216 157224
rect 264980 153128 265032 153134
rect 264980 153070 265032 153076
rect 265176 151814 265204 157218
rect 265452 153474 265480 163254
rect 266096 163146 266124 163254
rect 266174 163200 266230 164400
rect 267002 163200 267058 164400
rect 267830 163200 267886 164400
rect 268658 163200 268714 164400
rect 269224 163254 269436 163282
rect 266188 163146 266216 163200
rect 266096 163118 266216 163146
rect 266360 158772 266412 158778
rect 266360 158714 266412 158720
rect 266268 155848 266320 155854
rect 266268 155790 266320 155796
rect 265440 153468 265492 153474
rect 265440 153410 265492 153416
rect 264900 151786 265020 151814
rect 265176 151786 265664 151814
rect 264992 150226 265020 151786
rect 265636 150226 265664 151786
rect 266280 150226 266308 155790
rect 266372 152318 266400 158714
rect 266912 156256 266964 156262
rect 266912 156198 266964 156204
rect 266360 152312 266412 152318
rect 266360 152254 266412 152260
rect 266924 150226 266952 156198
rect 267016 155650 267044 163200
rect 267844 158778 267872 163200
rect 268672 159934 268700 163200
rect 269120 159996 269172 160002
rect 269120 159938 269172 159944
rect 268660 159928 268712 159934
rect 268660 159870 268712 159876
rect 267832 158772 267884 158778
rect 267832 158714 267884 158720
rect 267740 157820 267792 157826
rect 267740 157762 267792 157768
rect 267004 155644 267056 155650
rect 267004 155586 267056 155592
rect 267556 153060 267608 153066
rect 267556 153002 267608 153008
rect 267568 150226 267596 153002
rect 267752 151814 267780 157762
rect 268844 155916 268896 155922
rect 268844 155858 268896 155864
rect 267752 151786 268240 151814
rect 268212 150226 268240 151786
rect 268856 150226 268884 155858
rect 257942 150146 257994 150152
rect 257954 149940 257982 150146
rect 258598 149940 258626 150198
rect 259242 149940 259270 150198
rect 259886 149940 259914 150198
rect 260530 149940 260558 150198
rect 261174 149940 261202 150198
rect 261818 149940 261846 150198
rect 262462 149940 262490 150198
rect 263106 149940 263134 150198
rect 263600 150204 263652 150210
rect 263704 150198 263778 150226
rect 263600 150146 263652 150152
rect 263750 149940 263778 150198
rect 264382 150204 264434 150210
rect 264992 150198 265066 150226
rect 265636 150198 265710 150226
rect 266280 150198 266354 150226
rect 266924 150198 266998 150226
rect 267568 150198 267642 150226
rect 268212 150198 268286 150226
rect 268856 150198 268930 150226
rect 269132 150210 269160 159938
rect 269224 153270 269252 163254
rect 269408 163146 269436 163254
rect 269486 163200 269542 164400
rect 270314 163200 270370 164400
rect 271234 163200 271290 164400
rect 272062 163200 272118 164400
rect 272890 163200 272946 164400
rect 273718 163200 273774 164400
rect 274546 163200 274602 164400
rect 275374 163200 275430 164400
rect 276202 163200 276258 164400
rect 277122 163200 277178 164400
rect 277412 163254 277900 163282
rect 269500 163146 269528 163200
rect 269408 163118 269528 163146
rect 270328 155718 270356 163200
rect 271248 160002 271276 163200
rect 272076 161474 272104 163200
rect 272076 161446 272196 161474
rect 271236 159996 271288 160002
rect 271236 159938 271288 159944
rect 271880 159996 271932 160002
rect 271880 159938 271932 159944
rect 270500 156596 270552 156602
rect 270500 156538 270552 156544
rect 270316 155712 270368 155718
rect 270316 155654 270368 155660
rect 269488 155032 269540 155038
rect 269488 154974 269540 154980
rect 269212 153264 269264 153270
rect 269212 153206 269264 153212
rect 269500 150226 269528 154974
rect 270512 151814 270540 156538
rect 271420 155100 271472 155106
rect 271420 155042 271472 155048
rect 270512 151786 270816 151814
rect 270788 150226 270816 151786
rect 271432 150226 271460 155042
rect 271892 151842 271920 159938
rect 272064 156936 272116 156942
rect 272064 156878 272116 156884
rect 271880 151836 271932 151842
rect 271880 151778 271932 151784
rect 272076 150226 272104 156878
rect 272168 153066 272196 161446
rect 272904 153338 272932 163200
rect 273732 157010 273760 163200
rect 274560 159497 274588 163200
rect 275388 160002 275416 163200
rect 275376 159996 275428 160002
rect 275376 159938 275428 159944
rect 274546 159488 274602 159497
rect 274546 159423 274602 159432
rect 275190 159352 275246 159361
rect 275190 159287 275246 159296
rect 273720 157004 273772 157010
rect 273720 156946 273772 156952
rect 273904 156120 273956 156126
rect 273904 156062 273956 156068
rect 273260 156052 273312 156058
rect 273260 155994 273312 156000
rect 272892 153332 272944 153338
rect 272892 153274 272944 153280
rect 272156 153060 272208 153066
rect 272156 153002 272208 153008
rect 272708 151904 272760 151910
rect 272708 151846 272760 151852
rect 272720 150226 272748 151846
rect 273272 150226 273300 155994
rect 273916 150226 273944 156062
rect 274548 152108 274600 152114
rect 274548 152050 274600 152056
rect 274560 150226 274588 152050
rect 275204 150226 275232 159287
rect 276112 155780 276164 155786
rect 276112 155722 276164 155728
rect 275836 154420 275888 154426
rect 275836 154362 275888 154368
rect 275848 150226 275876 154362
rect 276124 151814 276152 155722
rect 276216 154426 276244 163200
rect 277136 156942 277164 163200
rect 277124 156936 277176 156942
rect 277124 156878 277176 156884
rect 277124 156188 277176 156194
rect 277124 156130 277176 156136
rect 276204 154420 276256 154426
rect 276204 154362 276256 154368
rect 276124 151786 276520 151814
rect 276492 150226 276520 151786
rect 277136 150226 277164 156130
rect 277412 152114 277440 163254
rect 277872 163146 277900 163254
rect 277950 163200 278006 164400
rect 278778 163200 278834 164400
rect 278884 163254 279556 163282
rect 277964 163146 277992 163200
rect 277872 163118 277992 163146
rect 278412 154352 278464 154358
rect 278412 154294 278464 154300
rect 277768 152924 277820 152930
rect 277768 152866 277820 152872
rect 277400 152108 277452 152114
rect 277400 152050 277452 152056
rect 277780 150226 277808 152866
rect 278424 150226 278452 154294
rect 278792 152930 278820 163200
rect 278884 154358 278912 163254
rect 279528 163146 279556 163254
rect 279606 163200 279662 164400
rect 280434 163200 280490 164400
rect 281262 163200 281318 164400
rect 282090 163200 282146 164400
rect 283010 163200 283066 164400
rect 283116 163254 283328 163282
rect 279620 163146 279648 163200
rect 279528 163118 279648 163146
rect 280344 160064 280396 160070
rect 280344 160006 280396 160012
rect 279056 156392 279108 156398
rect 279056 156334 279108 156340
rect 278872 154352 278924 154358
rect 278872 154294 278924 154300
rect 278780 152924 278832 152930
rect 278780 152866 278832 152872
rect 279068 150226 279096 156334
rect 279700 153196 279752 153202
rect 279700 153138 279752 153144
rect 279712 150226 279740 153138
rect 280356 150226 280384 160006
rect 280448 157078 280476 163200
rect 281276 160070 281304 163200
rect 281264 160064 281316 160070
rect 281264 160006 281316 160012
rect 282104 159322 282132 163200
rect 283024 163146 283052 163200
rect 283116 163146 283144 163254
rect 283024 163118 283144 163146
rect 281540 159316 281592 159322
rect 281540 159258 281592 159264
rect 282092 159316 282144 159322
rect 282092 159258 282144 159264
rect 280436 157072 280488 157078
rect 280436 157014 280488 157020
rect 280986 153776 281042 153785
rect 280986 153711 281042 153720
rect 281000 150226 281028 153711
rect 264382 150146 264434 150152
rect 264394 149940 264422 150146
rect 265038 149940 265066 150198
rect 265682 149940 265710 150198
rect 266326 149940 266354 150198
rect 266970 149940 266998 150198
rect 267614 149940 267642 150198
rect 268258 149940 268286 150198
rect 268902 149940 268930 150198
rect 269120 150204 269172 150210
rect 269500 150198 269574 150226
rect 269120 150146 269172 150152
rect 269546 149940 269574 150198
rect 270178 150204 270230 150210
rect 270788 150198 270862 150226
rect 271432 150198 271506 150226
rect 272076 150198 272150 150226
rect 272720 150198 272794 150226
rect 273272 150198 273346 150226
rect 273916 150198 273990 150226
rect 274560 150198 274634 150226
rect 275204 150198 275278 150226
rect 275848 150198 275922 150226
rect 276492 150198 276566 150226
rect 277136 150198 277210 150226
rect 277780 150198 277854 150226
rect 278424 150198 278498 150226
rect 279068 150198 279142 150226
rect 279712 150198 279786 150226
rect 280356 150198 280430 150226
rect 281000 150198 281074 150226
rect 281552 150210 281580 159258
rect 283196 159112 283248 159118
rect 283196 159054 283248 159060
rect 281632 157344 281684 157350
rect 281632 157286 281684 157292
rect 281644 150226 281672 157286
rect 283104 156664 283156 156670
rect 283104 156606 283156 156612
rect 282920 152244 282972 152250
rect 282920 152186 282972 152192
rect 282932 150226 282960 152186
rect 270178 150146 270230 150152
rect 270190 149940 270218 150146
rect 270834 149940 270862 150198
rect 271478 149940 271506 150198
rect 272122 149940 272150 150198
rect 272766 149940 272794 150198
rect 273318 149940 273346 150198
rect 273962 149940 273990 150198
rect 274606 149940 274634 150198
rect 275250 149940 275278 150198
rect 275894 149940 275922 150198
rect 276538 149940 276566 150198
rect 277182 149940 277210 150198
rect 277826 149940 277854 150198
rect 278470 149940 278498 150198
rect 279114 149940 279142 150198
rect 279758 149940 279786 150198
rect 280402 149940 280430 150198
rect 281046 149940 281074 150198
rect 281540 150204 281592 150210
rect 281644 150198 281718 150226
rect 281540 150146 281592 150152
rect 281690 149940 281718 150198
rect 282322 150204 282374 150210
rect 282932 150198 283006 150226
rect 283116 150210 283144 156606
rect 283208 151842 283236 159054
rect 283300 154494 283328 163254
rect 283838 163200 283894 164400
rect 284666 163200 284722 164400
rect 285494 163200 285550 164400
rect 285692 163254 286272 163282
rect 283852 157282 283880 163200
rect 284392 159248 284444 159254
rect 284392 159190 284444 159196
rect 283840 157276 283892 157282
rect 283840 157218 283892 157224
rect 283656 154556 283708 154562
rect 283656 154498 283708 154504
rect 283288 154488 283340 154494
rect 283288 154430 283340 154436
rect 283196 151836 283248 151842
rect 283196 151778 283248 151784
rect 283668 150226 283696 154498
rect 282322 150146 282374 150152
rect 282334 149940 282362 150146
rect 282978 149940 283006 150198
rect 283104 150204 283156 150210
rect 283104 150146 283156 150152
rect 283622 150198 283696 150226
rect 284404 150210 284432 159190
rect 284680 159118 284708 163200
rect 284668 159112 284720 159118
rect 284668 159054 284720 159060
rect 285508 153202 285536 163200
rect 285692 154562 285720 163254
rect 286244 163146 286272 163254
rect 286322 163200 286378 164400
rect 287150 163200 287206 164400
rect 287978 163200 288034 164400
rect 288898 163200 288954 164400
rect 289726 163200 289782 164400
rect 290554 163200 290610 164400
rect 291382 163200 291438 164400
rect 292210 163200 292266 164400
rect 293038 163200 293094 164400
rect 293866 163200 293922 164400
rect 294786 163200 294842 164400
rect 295614 163200 295670 164400
rect 296442 163200 296498 164400
rect 297270 163200 297326 164400
rect 298098 163200 298154 164400
rect 298664 163254 298876 163282
rect 286336 163146 286364 163200
rect 286244 163118 286364 163146
rect 285772 159112 285824 159118
rect 285772 159054 285824 159060
rect 285588 154556 285640 154562
rect 285588 154498 285640 154504
rect 285680 154556 285732 154562
rect 285680 154498 285732 154504
rect 285600 154442 285628 154498
rect 285600 154414 285720 154442
rect 285496 153196 285548 153202
rect 285496 153138 285548 153144
rect 284852 152992 284904 152998
rect 284852 152934 284904 152940
rect 284864 150226 284892 152934
rect 285692 151814 285720 154414
rect 285784 152250 285812 159054
rect 287164 157146 287192 163200
rect 287992 159254 288020 163200
rect 287980 159248 288032 159254
rect 287980 159190 288032 159196
rect 288912 159118 288940 163200
rect 288072 159112 288124 159118
rect 288072 159054 288124 159060
rect 288900 159112 288952 159118
rect 288900 159054 288952 159060
rect 287152 157140 287204 157146
rect 287152 157082 287204 157088
rect 286232 156324 286284 156330
rect 286232 156266 286284 156272
rect 285772 152244 285824 152250
rect 285772 152186 285824 152192
rect 286244 151814 286272 156266
rect 288084 152998 288112 159054
rect 289360 156732 289412 156738
rect 289360 156674 289412 156680
rect 288716 154012 288768 154018
rect 288716 153954 288768 153960
rect 288072 152992 288124 152998
rect 288072 152934 288124 152940
rect 288072 152380 288124 152386
rect 288072 152322 288124 152328
rect 287428 151836 287480 151842
rect 285692 151786 286180 151814
rect 286244 151786 286824 151814
rect 286152 150226 286180 151786
rect 286796 150226 286824 151786
rect 287428 151778 287480 151784
rect 287440 150226 287468 151778
rect 288084 150226 288112 152322
rect 288728 150226 288756 153954
rect 289372 150226 289400 156674
rect 289740 155786 289768 163200
rect 290568 157214 290596 163200
rect 290648 159180 290700 159186
rect 290648 159122 290700 159128
rect 290556 157208 290608 157214
rect 290556 157150 290608 157156
rect 289728 155780 289780 155786
rect 289728 155722 289780 155728
rect 290004 152992 290056 152998
rect 290004 152934 290056 152940
rect 290016 150226 290044 152934
rect 290660 150226 290688 159122
rect 291292 153944 291344 153950
rect 291292 153886 291344 153892
rect 291304 150226 291332 153886
rect 291396 152386 291424 163200
rect 291936 156868 291988 156874
rect 291936 156810 291988 156816
rect 291384 152380 291436 152386
rect 291384 152322 291436 152328
rect 291948 150226 291976 156810
rect 292224 152998 292252 163200
rect 293052 155854 293080 163200
rect 293880 156738 293908 163200
rect 294800 159526 294828 163200
rect 293960 159520 294012 159526
rect 293960 159462 294012 159468
rect 294788 159520 294840 159526
rect 294788 159462 294840 159468
rect 293972 159186 294000 159462
rect 295628 159390 295656 163200
rect 295524 159384 295576 159390
rect 295524 159326 295576 159332
rect 295616 159384 295668 159390
rect 295616 159326 295668 159332
rect 293960 159180 294012 159186
rect 293960 159122 294012 159128
rect 295156 159180 295208 159186
rect 295156 159122 295208 159128
rect 294052 156800 294104 156806
rect 294052 156742 294104 156748
rect 293868 156732 293920 156738
rect 293868 156674 293920 156680
rect 293040 155848 293092 155854
rect 293040 155790 293092 155796
rect 293868 153672 293920 153678
rect 293868 153614 293920 153620
rect 292212 152992 292264 152998
rect 292212 152934 292264 152940
rect 293224 152516 293276 152522
rect 293224 152458 293276 152464
rect 292578 152416 292634 152425
rect 292578 152351 292634 152360
rect 292592 150226 292620 152351
rect 293236 150226 293264 152458
rect 293880 150226 293908 153614
rect 294064 151814 294092 156742
rect 294064 151786 294552 151814
rect 294524 150226 294552 151786
rect 295168 150226 295196 159122
rect 295536 151814 295564 159326
rect 296456 155922 296484 163200
rect 297284 156806 297312 163200
rect 298008 159452 298060 159458
rect 298008 159394 298060 159400
rect 297272 156800 297324 156806
rect 297272 156742 297324 156748
rect 296444 155916 296496 155922
rect 296444 155858 296496 155864
rect 297088 155304 297140 155310
rect 297088 155246 297140 155252
rect 296444 153808 296496 153814
rect 296444 153750 296496 153756
rect 295536 151786 295840 151814
rect 295812 150226 295840 151786
rect 296456 150226 296484 153750
rect 297100 150226 297128 155246
rect 297732 152584 297784 152590
rect 297732 152526 297784 152532
rect 297744 150226 297772 152526
rect 298020 151814 298048 159394
rect 298112 159050 298140 163200
rect 298100 159044 298152 159050
rect 298100 158986 298152 158992
rect 298664 152522 298692 163254
rect 298848 163146 298876 163254
rect 298926 163200 298982 164400
rect 299754 163200 299810 164400
rect 300674 163200 300730 164400
rect 301502 163200 301558 164400
rect 302330 163200 302386 164400
rect 303158 163200 303214 164400
rect 303632 163254 303936 163282
rect 298940 163146 298968 163200
rect 298848 163118 298968 163146
rect 299480 158976 299532 158982
rect 299480 158918 299532 158924
rect 299020 153740 299072 153746
rect 299020 153682 299072 153688
rect 298652 152516 298704 152522
rect 298652 152458 298704 152464
rect 298020 151786 298416 151814
rect 298388 150226 298416 151786
rect 299032 150226 299060 153682
rect 284254 150204 284306 150210
rect 283622 149940 283650 150198
rect 284254 150146 284306 150152
rect 284392 150204 284444 150210
rect 284864 150198 284938 150226
rect 284392 150146 284444 150152
rect 284266 149940 284294 150146
rect 284910 149940 284938 150198
rect 285542 150204 285594 150210
rect 286152 150198 286226 150226
rect 286796 150198 286870 150226
rect 287440 150198 287514 150226
rect 288084 150198 288158 150226
rect 288728 150198 288802 150226
rect 289372 150198 289446 150226
rect 290016 150198 290090 150226
rect 290660 150198 290734 150226
rect 291304 150198 291378 150226
rect 291948 150198 292022 150226
rect 292592 150198 292666 150226
rect 293236 150198 293310 150226
rect 293880 150198 293954 150226
rect 294524 150198 294598 150226
rect 295168 150198 295242 150226
rect 295812 150198 295886 150226
rect 296456 150198 296530 150226
rect 297100 150198 297174 150226
rect 297744 150198 297818 150226
rect 298388 150198 298462 150226
rect 299032 150198 299106 150226
rect 299492 150210 299520 158918
rect 299664 158024 299716 158030
rect 299664 157966 299716 157972
rect 299676 150226 299704 157966
rect 299768 155310 299796 163200
rect 300400 159044 300452 159050
rect 300400 158986 300452 158992
rect 299756 155304 299808 155310
rect 299756 155246 299808 155252
rect 300412 151842 300440 158986
rect 300688 156874 300716 163200
rect 301516 159458 301544 163200
rect 301504 159452 301556 159458
rect 301504 159394 301556 159400
rect 302344 159186 302372 163200
rect 302332 159180 302384 159186
rect 302332 159122 302384 159128
rect 300676 156868 300728 156874
rect 300676 156810 300728 156816
rect 302516 155236 302568 155242
rect 302516 155178 302568 155184
rect 301596 153604 301648 153610
rect 301596 153546 301648 153552
rect 300952 152040 301004 152046
rect 300952 151982 301004 151988
rect 300400 151836 300452 151842
rect 300400 151778 300452 151784
rect 300964 150226 300992 151982
rect 301608 150226 301636 153546
rect 302528 151814 302556 155178
rect 303172 155106 303200 163200
rect 303528 158908 303580 158914
rect 303528 158850 303580 158856
rect 303160 155100 303212 155106
rect 303160 155042 303212 155048
rect 302884 151972 302936 151978
rect 302884 151914 302936 151920
rect 302344 151786 302556 151814
rect 302344 150226 302372 151786
rect 285542 150146 285594 150152
rect 285554 149940 285582 150146
rect 286198 149940 286226 150198
rect 286842 149940 286870 150198
rect 287486 149940 287514 150198
rect 288130 149940 288158 150198
rect 288774 149940 288802 150198
rect 289418 149940 289446 150198
rect 290062 149940 290090 150198
rect 290706 149940 290734 150198
rect 291350 149940 291378 150198
rect 291994 149940 292022 150198
rect 292638 149940 292666 150198
rect 293282 149940 293310 150198
rect 293926 149940 293954 150198
rect 294570 149940 294598 150198
rect 295214 149940 295242 150198
rect 295858 149940 295886 150198
rect 296502 149940 296530 150198
rect 297146 149940 297174 150198
rect 297790 149940 297818 150198
rect 298434 149940 298462 150198
rect 299078 149940 299106 150198
rect 299480 150204 299532 150210
rect 299676 150198 299750 150226
rect 299480 150146 299532 150152
rect 299722 149940 299750 150198
rect 300354 150204 300406 150210
rect 300964 150198 301038 150226
rect 301608 150198 301682 150226
rect 300354 150146 300406 150152
rect 300366 149940 300394 150146
rect 301010 149940 301038 150198
rect 301654 149940 301682 150198
rect 302298 150198 302372 150226
rect 302896 150226 302924 151914
rect 303540 150226 303568 158850
rect 303632 152590 303660 163254
rect 303908 163146 303936 163254
rect 303986 163200 304042 164400
rect 304184 163254 304764 163282
rect 304000 163146 304028 163200
rect 303908 163118 304028 163146
rect 304080 153876 304132 153882
rect 304080 153818 304132 153824
rect 303620 152584 303672 152590
rect 303620 152526 303672 152532
rect 304092 150226 304120 153818
rect 304184 152046 304212 163254
rect 304736 163146 304764 163254
rect 304814 163200 304870 164400
rect 305642 163200 305698 164400
rect 306562 163200 306618 164400
rect 307390 163200 307446 164400
rect 308218 163200 308274 164400
rect 309046 163200 309102 164400
rect 309152 163254 309824 163282
rect 304828 163146 304856 163200
rect 304736 163118 304856 163146
rect 305368 159656 305420 159662
rect 305368 159598 305420 159604
rect 304724 158092 304776 158098
rect 304724 158034 304776 158040
rect 304172 152040 304224 152046
rect 304172 151982 304224 151988
rect 304736 150226 304764 158034
rect 305380 150226 305408 159598
rect 305656 158914 305684 163200
rect 305644 158908 305696 158914
rect 305644 158850 305696 158856
rect 306576 155242 306604 163200
rect 307404 159050 307432 163200
rect 308232 159730 308260 163200
rect 308220 159724 308272 159730
rect 308220 159666 308272 159672
rect 309060 159662 309088 163200
rect 308588 159656 308640 159662
rect 308588 159598 308640 159604
rect 309048 159656 309100 159662
rect 309048 159598 309100 159604
rect 307392 159044 307444 159050
rect 307392 158986 307444 158992
rect 307668 158908 307720 158914
rect 307668 158850 307720 158856
rect 306932 158160 306984 158166
rect 306932 158102 306984 158108
rect 306564 155236 306616 155242
rect 306564 155178 306616 155184
rect 306656 154148 306708 154154
rect 306656 154090 306708 154096
rect 306012 152176 306064 152182
rect 306012 152118 306064 152124
rect 306024 150226 306052 152118
rect 306668 150226 306696 154090
rect 306944 151814 306972 158102
rect 307680 151978 307708 158850
rect 307944 152652 307996 152658
rect 307944 152594 307996 152600
rect 307668 151972 307720 151978
rect 307668 151914 307720 151920
rect 306944 151786 307340 151814
rect 307312 150226 307340 151786
rect 307956 150226 307984 152594
rect 308600 150226 308628 159598
rect 309152 153882 309180 163254
rect 309796 163146 309824 163254
rect 309874 163200 309930 164400
rect 310702 163200 310758 164400
rect 311530 163200 311586 164400
rect 312450 163200 312506 164400
rect 313278 163200 313334 164400
rect 314106 163200 314162 164400
rect 314934 163200 314990 164400
rect 315762 163200 315818 164400
rect 316052 163254 316540 163282
rect 309888 163146 309916 163200
rect 309796 163118 309916 163146
rect 310612 159588 310664 159594
rect 310612 159530 310664 159536
rect 309876 155372 309928 155378
rect 309876 155314 309928 155320
rect 309232 154080 309284 154086
rect 309232 154022 309284 154028
rect 309140 153876 309192 153882
rect 309140 153818 309192 153824
rect 309244 150226 309272 154022
rect 309888 150226 309916 155314
rect 310624 150226 310652 159530
rect 310716 158914 310744 163200
rect 310704 158908 310756 158914
rect 310704 158850 310756 158856
rect 311164 152720 311216 152726
rect 311164 152662 311216 152668
rect 302896 150198 302970 150226
rect 303540 150198 303614 150226
rect 304092 150198 304166 150226
rect 304736 150198 304810 150226
rect 305380 150198 305454 150226
rect 306024 150198 306098 150226
rect 306668 150198 306742 150226
rect 307312 150198 307386 150226
rect 307956 150198 308030 150226
rect 308600 150198 308674 150226
rect 309244 150198 309318 150226
rect 309888 150198 309962 150226
rect 302298 149940 302326 150198
rect 302942 149940 302970 150198
rect 303586 149940 303614 150198
rect 304138 149940 304166 150198
rect 304782 149940 304810 150198
rect 305426 149940 305454 150198
rect 306070 149940 306098 150198
rect 306714 149940 306742 150198
rect 307358 149940 307386 150198
rect 308002 149940 308030 150198
rect 308646 149940 308674 150198
rect 309290 149940 309318 150198
rect 309934 149940 309962 150198
rect 310578 150198 310652 150226
rect 311176 150226 311204 152662
rect 311544 152658 311572 163200
rect 312464 158914 312492 163200
rect 312176 158908 312228 158914
rect 312176 158850 312228 158856
rect 312452 158908 312504 158914
rect 312452 158850 312504 158856
rect 311808 153536 311860 153542
rect 311808 153478 311860 153484
rect 311532 152652 311584 152658
rect 311532 152594 311584 152600
rect 311820 150226 311848 153478
rect 312188 152726 312216 158850
rect 312452 155440 312504 155446
rect 312452 155382 312504 155388
rect 312176 152720 312228 152726
rect 312176 152662 312228 152668
rect 312464 150226 312492 155382
rect 313292 153950 313320 163200
rect 314120 159798 314148 163200
rect 313464 159792 313516 159798
rect 313464 159734 313516 159740
rect 314108 159792 314160 159798
rect 314108 159734 314160 159740
rect 313372 158908 313424 158914
rect 313372 158850 313424 158856
rect 313280 153944 313332 153950
rect 313280 153886 313332 153892
rect 313096 152856 313148 152862
rect 313096 152798 313148 152804
rect 313108 150226 313136 152798
rect 313384 152425 313412 158850
rect 313370 152416 313426 152425
rect 313370 152351 313426 152360
rect 313476 151814 313504 159734
rect 314948 158982 314976 163200
rect 315776 159594 315804 163200
rect 315764 159588 315816 159594
rect 315764 159530 315816 159536
rect 314936 158976 314988 158982
rect 314936 158918 314988 158924
rect 315028 158228 315080 158234
rect 315028 158170 315080 158176
rect 314384 154216 314436 154222
rect 314384 154158 314436 154164
rect 313476 151786 313780 151814
rect 313752 150226 313780 151786
rect 314396 150226 314424 154158
rect 315040 150226 315068 158170
rect 316052 154018 316080 163254
rect 316512 163146 316540 163254
rect 316590 163200 316646 164400
rect 317418 163200 317474 164400
rect 317524 163254 318288 163282
rect 316604 163146 316632 163200
rect 316512 163118 316632 163146
rect 317052 158840 317104 158846
rect 317052 158782 317104 158788
rect 316040 154012 316092 154018
rect 316040 153954 316092 153960
rect 316960 153400 317012 153406
rect 316960 153342 317012 153348
rect 315672 152788 315724 152794
rect 315672 152730 315724 152736
rect 315684 150226 315712 152730
rect 316316 152448 316368 152454
rect 316316 152390 316368 152396
rect 316328 150226 316356 152390
rect 316972 150226 317000 153342
rect 317064 152862 317092 158782
rect 317052 152856 317104 152862
rect 317052 152798 317104 152804
rect 317432 152794 317460 163200
rect 317420 152788 317472 152794
rect 317420 152730 317472 152736
rect 317524 152454 317552 163254
rect 318260 163146 318288 163254
rect 318338 163200 318394 164400
rect 319166 163200 319222 164400
rect 319994 163200 320050 164400
rect 320822 163200 320878 164400
rect 321650 163200 321706 164400
rect 322478 163200 322534 164400
rect 323306 163200 323362 164400
rect 324226 163200 324282 164400
rect 324332 163254 325004 163282
rect 318352 163146 318380 163200
rect 318260 163118 318380 163146
rect 318892 159860 318944 159866
rect 318892 159802 318944 159808
rect 317604 155508 317656 155514
rect 317604 155450 317656 155456
rect 317512 152448 317564 152454
rect 317512 152390 317564 152396
rect 317616 150226 317644 155450
rect 318248 152856 318300 152862
rect 318248 152798 318300 152804
rect 318260 150226 318288 152798
rect 318904 150226 318932 159802
rect 319180 158846 319208 163200
rect 319168 158840 319220 158846
rect 319168 158782 319220 158788
rect 320008 155378 320036 163200
rect 320836 159866 320864 163200
rect 320824 159860 320876 159866
rect 320824 159802 320876 159808
rect 321560 158840 321612 158846
rect 321560 158782 321612 158788
rect 320272 158772 320324 158778
rect 320272 158714 320324 158720
rect 320180 155576 320232 155582
rect 320180 155518 320232 155524
rect 319996 155372 320048 155378
rect 319996 155314 320048 155320
rect 319536 154284 319588 154290
rect 319536 154226 319588 154232
rect 319548 150226 319576 154226
rect 320192 150226 320220 155518
rect 320284 152862 320312 158714
rect 321468 153128 321520 153134
rect 321468 153070 321520 153076
rect 320272 152856 320324 152862
rect 320272 152798 320324 152804
rect 320652 152748 320956 152776
rect 320652 152454 320680 152748
rect 320928 152658 320956 152748
rect 320824 152652 320876 152658
rect 320824 152594 320876 152600
rect 320916 152652 320968 152658
rect 320916 152594 320968 152600
rect 320640 152448 320692 152454
rect 320640 152390 320692 152396
rect 320732 152448 320784 152454
rect 320732 152390 320784 152396
rect 320744 151910 320772 152390
rect 320836 152182 320864 152594
rect 320916 152312 320968 152318
rect 320916 152254 320968 152260
rect 320824 152176 320876 152182
rect 320824 152118 320876 152124
rect 320732 151904 320784 151910
rect 320732 151846 320784 151852
rect 320928 150226 320956 152254
rect 311176 150198 311250 150226
rect 311820 150198 311894 150226
rect 312464 150198 312538 150226
rect 313108 150198 313182 150226
rect 313752 150198 313826 150226
rect 314396 150198 314470 150226
rect 315040 150198 315114 150226
rect 315684 150198 315758 150226
rect 316328 150198 316402 150226
rect 316972 150198 317046 150226
rect 317616 150198 317690 150226
rect 318260 150198 318334 150226
rect 318904 150198 318978 150226
rect 319548 150198 319622 150226
rect 320192 150198 320266 150226
rect 310578 149940 310606 150198
rect 311222 149940 311250 150198
rect 311866 149940 311894 150198
rect 312510 149940 312538 150198
rect 313154 149940 313182 150198
rect 313798 149940 313826 150198
rect 314442 149940 314470 150198
rect 315086 149940 315114 150198
rect 315730 149940 315758 150198
rect 316374 149940 316402 150198
rect 317018 149940 317046 150198
rect 317662 149940 317690 150198
rect 318306 149940 318334 150198
rect 318950 149940 318978 150198
rect 319594 149940 319622 150198
rect 320238 149940 320266 150198
rect 320882 150198 320956 150226
rect 321480 150226 321508 153070
rect 321572 151910 321600 158782
rect 321664 158778 321692 163200
rect 322492 158914 322520 163200
rect 322480 158908 322532 158914
rect 322480 158850 322532 158856
rect 321652 158772 321704 158778
rect 321652 158714 321704 158720
rect 322112 155644 322164 155650
rect 322112 155586 322164 155592
rect 322020 153468 322072 153474
rect 322020 153410 322072 153416
rect 321560 151904 321612 151910
rect 321560 151846 321612 151852
rect 322032 150498 322060 153410
rect 322124 151814 322152 155586
rect 323320 154086 323348 163200
rect 324044 159928 324096 159934
rect 324044 159870 324096 159876
rect 323308 154080 323360 154086
rect 323308 154022 323360 154028
rect 323124 152856 323176 152862
rect 323124 152798 323176 152804
rect 323136 151814 323164 152798
rect 322124 151786 322796 151814
rect 323136 151786 323440 151814
rect 322032 150470 322152 150498
rect 322124 150226 322152 150470
rect 322768 150226 322796 151786
rect 323412 150226 323440 151786
rect 324056 150226 324084 159870
rect 324240 152862 324268 163200
rect 324332 153134 324360 163254
rect 324976 163146 325004 163254
rect 325054 163200 325110 164400
rect 325882 163200 325938 164400
rect 326710 163200 326766 164400
rect 327538 163200 327594 164400
rect 328366 163200 328422 164400
rect 329194 163200 329250 164400
rect 330114 163200 330170 164400
rect 330942 163200 330998 164400
rect 331232 163254 331720 163282
rect 325068 163146 325096 163200
rect 324976 163118 325096 163146
rect 325896 161474 325924 163200
rect 325896 161446 326108 161474
rect 325332 155712 325384 155718
rect 325332 155654 325384 155660
rect 324688 153264 324740 153270
rect 324688 153206 324740 153212
rect 324320 153128 324372 153134
rect 324320 153070 324372 153076
rect 324228 152856 324280 152862
rect 324228 152798 324280 152804
rect 324700 150226 324728 153206
rect 325344 150226 325372 155654
rect 326080 152454 326108 161446
rect 326724 154154 326752 163200
rect 327552 158846 327580 163200
rect 328380 159934 328408 163200
rect 329208 160002 329236 163200
rect 329104 159996 329156 160002
rect 329104 159938 329156 159944
rect 329196 159996 329248 160002
rect 329196 159938 329248 159944
rect 328368 159928 328420 159934
rect 328368 159870 328420 159876
rect 328550 159488 328606 159497
rect 328550 159423 328606 159432
rect 327540 158840 327592 158846
rect 327540 158782 327592 158788
rect 327908 157004 327960 157010
rect 327908 156946 327960 156952
rect 326712 154148 326764 154154
rect 326712 154090 326764 154096
rect 327264 153332 327316 153338
rect 327264 153274 327316 153280
rect 326620 153060 326672 153066
rect 326620 153002 326672 153008
rect 325976 152448 326028 152454
rect 325976 152390 326028 152396
rect 326068 152448 326120 152454
rect 326068 152390 326120 152396
rect 325988 150226 326016 152390
rect 326632 150226 326660 153002
rect 327276 150226 327304 153274
rect 327920 150226 327948 156946
rect 328564 150226 328592 159423
rect 329116 151814 329144 159938
rect 330128 155446 330156 163200
rect 330484 158840 330536 158846
rect 330536 158788 330708 158794
rect 330484 158782 330708 158788
rect 330496 158778 330708 158782
rect 330496 158772 330720 158778
rect 330496 158766 330668 158772
rect 330668 158714 330720 158720
rect 330484 156936 330536 156942
rect 330484 156878 330536 156884
rect 330116 155440 330168 155446
rect 330116 155382 330168 155388
rect 329932 154420 329984 154426
rect 329932 154362 329984 154368
rect 329116 151786 329236 151814
rect 329208 150226 329236 151786
rect 329944 150226 329972 154362
rect 321480 150198 321554 150226
rect 322124 150198 322198 150226
rect 322768 150198 322842 150226
rect 323412 150198 323486 150226
rect 324056 150198 324130 150226
rect 324700 150198 324774 150226
rect 325344 150198 325418 150226
rect 325988 150198 326062 150226
rect 326632 150198 326706 150226
rect 327276 150198 327350 150226
rect 327920 150198 327994 150226
rect 328564 150198 328638 150226
rect 329208 150198 329282 150226
rect 320882 149940 320910 150198
rect 321526 149940 321554 150198
rect 322170 149940 322198 150198
rect 322814 149940 322842 150198
rect 323458 149940 323486 150198
rect 324102 149940 324130 150198
rect 324746 149940 324774 150198
rect 325390 149940 325418 150198
rect 326034 149940 326062 150198
rect 326678 149940 326706 150198
rect 327322 149940 327350 150198
rect 327966 149940 327994 150198
rect 328610 149940 328638 150198
rect 329254 149940 329282 150198
rect 329898 150198 329972 150226
rect 330496 150226 330524 156878
rect 330956 153066 330984 163200
rect 330944 153060 330996 153066
rect 330944 153002 330996 153008
rect 331232 152318 331260 163254
rect 331692 163146 331720 163254
rect 331770 163200 331826 164400
rect 332598 163200 332654 164400
rect 333426 163200 333482 164400
rect 334254 163200 334310 164400
rect 335082 163200 335138 164400
rect 335372 163254 335952 163282
rect 331784 163146 331812 163200
rect 331692 163118 331812 163146
rect 332416 154352 332468 154358
rect 332416 154294 332468 154300
rect 331772 152924 331824 152930
rect 331772 152866 331824 152872
rect 331220 152312 331272 152318
rect 331220 152254 331272 152260
rect 331128 152108 331180 152114
rect 331128 152050 331180 152056
rect 331140 150226 331168 152050
rect 331784 150226 331812 152866
rect 332428 150226 332456 154294
rect 332612 152930 332640 163200
rect 332692 160064 332744 160070
rect 332692 160006 332744 160012
rect 332600 152924 332652 152930
rect 332600 152866 332652 152872
rect 330496 150198 330570 150226
rect 331140 150198 331214 150226
rect 331784 150198 331858 150226
rect 332428 150198 332502 150226
rect 332704 150210 332732 160006
rect 333060 157072 333112 157078
rect 333060 157014 333112 157020
rect 333072 150226 333100 157014
rect 333440 155514 333468 163200
rect 334268 160070 334296 163200
rect 334256 160064 334308 160070
rect 334256 160006 334308 160012
rect 335096 159322 335124 163200
rect 334348 159316 334400 159322
rect 334348 159258 334400 159264
rect 335084 159316 335136 159322
rect 335084 159258 335136 159264
rect 333428 155508 333480 155514
rect 333428 155450 333480 155456
rect 334360 150226 334388 159258
rect 334900 154488 334952 154494
rect 334900 154430 334952 154436
rect 334912 150226 334940 154430
rect 335372 152114 335400 163254
rect 335924 163146 335952 163254
rect 336002 163200 336058 164400
rect 336830 163200 336886 164400
rect 337658 163200 337714 164400
rect 338486 163200 338542 164400
rect 339314 163200 339370 164400
rect 339512 163254 340092 163282
rect 336016 163146 336044 163200
rect 335924 163118 336044 163146
rect 335544 157276 335596 157282
rect 335544 157218 335596 157224
rect 335360 152108 335412 152114
rect 335360 152050 335412 152056
rect 335556 150226 335584 157218
rect 336844 154222 336872 163200
rect 337672 155582 337700 163200
rect 338500 159118 338528 163200
rect 339328 159254 339356 163200
rect 338764 159248 338816 159254
rect 338764 159190 338816 159196
rect 339316 159248 339368 159254
rect 339316 159190 339368 159196
rect 338304 159112 338356 159118
rect 338304 159054 338356 159060
rect 338488 159112 338540 159118
rect 338488 159054 338540 159060
rect 338120 157140 338172 157146
rect 338120 157082 338172 157088
rect 337660 155576 337712 155582
rect 337660 155518 337712 155524
rect 337476 154556 337528 154562
rect 337476 154498 337528 154504
rect 336832 154216 336884 154222
rect 336832 154158 336884 154164
rect 336832 153196 336884 153202
rect 336832 153138 336884 153144
rect 336188 152244 336240 152250
rect 336188 152186 336240 152192
rect 336200 150226 336228 152186
rect 336844 150226 336872 153138
rect 337488 150226 337516 154498
rect 338132 150226 338160 157082
rect 329898 149940 329926 150198
rect 330542 149940 330570 150198
rect 331186 149940 331214 150198
rect 331830 149940 331858 150198
rect 332474 149940 332502 150198
rect 332692 150204 332744 150210
rect 333072 150198 333146 150226
rect 332692 150146 332744 150152
rect 333118 149940 333146 150198
rect 333750 150204 333802 150210
rect 334360 150198 334434 150226
rect 334912 150198 334986 150226
rect 335556 150198 335630 150226
rect 336200 150198 336274 150226
rect 336844 150198 336918 150226
rect 337488 150198 337562 150226
rect 338132 150198 338206 150226
rect 338316 150210 338344 159054
rect 338776 150226 338804 159190
rect 339512 154290 339540 163254
rect 340064 163146 340092 163254
rect 340142 163200 340198 164400
rect 340970 163200 341026 164400
rect 341890 163200 341946 164400
rect 341996 163254 342208 163282
rect 340156 163146 340184 163200
rect 340064 163118 340184 163146
rect 339684 159112 339736 159118
rect 339684 159054 339736 159060
rect 339592 155780 339644 155786
rect 339592 155722 339644 155728
rect 339500 154284 339552 154290
rect 339500 154226 339552 154232
rect 339604 151814 339632 155722
rect 339696 153202 339724 159054
rect 340052 157208 340104 157214
rect 340052 157150 340104 157156
rect 339684 153196 339736 153202
rect 339684 153138 339736 153144
rect 340064 151814 340092 157150
rect 340984 155650 341012 163200
rect 341904 163146 341932 163200
rect 341996 163146 342024 163254
rect 341904 163118 342024 163146
rect 341616 159656 341668 159662
rect 341616 159598 341668 159604
rect 342180 159610 342208 163254
rect 342718 163200 342774 164400
rect 343546 163200 343602 164400
rect 344374 163200 344430 164400
rect 345202 163200 345258 164400
rect 346030 163200 346086 164400
rect 346412 163254 346808 163282
rect 342732 159730 342760 163200
rect 342628 159724 342680 159730
rect 342628 159666 342680 159672
rect 342720 159724 342772 159730
rect 342720 159666 342772 159672
rect 342640 159610 342668 159666
rect 342812 159656 342864 159662
rect 341628 159526 341656 159598
rect 342180 159582 342392 159610
rect 342640 159604 342812 159610
rect 342640 159598 342864 159604
rect 342640 159582 342852 159598
rect 341616 159520 341668 159526
rect 341616 159462 341668 159468
rect 342364 159458 342392 159582
rect 341432 159452 341484 159458
rect 341432 159394 341484 159400
rect 342260 159452 342312 159458
rect 342260 159394 342312 159400
rect 342352 159452 342404 159458
rect 342352 159394 342404 159400
rect 341444 159186 341472 159394
rect 341432 159180 341484 159186
rect 341432 159122 341484 159128
rect 340972 155644 341024 155650
rect 340972 155586 341024 155592
rect 342272 152998 342300 159394
rect 342444 159384 342496 159390
rect 342444 159326 342496 159332
rect 342352 155848 342404 155854
rect 342352 155790 342404 155796
rect 341984 152992 342036 152998
rect 341984 152934 342036 152940
rect 342260 152992 342312 152998
rect 342260 152934 342312 152940
rect 341340 152380 341392 152386
rect 341340 152322 341392 152328
rect 339604 151786 340000 151814
rect 340064 151786 340736 151814
rect 339972 150226 340000 151786
rect 340708 150226 340736 151786
rect 341352 150226 341380 152322
rect 341996 150226 342024 152934
rect 342364 151814 342392 155790
rect 342456 152250 342484 159326
rect 342536 156732 342588 156738
rect 342536 156674 342588 156680
rect 342444 152244 342496 152250
rect 342444 152186 342496 152192
rect 342548 151814 342576 156674
rect 343560 154358 343588 163200
rect 343824 159724 343876 159730
rect 343824 159666 343876 159672
rect 343548 154352 343600 154358
rect 343548 154294 343600 154300
rect 343836 152386 343864 159666
rect 344388 155718 344416 163200
rect 345216 157334 345244 163200
rect 346044 159390 346072 163200
rect 346032 159384 346084 159390
rect 345584 159310 345796 159338
rect 346032 159326 346084 159332
rect 345584 159050 345612 159310
rect 345768 159186 345796 159310
rect 345664 159180 345716 159186
rect 345664 159122 345716 159128
rect 345756 159180 345808 159186
rect 345756 159122 345808 159128
rect 345676 159066 345704 159122
rect 345676 159050 345888 159066
rect 345572 159044 345624 159050
rect 345676 159044 345900 159050
rect 345676 159038 345848 159044
rect 345572 158986 345624 158992
rect 345848 158986 345900 158992
rect 345216 157306 345336 157334
rect 345112 156800 345164 156806
rect 345112 156742 345164 156748
rect 344376 155712 344428 155718
rect 344376 155654 344428 155660
rect 343916 152992 343968 152998
rect 343916 152934 343968 152940
rect 343824 152380 343876 152386
rect 343824 152322 343876 152328
rect 342364 151786 342484 151814
rect 342548 151786 343312 151814
rect 342456 150226 342484 151786
rect 343284 150226 343312 151786
rect 343928 150226 343956 152934
rect 344560 152244 344612 152250
rect 344560 152186 344612 152192
rect 344572 150226 344600 152186
rect 333750 150146 333802 150152
rect 333762 149940 333790 150146
rect 334406 149940 334434 150198
rect 334958 149940 334986 150198
rect 335602 149940 335630 150198
rect 336246 149940 336274 150198
rect 336890 149940 336918 150198
rect 337534 149940 337562 150198
rect 338178 149940 338206 150198
rect 338304 150204 338356 150210
rect 338776 150198 338850 150226
rect 338304 150146 338356 150152
rect 338822 149940 338850 150198
rect 339454 150204 339506 150210
rect 339972 150198 340138 150226
rect 340708 150198 340782 150226
rect 341352 150198 341426 150226
rect 341996 150198 342070 150226
rect 342456 150198 342714 150226
rect 343284 150198 343358 150226
rect 343928 150198 344002 150226
rect 344572 150198 344646 150226
rect 345124 150210 345152 156742
rect 345204 155916 345256 155922
rect 345204 155858 345256 155864
rect 345216 150226 345244 155858
rect 345308 152998 345336 157306
rect 346412 154426 346440 163254
rect 346780 163146 346808 163254
rect 346858 163200 346914 164400
rect 347778 163200 347834 164400
rect 348160 163254 348556 163282
rect 346872 163146 346900 163200
rect 346780 163118 346900 163146
rect 347792 159730 347820 163200
rect 347780 159724 347832 159730
rect 347780 159666 347832 159672
rect 348056 156868 348108 156874
rect 348056 156810 348108 156816
rect 347872 155304 347924 155310
rect 347872 155246 347924 155252
rect 346400 154420 346452 154426
rect 346400 154362 346452 154368
rect 345296 152992 345348 152998
rect 345296 152934 345348 152940
rect 347136 152516 347188 152522
rect 347136 152458 347188 152464
rect 346492 151836 346544 151842
rect 346492 151778 346544 151784
rect 346504 150226 346532 151778
rect 347148 150226 347176 152458
rect 347884 150226 347912 155246
rect 348068 151814 348096 156810
rect 348160 152522 348188 163254
rect 348528 163146 348556 163254
rect 348606 163200 348662 164400
rect 349172 163254 349384 163282
rect 348620 163146 348648 163200
rect 348528 163118 348648 163146
rect 349068 159044 349120 159050
rect 349068 158986 349120 158992
rect 348148 152516 348200 152522
rect 348148 152458 348200 152464
rect 348068 151786 348464 151814
rect 339454 150146 339506 150152
rect 339466 149940 339494 150146
rect 340110 149940 340138 150198
rect 340754 149940 340782 150198
rect 341398 149940 341426 150198
rect 342042 149940 342070 150198
rect 342686 149940 342714 150198
rect 343330 149940 343358 150198
rect 343974 149940 344002 150198
rect 344618 149940 344646 150198
rect 345112 150204 345164 150210
rect 345216 150198 345290 150226
rect 345112 150146 345164 150152
rect 345262 149940 345290 150198
rect 345894 150204 345946 150210
rect 346504 150198 346578 150226
rect 347148 150198 347222 150226
rect 345894 150146 345946 150152
rect 345906 149940 345934 150146
rect 346550 149940 346578 150198
rect 347194 149940 347222 150198
rect 347838 150198 347912 150226
rect 348436 150226 348464 151786
rect 349080 150226 349108 158986
rect 349172 152250 349200 163254
rect 349356 163146 349384 163254
rect 349434 163200 349490 164400
rect 349540 163254 350212 163282
rect 349448 163146 349476 163200
rect 349356 163118 349476 163146
rect 349344 159452 349396 159458
rect 349344 159394 349396 159400
rect 349356 159118 349384 159394
rect 349252 159112 349304 159118
rect 349252 159054 349304 159060
rect 349344 159112 349396 159118
rect 349344 159054 349396 159060
rect 349160 152244 349212 152250
rect 349160 152186 349212 152192
rect 349264 151814 349292 159054
rect 349540 154494 349568 163254
rect 350184 163146 350212 163254
rect 350262 163200 350318 164400
rect 351090 163200 351146 164400
rect 351918 163200 351974 164400
rect 352024 163254 352696 163282
rect 350276 163146 350304 163200
rect 350184 163118 350304 163146
rect 351104 159050 351132 163200
rect 351932 159186 351960 163200
rect 351828 159180 351880 159186
rect 351828 159122 351880 159128
rect 351920 159180 351972 159186
rect 351920 159122 351972 159128
rect 351840 159066 351868 159122
rect 351092 159044 351144 159050
rect 351840 159038 351960 159066
rect 351092 158986 351144 158992
rect 350356 155100 350408 155106
rect 350356 155042 350408 155048
rect 349528 154488 349580 154494
rect 349528 154430 349580 154436
rect 349804 152380 349856 152386
rect 349804 152322 349856 152328
rect 349896 152380 349948 152386
rect 349896 152322 349948 152328
rect 349816 151842 349844 152322
rect 349908 152250 349936 152322
rect 349896 152244 349948 152250
rect 349896 152186 349948 152192
rect 349804 151836 349856 151842
rect 349264 151786 349752 151814
rect 349724 150226 349752 151786
rect 349804 151778 349856 151784
rect 350368 150226 350396 155042
rect 351932 152590 351960 159038
rect 351000 152584 351052 152590
rect 351000 152526 351052 152532
rect 351920 152584 351972 152590
rect 351920 152526 351972 152532
rect 351012 150226 351040 152526
rect 352024 152250 352052 163254
rect 352668 163146 352696 163254
rect 352746 163200 352802 164400
rect 353666 163200 353722 164400
rect 354494 163200 354550 164400
rect 354692 163254 355272 163282
rect 352760 163146 352788 163200
rect 352668 163118 352788 163146
rect 352472 155236 352524 155242
rect 352472 155178 352524 155184
rect 352012 152244 352064 152250
rect 352012 152186 352064 152192
rect 351644 152040 351696 152046
rect 351644 151982 351696 151988
rect 351656 150226 351684 151982
rect 352288 151972 352340 151978
rect 352288 151914 352340 151920
rect 352300 150226 352328 151914
rect 352484 151814 352512 155178
rect 353680 154562 353708 163200
rect 354220 159656 354272 159662
rect 354220 159598 354272 159604
rect 353668 154556 353720 154562
rect 353668 154498 353720 154504
rect 353484 152584 353536 152590
rect 353484 152526 353536 152532
rect 353496 151814 353524 152526
rect 352484 151786 352972 151814
rect 353496 151786 353616 151814
rect 352944 150226 352972 151786
rect 353588 150226 353616 151786
rect 354232 150226 354260 159598
rect 354508 152590 354536 163200
rect 354496 152584 354548 152590
rect 354496 152526 354548 152532
rect 354692 152046 354720 163254
rect 355244 163146 355272 163254
rect 355322 163200 355378 164400
rect 356150 163200 356206 164400
rect 356256 163254 356928 163282
rect 355336 163146 355364 163200
rect 355244 163118 355364 163146
rect 356164 159526 356192 163200
rect 354864 159520 354916 159526
rect 354864 159462 354916 159468
rect 356152 159520 356204 159526
rect 356152 159462 356204 159468
rect 354680 152040 354732 152046
rect 354680 151982 354732 151988
rect 354876 150226 354904 159462
rect 356256 153882 356284 163254
rect 356900 163146 356928 163254
rect 356978 163200 357034 164400
rect 357806 163200 357862 164400
rect 358634 163200 358690 164400
rect 358832 163254 359504 163282
rect 356992 163146 357020 163200
rect 356900 163118 357020 163146
rect 357820 159662 357848 163200
rect 357992 159792 358044 159798
rect 357992 159734 358044 159740
rect 357808 159656 357860 159662
rect 357808 159598 357860 159604
rect 357532 158976 357584 158982
rect 357532 158918 357584 158924
rect 355508 153876 355560 153882
rect 355508 153818 355560 153824
rect 356244 153876 356296 153882
rect 356244 153818 356296 153824
rect 355520 150226 355548 153818
rect 356152 152720 356204 152726
rect 356152 152662 356204 152668
rect 356164 150226 356192 152662
rect 357438 152416 357494 152425
rect 357438 152351 357494 152360
rect 356796 152176 356848 152182
rect 356796 152118 356848 152124
rect 356808 150226 356836 152118
rect 357452 150226 357480 152351
rect 357544 152182 357572 158918
rect 357900 153944 357952 153950
rect 357900 153886 357952 153892
rect 357532 152176 357584 152182
rect 357532 152118 357584 152124
rect 357912 150498 357940 153886
rect 358004 151814 358032 159734
rect 358648 159458 358676 163200
rect 358636 159452 358688 159458
rect 358636 159394 358688 159400
rect 358832 152726 358860 163254
rect 359476 163146 359504 163254
rect 359554 163200 359610 164400
rect 360382 163200 360438 164400
rect 361210 163200 361266 164400
rect 361592 163254 361988 163282
rect 359568 163146 359596 163200
rect 359476 163118 359596 163146
rect 358912 159588 358964 159594
rect 358912 159530 358964 159536
rect 358820 152720 358872 152726
rect 358820 152662 358872 152668
rect 358004 151786 358768 151814
rect 357912 150470 358124 150498
rect 358096 150226 358124 150470
rect 358740 150226 358768 151786
rect 348436 150198 348510 150226
rect 349080 150198 349154 150226
rect 349724 150198 349798 150226
rect 350368 150198 350442 150226
rect 351012 150198 351086 150226
rect 351656 150198 351730 150226
rect 352300 150198 352374 150226
rect 352944 150198 353018 150226
rect 353588 150198 353662 150226
rect 354232 150198 354306 150226
rect 354876 150198 354950 150226
rect 355520 150198 355594 150226
rect 356164 150198 356238 150226
rect 356808 150198 356882 150226
rect 357452 150198 357526 150226
rect 358096 150198 358170 150226
rect 358740 150198 358814 150226
rect 358924 150210 358952 159530
rect 360396 153814 360424 163200
rect 361224 158982 361252 163200
rect 361212 158976 361264 158982
rect 361212 158918 361264 158924
rect 360660 154012 360712 154018
rect 360660 153954 360712 153960
rect 360384 153808 360436 153814
rect 360384 153750 360436 153756
rect 359372 152176 359424 152182
rect 359372 152118 359424 152124
rect 359384 150226 359412 152118
rect 360672 150226 360700 153954
rect 361592 152794 361620 163254
rect 361960 163146 361988 163254
rect 362038 163200 362094 164400
rect 362866 163200 362922 164400
rect 363064 163254 363644 163282
rect 362052 163146 362080 163200
rect 361960 163118 362080 163146
rect 362880 159594 362908 163200
rect 362960 159860 363012 159866
rect 362960 159802 363012 159808
rect 362868 159588 362920 159594
rect 362868 159530 362920 159536
rect 361304 152788 361356 152794
rect 361304 152730 361356 152736
rect 361580 152788 361632 152794
rect 361580 152730 361632 152736
rect 361316 150226 361344 152730
rect 361948 152652 362000 152658
rect 361948 152594 362000 152600
rect 361960 150226 361988 152594
rect 362592 151904 362644 151910
rect 362592 151846 362644 151852
rect 362604 150226 362632 151846
rect 347838 149940 347866 150198
rect 348482 149940 348510 150198
rect 349126 149940 349154 150198
rect 349770 149940 349798 150198
rect 350414 149940 350442 150198
rect 351058 149940 351086 150198
rect 351702 149940 351730 150198
rect 352346 149940 352374 150198
rect 352990 149940 353018 150198
rect 353634 149940 353662 150198
rect 354278 149940 354306 150198
rect 354922 149940 354950 150198
rect 355566 149940 355594 150198
rect 356210 149940 356238 150198
rect 356854 149940 356882 150198
rect 357498 149940 357526 150198
rect 358142 149940 358170 150198
rect 358786 149940 358814 150198
rect 358912 150204 358964 150210
rect 359384 150198 359458 150226
rect 358912 150146 358964 150152
rect 359430 149940 359458 150198
rect 360062 150204 360114 150210
rect 360672 150198 360746 150226
rect 361316 150198 361390 150226
rect 361960 150198 362034 150226
rect 362604 150198 362678 150226
rect 362972 150210 363000 159802
rect 363064 153950 363092 163254
rect 363616 163146 363644 163254
rect 363694 163200 363750 164400
rect 364522 163200 364578 164400
rect 365442 163200 365498 164400
rect 365732 163254 366220 163282
rect 363708 163146 363736 163200
rect 363616 163118 363736 163146
rect 364536 161474 364564 163200
rect 364536 161446 364656 161474
rect 363144 158840 363196 158846
rect 363144 158782 363196 158788
rect 363052 153944 363104 153950
rect 363052 153886 363104 153892
rect 363156 151910 363184 158782
rect 363236 155372 363288 155378
rect 363236 155314 363288 155320
rect 363144 151904 363196 151910
rect 363144 151846 363196 151852
rect 363248 150226 363276 155314
rect 364628 151978 364656 161446
rect 365456 159798 365484 163200
rect 365444 159792 365496 159798
rect 365444 159734 365496 159740
rect 365168 158908 365220 158914
rect 365168 158850 365220 158856
rect 364616 151972 364668 151978
rect 364616 151914 364668 151920
rect 364524 151904 364576 151910
rect 364524 151846 364576 151852
rect 364536 150226 364564 151846
rect 365180 150226 365208 158850
rect 365732 152182 365760 163254
rect 366192 163146 366220 163254
rect 366270 163200 366326 164400
rect 367098 163200 367154 164400
rect 367926 163200 367982 164400
rect 368492 163254 368704 163282
rect 366284 163146 366312 163200
rect 366192 163118 366312 163146
rect 365812 154080 365864 154086
rect 365812 154022 365864 154028
rect 365720 152176 365772 152182
rect 365720 152118 365772 152124
rect 365824 150226 365852 154022
rect 367112 154018 367140 163200
rect 367940 158778 367968 163200
rect 367192 158772 367244 158778
rect 367192 158714 367244 158720
rect 367928 158772 367980 158778
rect 367928 158714 367980 158720
rect 367100 154012 367152 154018
rect 367100 153954 367152 153960
rect 367204 153134 367232 158714
rect 368296 154148 368348 154154
rect 368296 154090 368348 154096
rect 367008 153128 367060 153134
rect 367008 153070 367060 153076
rect 367192 153128 367244 153134
rect 367192 153070 367244 153076
rect 366364 152856 366416 152862
rect 366364 152798 366416 152804
rect 360062 150146 360114 150152
rect 360074 149940 360102 150146
rect 360718 149940 360746 150198
rect 361362 149940 361390 150198
rect 362006 149940 362034 150198
rect 362650 149940 362678 150198
rect 362960 150204 363012 150210
rect 363248 150198 363322 150226
rect 362960 150146 363012 150152
rect 363294 149940 363322 150198
rect 363926 150204 363978 150210
rect 364536 150198 364610 150226
rect 365180 150198 365254 150226
rect 363926 150146 363978 150152
rect 363938 149940 363966 150146
rect 364582 149940 364610 150198
rect 365226 149940 365254 150198
rect 365778 150198 365852 150226
rect 366376 150226 366404 152798
rect 367020 150226 367048 153070
rect 367652 152448 367704 152454
rect 367652 152390 367704 152396
rect 367664 150226 367692 152390
rect 368308 150226 368336 154090
rect 368492 152658 368520 163254
rect 368676 163146 368704 163254
rect 368754 163200 368810 164400
rect 369582 163200 369638 164400
rect 370410 163200 370466 164400
rect 371330 163200 371386 164400
rect 372158 163200 372214 164400
rect 372632 163254 372936 163282
rect 368768 163146 368796 163200
rect 368676 163118 368796 163146
rect 369492 159928 369544 159934
rect 369492 159870 369544 159876
rect 369216 159656 369268 159662
rect 369216 159598 369268 159604
rect 369228 158982 369256 159598
rect 369216 158976 369268 158982
rect 369216 158918 369268 158924
rect 368940 153128 368992 153134
rect 368940 153070 368992 153076
rect 368480 152652 368532 152658
rect 368480 152594 368532 152600
rect 368952 150226 368980 153070
rect 369504 151814 369532 159870
rect 369596 159662 369624 163200
rect 369952 159996 370004 160002
rect 369952 159938 370004 159944
rect 369584 159656 369636 159662
rect 369584 159598 369636 159604
rect 369964 151814 369992 159938
rect 370424 155242 370452 163200
rect 370872 155440 370924 155446
rect 370872 155382 370924 155388
rect 370412 155236 370464 155242
rect 370412 155178 370464 155184
rect 369504 151786 369624 151814
rect 369964 151786 370268 151814
rect 369596 150226 369624 151786
rect 370240 150226 370268 151786
rect 370884 150226 370912 155382
rect 371344 152862 371372 163200
rect 372172 159934 372200 163200
rect 372160 159928 372212 159934
rect 372160 159870 372212 159876
rect 372632 153066 372660 163254
rect 372908 163146 372936 163254
rect 372986 163200 373042 164400
rect 373814 163200 373870 164400
rect 374642 163200 374698 164400
rect 375470 163200 375526 164400
rect 376298 163200 376354 164400
rect 376864 163254 377168 163282
rect 373000 163146 373028 163200
rect 372908 163118 373028 163146
rect 373448 155508 373500 155514
rect 373448 155450 373500 155456
rect 371516 153060 371568 153066
rect 371516 153002 371568 153008
rect 372620 153060 372672 153066
rect 372620 153002 372672 153008
rect 371332 152856 371384 152862
rect 371332 152798 371384 152804
rect 371528 150226 371556 153002
rect 372804 152924 372856 152930
rect 372804 152866 372856 152872
rect 372160 152312 372212 152318
rect 372160 152254 372212 152260
rect 372172 150226 372200 152254
rect 372816 150226 372844 152866
rect 373460 150226 373488 155450
rect 373828 155310 373856 163200
rect 374092 160064 374144 160070
rect 374092 160006 374144 160012
rect 374000 159316 374052 159322
rect 374000 159258 374052 159264
rect 373816 155304 373868 155310
rect 373816 155246 373868 155252
rect 366376 150198 366450 150226
rect 367020 150198 367094 150226
rect 367664 150198 367738 150226
rect 368308 150198 368382 150226
rect 368952 150198 369026 150226
rect 369596 150198 369670 150226
rect 370240 150198 370314 150226
rect 370884 150198 370958 150226
rect 371528 150198 371602 150226
rect 372172 150198 372246 150226
rect 372816 150198 372890 150226
rect 373460 150198 373534 150226
rect 374012 150210 374040 159258
rect 374104 150226 374132 160006
rect 374656 160002 374684 163200
rect 374644 159996 374696 160002
rect 374644 159938 374696 159944
rect 374644 159316 374696 159322
rect 374644 159258 374696 159264
rect 374656 159050 374684 159258
rect 374644 159044 374696 159050
rect 374644 158986 374696 158992
rect 374552 158840 374604 158846
rect 374736 158840 374788 158846
rect 374604 158788 374736 158794
rect 374552 158782 374788 158788
rect 374564 158766 374776 158782
rect 375484 152930 375512 163200
rect 376312 159866 376340 163200
rect 376300 159860 376352 159866
rect 376300 159802 376352 159808
rect 375564 155576 375616 155582
rect 375564 155518 375616 155524
rect 375472 152924 375524 152930
rect 375472 152866 375524 152872
rect 375380 152108 375432 152114
rect 375380 152050 375432 152056
rect 375392 150226 375420 152050
rect 365778 149940 365806 150198
rect 366422 149940 366450 150198
rect 367066 149940 367094 150198
rect 367710 149940 367738 150198
rect 368354 149940 368382 150198
rect 368998 149940 369026 150198
rect 369642 149940 369670 150198
rect 370286 149940 370314 150198
rect 370930 149940 370958 150198
rect 371574 149940 371602 150198
rect 372218 149940 372246 150198
rect 372862 149940 372890 150198
rect 373506 149940 373534 150198
rect 374000 150204 374052 150210
rect 374104 150198 374178 150226
rect 374000 150146 374052 150152
rect 374150 149940 374178 150198
rect 374782 150204 374834 150210
rect 375392 150198 375466 150226
rect 375576 150210 375604 155518
rect 376024 154216 376076 154222
rect 376024 154158 376076 154164
rect 376036 150226 376064 154158
rect 376864 154154 376892 163254
rect 377140 163146 377168 163254
rect 377218 163200 377274 164400
rect 378046 163200 378102 164400
rect 378874 163200 378930 164400
rect 379702 163200 379758 164400
rect 380176 163254 380480 163282
rect 377232 163146 377260 163200
rect 377140 163118 377260 163146
rect 377956 159248 378008 159254
rect 377956 159190 378008 159196
rect 376852 154148 376904 154154
rect 376852 154090 376904 154096
rect 377312 153196 377364 153202
rect 377312 153138 377364 153144
rect 377324 150226 377352 153138
rect 377968 150226 377996 159190
rect 378060 159118 378088 163200
rect 378888 160070 378916 163200
rect 378876 160064 378928 160070
rect 378876 160006 378928 160012
rect 379716 159730 379744 163200
rect 378784 159724 378836 159730
rect 378784 159666 378836 159672
rect 379704 159724 379756 159730
rect 379704 159666 379756 159672
rect 378048 159112 378100 159118
rect 378048 159054 378100 159060
rect 378232 159044 378284 159050
rect 378232 158986 378284 158992
rect 378140 155644 378192 155650
rect 378140 155586 378192 155592
rect 374782 150146 374834 150152
rect 374794 149940 374822 150146
rect 375438 149940 375466 150198
rect 375564 150204 375616 150210
rect 376036 150198 376110 150226
rect 375564 150146 375616 150152
rect 376082 149940 376110 150198
rect 376714 150204 376766 150210
rect 377324 150198 377398 150226
rect 377968 150198 378042 150226
rect 378152 150210 378180 155586
rect 378244 153202 378272 158986
rect 378600 154284 378652 154290
rect 378600 154226 378652 154232
rect 378232 153196 378284 153202
rect 378232 153138 378284 153144
rect 378612 150226 378640 154226
rect 378796 152114 378824 159666
rect 380176 154086 380204 163254
rect 380452 163146 380480 163254
rect 380530 163200 380586 164400
rect 381004 163254 381308 163282
rect 380544 163146 380572 163200
rect 380452 163118 380572 163146
rect 380164 154080 380216 154086
rect 380164 154022 380216 154028
rect 379888 153196 379940 153202
rect 379888 153138 379940 153144
rect 378784 152108 378836 152114
rect 378784 152050 378836 152056
rect 379900 150226 379928 153138
rect 381004 152454 381032 163254
rect 381280 163146 381308 163254
rect 381358 163200 381414 164400
rect 382186 163200 382242 164400
rect 383106 163200 383162 164400
rect 383672 163254 383884 163282
rect 381372 163146 381400 163200
rect 381280 163118 381400 163146
rect 381820 155712 381872 155718
rect 381820 155654 381872 155660
rect 381176 154352 381228 154358
rect 381176 154294 381228 154300
rect 380992 152448 381044 152454
rect 380992 152390 381044 152396
rect 380532 151836 380584 151842
rect 380532 151778 380584 151784
rect 380544 150226 380572 151778
rect 381188 150226 381216 154294
rect 381832 150226 381860 155654
rect 382200 153134 382228 163200
rect 383120 159390 383148 163200
rect 382832 159384 382884 159390
rect 382832 159326 382884 159332
rect 383108 159384 383160 159390
rect 383108 159326 383160 159332
rect 382280 159316 382332 159322
rect 382280 159258 382332 159264
rect 382188 153128 382240 153134
rect 382188 153070 382240 153076
rect 382292 152318 382320 159258
rect 382464 152992 382516 152998
rect 382464 152934 382516 152940
rect 382280 152312 382332 152318
rect 382280 152254 382332 152260
rect 382476 150226 382504 152934
rect 382844 151814 382872 159326
rect 383672 154222 383700 163254
rect 383856 163146 383884 163254
rect 383934 163200 383990 164400
rect 384762 163200 384818 164400
rect 385590 163200 385646 164400
rect 386418 163200 386474 164400
rect 386524 163254 387196 163282
rect 383948 163146 383976 163200
rect 383856 163118 383976 163146
rect 384776 158846 384804 163200
rect 385604 159254 385632 163200
rect 385500 159248 385552 159254
rect 385500 159190 385552 159196
rect 385592 159248 385644 159254
rect 385592 159190 385644 159196
rect 384948 158976 385000 158982
rect 384948 158918 385000 158924
rect 384764 158840 384816 158846
rect 384764 158782 384816 158788
rect 383752 154420 383804 154426
rect 383752 154362 383804 154368
rect 383660 154216 383712 154222
rect 383660 154158 383712 154164
rect 382844 151786 383148 151814
rect 383120 150226 383148 151786
rect 383764 150226 383792 154362
rect 384960 152998 384988 158918
rect 385512 153202 385540 159190
rect 386144 158908 386196 158914
rect 386144 158850 386196 158856
rect 385500 153196 385552 153202
rect 385500 153138 385552 153144
rect 384948 152992 385000 152998
rect 384948 152934 385000 152940
rect 385040 152516 385092 152522
rect 385040 152458 385092 152464
rect 384396 152108 384448 152114
rect 384396 152050 384448 152056
rect 384408 150226 384436 152050
rect 385052 150226 385080 152458
rect 385684 152380 385736 152386
rect 385684 152322 385736 152328
rect 385696 150226 385724 152322
rect 386156 151842 386184 158850
rect 386236 158772 386288 158778
rect 386236 158714 386288 158720
rect 386248 152386 386276 158714
rect 386328 154488 386380 154494
rect 386328 154430 386380 154436
rect 386236 152380 386288 152386
rect 386236 152322 386288 152328
rect 386144 151836 386196 151842
rect 386144 151778 386196 151784
rect 386340 150226 386368 154430
rect 386432 152522 386460 163200
rect 386524 154290 386552 163254
rect 387168 163146 387196 163254
rect 387246 163200 387302 164400
rect 388074 163200 388130 164400
rect 388994 163200 389050 164400
rect 389822 163200 389878 164400
rect 390650 163200 390706 164400
rect 391478 163200 391534 164400
rect 392306 163200 392362 164400
rect 393134 163200 393190 164400
rect 393332 163254 393912 163282
rect 387260 163146 387288 163200
rect 387168 163118 387288 163146
rect 388088 158778 388116 163200
rect 388168 159996 388220 160002
rect 388168 159938 388220 159944
rect 388076 158772 388128 158778
rect 388076 158714 388128 158720
rect 386512 154284 386564 154290
rect 386512 154226 386564 154232
rect 387616 153196 387668 153202
rect 387616 153138 387668 153144
rect 386420 152516 386472 152522
rect 386420 152458 386472 152464
rect 386972 152312 387024 152318
rect 386972 152254 387024 152260
rect 386984 150226 387012 152254
rect 387628 150226 387656 153138
rect 388180 151910 388208 159938
rect 389008 159322 389036 163200
rect 389836 160002 389864 163200
rect 389824 159996 389876 160002
rect 389824 159938 389876 159944
rect 390560 159520 390612 159526
rect 390560 159462 390612 159468
rect 388996 159316 389048 159322
rect 388996 159258 389048 159264
rect 388444 159180 388496 159186
rect 388444 159122 388496 159128
rect 388260 152244 388312 152250
rect 388260 152186 388312 152192
rect 388168 151904 388220 151910
rect 388168 151846 388220 151852
rect 388272 150226 388300 152186
rect 388456 152114 388484 159122
rect 389180 158840 389232 158846
rect 389180 158782 389232 158788
rect 388904 154556 388956 154562
rect 388904 154498 388956 154504
rect 388444 152108 388496 152114
rect 388444 152050 388496 152056
rect 388916 150226 388944 154498
rect 389192 153202 389220 158782
rect 390376 158772 390428 158778
rect 390376 158714 390428 158720
rect 389180 153196 389232 153202
rect 389180 153138 389232 153144
rect 390388 152590 390416 158714
rect 389548 152584 389600 152590
rect 389548 152526 389600 152532
rect 390376 152584 390428 152590
rect 390376 152526 390428 152532
rect 376714 150146 376766 150152
rect 376726 149940 376754 150146
rect 377370 149940 377398 150198
rect 378014 149940 378042 150198
rect 378140 150204 378192 150210
rect 378612 150198 378686 150226
rect 378140 150146 378192 150152
rect 378658 149940 378686 150198
rect 379290 150204 379342 150210
rect 379900 150198 379974 150226
rect 380544 150198 380618 150226
rect 381188 150198 381262 150226
rect 381832 150198 381906 150226
rect 382476 150198 382550 150226
rect 383120 150198 383194 150226
rect 383764 150198 383838 150226
rect 384408 150198 384482 150226
rect 385052 150198 385126 150226
rect 385696 150198 385770 150226
rect 386340 150198 386414 150226
rect 386984 150198 387058 150226
rect 387628 150198 387702 150226
rect 388272 150198 388346 150226
rect 388916 150198 388990 150226
rect 379290 150146 379342 150152
rect 379302 149940 379330 150146
rect 379946 149940 379974 150198
rect 380590 149940 380618 150198
rect 381234 149940 381262 150198
rect 381878 149940 381906 150198
rect 382522 149940 382550 150198
rect 383166 149940 383194 150198
rect 383810 149940 383838 150198
rect 384454 149940 384482 150198
rect 385098 149940 385126 150198
rect 385742 149940 385770 150198
rect 386386 149940 386414 150198
rect 387030 149940 387058 150198
rect 387674 149940 387702 150198
rect 388318 149940 388346 150198
rect 388962 149940 388990 150198
rect 389560 150090 389588 152526
rect 390192 152040 390244 152046
rect 390192 151982 390244 151988
rect 390204 150090 390232 151982
rect 390572 150226 390600 159462
rect 390664 154494 390692 163200
rect 391492 158914 391520 163200
rect 392320 159186 392348 163200
rect 392768 159452 392820 159458
rect 392768 159394 392820 159400
rect 392308 159180 392360 159186
rect 392308 159122 392360 159128
rect 391480 158908 391532 158914
rect 391480 158850 391532 158856
rect 390652 154488 390704 154494
rect 390652 154430 390704 154436
rect 391480 153876 391532 153882
rect 391480 153818 391532 153824
rect 390572 150198 390922 150226
rect 389560 150062 389634 150090
rect 390204 150062 390278 150090
rect 389606 149940 389634 150062
rect 390250 149940 390278 150062
rect 390894 149940 390922 150198
rect 391492 150090 391520 153818
rect 392124 152992 392176 152998
rect 392124 152934 392176 152940
rect 392136 150090 392164 152934
rect 392780 150226 392808 159394
rect 393148 152318 393176 163200
rect 393332 154358 393360 163254
rect 393884 163146 393912 163254
rect 393962 163200 394018 164400
rect 394882 163200 394938 164400
rect 395710 163200 395766 164400
rect 396538 163200 396594 164400
rect 397366 163200 397422 164400
rect 397472 163254 398144 163282
rect 393976 163146 394004 163200
rect 393884 163118 394004 163146
rect 394332 158908 394384 158914
rect 394332 158850 394384 158856
rect 393320 154352 393372 154358
rect 393320 154294 393372 154300
rect 394056 153808 394108 153814
rect 394056 153750 394108 153756
rect 393504 153196 393556 153202
rect 393504 153138 393556 153144
rect 393516 152726 393544 153138
rect 393412 152720 393464 152726
rect 393412 152662 393464 152668
rect 393504 152720 393556 152726
rect 393504 152662 393556 152668
rect 393136 152312 393188 152318
rect 393136 152254 393188 152260
rect 392780 150198 392854 150226
rect 391492 150062 391566 150090
rect 392136 150062 392210 150090
rect 391538 149940 391566 150062
rect 392182 149940 392210 150062
rect 392826 149940 392854 150198
rect 393424 150090 393452 152662
rect 394068 150090 394096 153750
rect 394344 152250 394372 158850
rect 394896 152998 394924 163200
rect 395528 159792 395580 159798
rect 395528 159734 395580 159740
rect 394976 159588 395028 159594
rect 394976 159530 395028 159536
rect 394988 157334 395016 159530
rect 394988 157306 395476 157334
rect 394884 152992 394936 152998
rect 394884 152934 394936 152940
rect 395344 152788 395396 152794
rect 395344 152730 395396 152736
rect 394332 152244 394384 152250
rect 394332 152186 394384 152192
rect 394700 151836 394752 151842
rect 394700 151778 394752 151784
rect 394712 150090 394740 151778
rect 395356 150090 395384 152730
rect 395448 152538 395476 157306
rect 395540 153202 395568 159734
rect 395724 159118 395752 163200
rect 396172 159928 396224 159934
rect 396172 159870 396224 159876
rect 395712 159112 395764 159118
rect 395712 159054 395764 159060
rect 395528 153196 395580 153202
rect 395528 153138 395580 153144
rect 395448 152510 396028 152538
rect 396000 150226 396028 152510
rect 396184 151910 396212 159870
rect 396552 159798 396580 163200
rect 396540 159792 396592 159798
rect 396540 159734 396592 159740
rect 397380 154426 397408 163200
rect 397368 154420 397420 154426
rect 397368 154362 397420 154368
rect 396540 153944 396592 153950
rect 396540 153886 396592 153892
rect 396172 151904 396224 151910
rect 396172 151846 396224 151852
rect 396000 150198 396074 150226
rect 393424 150062 393498 150090
rect 394068 150062 394142 150090
rect 394712 150062 394786 150090
rect 395356 150062 395430 150090
rect 393470 149940 393498 150062
rect 394114 149940 394142 150062
rect 394758 149940 394786 150062
rect 395402 149940 395430 150062
rect 396046 149940 396074 150198
rect 396552 150090 396580 153886
rect 397472 153882 397500 163254
rect 398116 163146 398144 163254
rect 398194 163200 398250 164400
rect 399022 163200 399078 164400
rect 399128 163254 399800 163282
rect 398208 163146 398236 163200
rect 398116 163118 398236 163146
rect 398564 160064 398616 160070
rect 398564 160006 398616 160012
rect 397460 153876 397512 153882
rect 397460 153818 397512 153824
rect 397828 153196 397880 153202
rect 397828 153138 397880 153144
rect 397920 153196 397972 153202
rect 397920 153138 397972 153144
rect 397184 152040 397236 152046
rect 397184 151982 397236 151988
rect 397196 150090 397224 151982
rect 397840 150090 397868 153138
rect 397932 152590 397960 153138
rect 398104 152720 398156 152726
rect 398104 152662 398156 152668
rect 397920 152584 397972 152590
rect 397920 152526 397972 152532
rect 398012 152584 398064 152590
rect 398012 152526 398064 152532
rect 398024 152318 398052 152526
rect 398116 152318 398144 152662
rect 398012 152312 398064 152318
rect 398012 152254 398064 152260
rect 398104 152312 398156 152318
rect 398104 152254 398156 152260
rect 398576 152182 398604 160006
rect 399036 159594 399064 163200
rect 399024 159588 399076 159594
rect 399024 159530 399076 159536
rect 398840 159248 398892 159254
rect 398840 159190 398892 159196
rect 398852 152794 398880 159190
rect 399128 157334 399156 163254
rect 399772 163146 399800 163254
rect 399850 163200 399906 164400
rect 400770 163200 400826 164400
rect 401598 163200 401654 164400
rect 402426 163200 402482 164400
rect 403254 163200 403310 164400
rect 404082 163200 404138 164400
rect 404372 163254 404860 163282
rect 399864 163146 399892 163200
rect 399772 163118 399892 163146
rect 400784 159526 400812 163200
rect 401048 159656 401100 159662
rect 401048 159598 401100 159604
rect 400772 159520 400824 159526
rect 400772 159462 400824 159468
rect 399128 157306 399248 157334
rect 399116 154012 399168 154018
rect 399116 153954 399168 153960
rect 398840 152788 398892 152794
rect 398840 152730 398892 152736
rect 398472 152176 398524 152182
rect 398472 152118 398524 152124
rect 398564 152176 398616 152182
rect 398564 152118 398616 152124
rect 398484 150090 398512 152118
rect 399128 150090 399156 153954
rect 399220 152726 399248 157306
rect 399208 152720 399260 152726
rect 399208 152662 399260 152668
rect 400404 152652 400456 152658
rect 400404 152594 400456 152600
rect 399760 152380 399812 152386
rect 399760 152322 399812 152328
rect 399772 150090 399800 152322
rect 400416 150090 400444 152594
rect 401060 150226 401088 159598
rect 401612 153950 401640 163200
rect 401692 155236 401744 155242
rect 401692 155178 401744 155184
rect 401600 153944 401652 153950
rect 401600 153886 401652 153892
rect 401060 150198 401134 150226
rect 396552 150062 396626 150090
rect 397196 150062 397270 150090
rect 397840 150062 397914 150090
rect 398484 150062 398558 150090
rect 399128 150062 399202 150090
rect 399772 150062 399846 150090
rect 400416 150062 400490 150090
rect 396598 149940 396626 150062
rect 397242 149940 397270 150062
rect 397886 149940 397914 150062
rect 398530 149940 398558 150062
rect 399174 149940 399202 150062
rect 399818 149940 399846 150062
rect 400462 149940 400490 150062
rect 401106 149940 401134 150198
rect 401704 150090 401732 155178
rect 402336 152856 402388 152862
rect 402336 152798 402388 152804
rect 402348 150090 402376 152798
rect 402440 152386 402468 163200
rect 403268 159934 403296 163200
rect 403256 159928 403308 159934
rect 403256 159870 403308 159876
rect 404096 159458 404124 163200
rect 404084 159452 404136 159458
rect 404084 159394 404136 159400
rect 404268 159316 404320 159322
rect 404268 159258 404320 159264
rect 404176 159180 404228 159186
rect 404176 159122 404228 159128
rect 404084 155304 404136 155310
rect 404084 155246 404136 155252
rect 403624 153060 403676 153066
rect 403624 153002 403676 153008
rect 403348 152584 403400 152590
rect 403532 152584 403584 152590
rect 403400 152532 403532 152538
rect 403348 152526 403584 152532
rect 403360 152510 403572 152526
rect 402428 152380 402480 152386
rect 402428 152322 402480 152328
rect 402980 151904 403032 151910
rect 402980 151846 403032 151852
rect 402992 150090 403020 151846
rect 403636 150090 403664 153002
rect 403808 152788 403860 152794
rect 403808 152730 403860 152736
rect 403716 152448 403768 152454
rect 403716 152390 403768 152396
rect 403728 152318 403756 152390
rect 403820 152318 403848 152730
rect 403716 152312 403768 152318
rect 403716 152254 403768 152260
rect 403808 152312 403860 152318
rect 403808 152254 403860 152260
rect 404096 150226 404124 155246
rect 404188 151978 404216 159122
rect 404176 151972 404228 151978
rect 404176 151914 404228 151920
rect 404280 151842 404308 159258
rect 404372 152794 404400 163254
rect 404832 163146 404860 163254
rect 404910 163200 404966 164400
rect 405738 163200 405794 164400
rect 406658 163200 406714 164400
rect 407486 163200 407542 164400
rect 407684 163254 408264 163282
rect 404924 163146 404952 163200
rect 404832 163118 404952 163146
rect 405752 159118 405780 163200
rect 406200 159860 406252 159866
rect 406200 159802 406252 159808
rect 405832 159724 405884 159730
rect 405832 159666 405884 159672
rect 405372 159112 405424 159118
rect 405372 159054 405424 159060
rect 405740 159112 405792 159118
rect 405740 159054 405792 159060
rect 404360 152788 404412 152794
rect 404360 152730 404412 152736
rect 405384 152046 405412 159054
rect 405844 153066 405872 159666
rect 405832 153060 405884 153066
rect 405832 153002 405884 153008
rect 405556 152924 405608 152930
rect 405556 152866 405608 152872
rect 404912 152040 404964 152046
rect 404912 151982 404964 151988
rect 405372 152040 405424 152046
rect 405372 151982 405424 151988
rect 404268 151836 404320 151842
rect 404268 151778 404320 151784
rect 404096 150198 404354 150226
rect 401704 150062 401778 150090
rect 402348 150062 402422 150090
rect 402992 150062 403066 150090
rect 403636 150062 403710 150090
rect 401750 149940 401778 150062
rect 402394 149940 402422 150062
rect 403038 149940 403066 150062
rect 403682 149940 403710 150062
rect 404326 149940 404354 150198
rect 404924 150090 404952 151982
rect 405568 150090 405596 152866
rect 406212 150226 406240 159802
rect 406672 152930 406700 163200
rect 407500 159662 407528 163200
rect 407488 159656 407540 159662
rect 407488 159598 407540 159604
rect 406844 154148 406896 154154
rect 406844 154090 406896 154096
rect 406660 152924 406712 152930
rect 406660 152866 406712 152872
rect 406212 150198 406286 150226
rect 404924 150062 404998 150090
rect 405568 150062 405642 150090
rect 404970 149940 404998 150062
rect 405614 149940 405642 150062
rect 406258 149940 406286 150198
rect 406856 150090 406884 154090
rect 407684 152425 407712 163254
rect 408236 163146 408264 163254
rect 408314 163200 408370 164400
rect 409142 163200 409198 164400
rect 409970 163200 410026 164400
rect 410798 163200 410854 164400
rect 411272 163254 411576 163282
rect 408328 163146 408356 163200
rect 408236 163118 408356 163146
rect 408500 159588 408552 159594
rect 408500 159530 408552 159536
rect 407670 152416 407726 152425
rect 407670 152351 407726 152360
rect 408132 152176 408184 152182
rect 408132 152118 408184 152124
rect 407488 152108 407540 152114
rect 407488 152050 407540 152056
rect 407500 150090 407528 152050
rect 408144 150090 408172 152118
rect 408512 152114 408540 159530
rect 409156 158778 409184 163200
rect 409984 159866 410012 163200
rect 409972 159860 410024 159866
rect 409972 159802 410024 159808
rect 410812 159594 410840 163200
rect 410800 159588 410852 159594
rect 410800 159530 410852 159536
rect 409236 159112 409288 159118
rect 409236 159054 409288 159060
rect 409144 158772 409196 158778
rect 409144 158714 409196 158720
rect 408776 153060 408828 153066
rect 408776 153002 408828 153008
rect 408500 152108 408552 152114
rect 408500 152050 408552 152056
rect 408788 150226 408816 153002
rect 409248 152182 409276 159054
rect 410524 158772 410576 158778
rect 410524 158714 410576 158720
rect 409420 154080 409472 154086
rect 409420 154022 409472 154028
rect 409236 152176 409288 152182
rect 409236 152118 409288 152124
rect 409432 150226 409460 154022
rect 410536 153066 410564 158714
rect 410708 153128 410760 153134
rect 410708 153070 410760 153076
rect 410524 153060 410576 153066
rect 410524 153002 410576 153008
rect 410064 152516 410116 152522
rect 410064 152458 410116 152464
rect 410076 150226 410104 152458
rect 410720 150226 410748 153070
rect 411272 152862 411300 163254
rect 411548 163146 411576 163254
rect 411626 163200 411682 164400
rect 412546 163200 412602 164400
rect 413374 163200 413430 164400
rect 414202 163200 414258 164400
rect 414308 163254 414980 163282
rect 411640 163146 411668 163200
rect 411548 163118 411668 163146
rect 411352 159384 411404 159390
rect 411352 159326 411404 159332
rect 411260 152856 411312 152862
rect 411260 152798 411312 152804
rect 411364 150226 411392 159326
rect 412560 158914 412588 163200
rect 412548 158908 412600 158914
rect 412548 158850 412600 158856
rect 412916 158908 412968 158914
rect 412916 158850 412968 158856
rect 411996 154216 412048 154222
rect 411996 154158 412048 154164
rect 412008 150226 412036 154158
rect 412928 153134 412956 158850
rect 413388 158778 413416 163200
rect 413836 159996 413888 160002
rect 413836 159938 413888 159944
rect 413376 158772 413428 158778
rect 413376 158714 413428 158720
rect 412916 153128 412968 153134
rect 412916 153070 412968 153076
rect 413848 152522 413876 159938
rect 413928 159792 413980 159798
rect 413928 159734 413980 159740
rect 413940 152810 413968 159734
rect 414216 159390 414244 163200
rect 414204 159384 414256 159390
rect 414204 159326 414256 159332
rect 413940 152782 414060 152810
rect 414032 152658 414060 152782
rect 413928 152652 413980 152658
rect 413928 152594 413980 152600
rect 414020 152652 414072 152658
rect 414020 152594 414072 152600
rect 413836 152516 413888 152522
rect 413836 152458 413888 152464
rect 412640 152448 412692 152454
rect 412640 152390 412692 152396
rect 412652 150226 412680 152390
rect 413284 152312 413336 152318
rect 413284 152254 413336 152260
rect 413296 150226 413324 152254
rect 413940 150226 413968 152594
rect 414308 152318 414336 163254
rect 414952 163146 414980 163254
rect 415030 163200 415086 164400
rect 415412 163254 415808 163282
rect 415044 163146 415072 163200
rect 414952 163118 415072 163146
rect 414572 154284 414624 154290
rect 414572 154226 414624 154232
rect 414296 152312 414348 152318
rect 414296 152254 414348 152260
rect 414584 150226 414612 154226
rect 415216 153196 415268 153202
rect 415216 153138 415268 153144
rect 415228 150226 415256 153138
rect 415412 152998 415440 163254
rect 415780 163146 415808 163254
rect 415858 163200 415914 164400
rect 416686 163200 416742 164400
rect 417514 163200 417570 164400
rect 418172 163254 418384 163282
rect 415872 163146 415900 163200
rect 415780 163118 415900 163146
rect 416596 159928 416648 159934
rect 416596 159870 416648 159876
rect 415308 152992 415360 152998
rect 415308 152934 415360 152940
rect 415400 152992 415452 152998
rect 415400 152934 415452 152940
rect 415320 152454 415348 152934
rect 416504 152516 416556 152522
rect 416504 152458 416556 152464
rect 415308 152448 415360 152454
rect 415308 152390 415360 152396
rect 415860 151836 415912 151842
rect 415860 151778 415912 151784
rect 415872 150226 415900 151778
rect 416516 150226 416544 152458
rect 416608 151910 416636 159870
rect 416700 158982 416728 163200
rect 417528 159730 417556 163200
rect 417884 159860 417936 159866
rect 417884 159802 417936 159808
rect 417516 159724 417568 159730
rect 417516 159666 417568 159672
rect 416688 158976 416740 158982
rect 416688 158918 416740 158924
rect 417148 154488 417200 154494
rect 417148 154430 417200 154436
rect 416596 151904 416648 151910
rect 416596 151846 416648 151852
rect 417160 150226 417188 154430
rect 417608 152924 417660 152930
rect 417608 152866 417660 152872
rect 417332 152720 417384 152726
rect 417332 152662 417384 152668
rect 417344 151842 417372 152662
rect 417620 152658 417648 152866
rect 417608 152652 417660 152658
rect 417608 152594 417660 152600
rect 417896 152250 417924 159802
rect 418172 153202 418200 163254
rect 418356 163146 418384 163254
rect 418434 163200 418490 164400
rect 418632 163254 419212 163282
rect 418448 163146 418476 163200
rect 418356 163118 418476 163146
rect 418160 153196 418212 153202
rect 418160 153138 418212 153144
rect 418632 152522 418660 163254
rect 419184 163146 419212 163254
rect 419262 163200 419318 164400
rect 420090 163200 420146 164400
rect 420918 163200 420974 164400
rect 421024 163254 421696 163282
rect 419276 163146 419304 163200
rect 419184 163118 419304 163146
rect 419540 158976 419592 158982
rect 419540 158918 419592 158924
rect 419080 152584 419132 152590
rect 419080 152526 419132 152532
rect 418620 152516 418672 152522
rect 418620 152458 418672 152464
rect 417792 152244 417844 152250
rect 417792 152186 417844 152192
rect 417884 152244 417936 152250
rect 417884 152186 417936 152192
rect 417332 151836 417384 151842
rect 417332 151778 417384 151784
rect 417804 150226 417832 152186
rect 418436 151972 418488 151978
rect 418436 151914 418488 151920
rect 408788 150198 408862 150226
rect 409432 150198 409506 150226
rect 410076 150198 410150 150226
rect 410720 150198 410794 150226
rect 411364 150198 411438 150226
rect 412008 150198 412082 150226
rect 412652 150198 412726 150226
rect 413296 150198 413370 150226
rect 413940 150198 414014 150226
rect 414584 150198 414658 150226
rect 415228 150198 415302 150226
rect 415872 150198 415946 150226
rect 416516 150198 416590 150226
rect 417160 150198 417234 150226
rect 417804 150198 417878 150226
rect 406856 150062 406930 150090
rect 407500 150062 407574 150090
rect 408144 150062 408218 150090
rect 406902 149940 406930 150062
rect 407546 149940 407574 150062
rect 408190 149940 408218 150062
rect 408834 149940 408862 150198
rect 409478 149940 409506 150198
rect 410122 149940 410150 150198
rect 410766 149940 410794 150198
rect 411410 149940 411438 150198
rect 412054 149940 412082 150198
rect 412698 149940 412726 150198
rect 413342 149940 413370 150198
rect 413986 149940 414014 150198
rect 414630 149940 414658 150198
rect 415274 149940 415302 150198
rect 415918 149940 415946 150198
rect 416562 149940 416590 150198
rect 417206 149940 417234 150198
rect 417850 149940 417878 150198
rect 418448 150090 418476 151914
rect 419092 150090 419120 152526
rect 419552 152522 419580 158918
rect 420104 158914 420132 163200
rect 420932 159798 420960 163200
rect 420920 159792 420972 159798
rect 420920 159734 420972 159740
rect 420092 158908 420144 158914
rect 420092 158850 420144 158856
rect 419632 158772 419684 158778
rect 419632 158714 419684 158720
rect 419540 152516 419592 152522
rect 419540 152458 419592 152464
rect 419644 151978 419672 158714
rect 419724 154352 419776 154358
rect 419724 154294 419776 154300
rect 419632 151972 419684 151978
rect 419632 151914 419684 151920
rect 419736 150090 419764 154294
rect 421024 152998 421052 163254
rect 421668 163146 421696 163254
rect 421746 163200 421802 164400
rect 422312 163254 422524 163282
rect 421760 163146 421788 163200
rect 421668 163118 421788 163146
rect 422312 153134 422340 163254
rect 422496 163146 422524 163254
rect 422574 163200 422630 164400
rect 422772 163254 423352 163282
rect 422588 163146 422616 163200
rect 422496 163118 422616 163146
rect 422772 157334 422800 163254
rect 423324 163146 423352 163254
rect 423402 163200 423458 164400
rect 424322 163200 424378 164400
rect 425150 163200 425206 164400
rect 425978 163200 426034 164400
rect 426452 163254 426756 163282
rect 423416 163146 423444 163200
rect 423324 163118 423444 163146
rect 424336 159866 424364 163200
rect 424324 159860 424376 159866
rect 424324 159802 424376 159808
rect 424876 159520 424928 159526
rect 424876 159462 424928 159468
rect 423220 158908 423272 158914
rect 423220 158850 423272 158856
rect 422772 157306 423076 157334
rect 422392 154420 422444 154426
rect 422392 154362 422444 154368
rect 422208 153128 422260 153134
rect 422208 153070 422260 153076
rect 422300 153128 422352 153134
rect 422300 153070 422352 153076
rect 421012 152992 421064 152998
rect 421012 152934 421064 152940
rect 421656 152720 421708 152726
rect 421656 152662 421708 152668
rect 420368 152448 420420 152454
rect 420368 152390 420420 152396
rect 420380 150090 420408 152390
rect 421012 152040 421064 152046
rect 421012 151982 421064 151988
rect 421024 150090 421052 151982
rect 421668 150090 421696 152662
rect 421760 152658 421972 152674
rect 421748 152652 421984 152658
rect 421800 152646 421932 152652
rect 421748 152594 421800 152600
rect 421932 152594 421984 152600
rect 421930 152552 421986 152561
rect 421930 152487 421932 152496
rect 421984 152487 421986 152496
rect 421932 152458 421984 152464
rect 422220 152454 422248 153070
rect 422208 152448 422260 152454
rect 422208 152390 422260 152396
rect 422404 150090 422432 154362
rect 422944 153876 422996 153882
rect 422944 153818 422996 153824
rect 422852 152516 422904 152522
rect 422852 152458 422904 152464
rect 422864 152318 422892 152458
rect 422852 152312 422904 152318
rect 422852 152254 422904 152260
rect 418448 150062 418522 150090
rect 419092 150062 419166 150090
rect 419736 150062 419810 150090
rect 420380 150062 420454 150090
rect 421024 150062 421098 150090
rect 421668 150062 421742 150090
rect 418494 149940 418522 150062
rect 419138 149940 419166 150062
rect 419782 149940 419810 150062
rect 420426 149940 420454 150062
rect 421070 149940 421098 150062
rect 421714 149940 421742 150062
rect 422358 150062 422432 150090
rect 422956 150090 422984 153818
rect 423048 152454 423076 157306
rect 423128 153128 423180 153134
rect 423128 153070 423180 153076
rect 423036 152448 423088 152454
rect 423036 152390 423088 152396
rect 423140 152318 423168 153070
rect 423128 152312 423180 152318
rect 423128 152254 423180 152260
rect 423232 151978 423260 158850
rect 424506 152552 424562 152561
rect 424506 152487 424562 152496
rect 424520 152386 424548 152487
rect 424416 152380 424468 152386
rect 424416 152322 424468 152328
rect 424508 152380 424560 152386
rect 424508 152322 424560 152328
rect 424324 152244 424376 152250
rect 424324 152186 424376 152192
rect 423588 152108 423640 152114
rect 423588 152050 423640 152056
rect 423220 151972 423272 151978
rect 423220 151914 423272 151920
rect 423600 150090 423628 152050
rect 424336 151842 424364 152186
rect 424428 152114 424456 152322
rect 424416 152108 424468 152114
rect 424416 152050 424468 152056
rect 424232 151836 424284 151842
rect 424232 151778 424284 151784
rect 424324 151836 424376 151842
rect 424324 151778 424376 151784
rect 424244 150090 424272 151778
rect 424888 150226 424916 159462
rect 425164 153134 425192 163200
rect 425520 153944 425572 153950
rect 425520 153886 425572 153892
rect 425152 153128 425204 153134
rect 425152 153070 425204 153076
rect 424888 150198 424962 150226
rect 422956 150062 423030 150090
rect 423600 150062 423674 150090
rect 424244 150062 424318 150090
rect 422358 149940 422386 150062
rect 423002 149940 423030 150062
rect 423646 149940 423674 150062
rect 424290 149940 424318 150062
rect 424934 149940 424962 150198
rect 425532 150090 425560 153886
rect 425992 152250 426020 163200
rect 426452 152726 426480 163254
rect 426728 163146 426756 163254
rect 426806 163200 426862 164400
rect 427634 163200 427690 164400
rect 427832 163254 428412 163282
rect 426820 163146 426848 163200
rect 426728 163118 426848 163146
rect 427648 159458 427676 163200
rect 427360 159452 427412 159458
rect 427360 159394 427412 159400
rect 427636 159452 427688 159458
rect 427636 159394 427688 159400
rect 426348 152720 426400 152726
rect 426348 152662 426400 152668
rect 426440 152720 426492 152726
rect 426440 152662 426492 152668
rect 426072 152584 426124 152590
rect 426072 152526 426124 152532
rect 426360 152538 426388 152662
rect 426532 152584 426584 152590
rect 426360 152532 426532 152538
rect 426360 152526 426584 152532
rect 425980 152244 426032 152250
rect 425980 152186 426032 152192
rect 426084 150226 426112 152526
rect 426360 152510 426572 152526
rect 426900 152380 426952 152386
rect 426900 152322 426952 152328
rect 426912 151910 426940 152322
rect 426808 151904 426860 151910
rect 426808 151846 426860 151852
rect 426900 151904 426952 151910
rect 426900 151846 426952 151852
rect 426084 150198 426250 150226
rect 425532 150062 425606 150090
rect 425578 149940 425606 150062
rect 426222 149940 426250 150198
rect 426820 150090 426848 151846
rect 427372 150226 427400 159394
rect 427832 152386 427860 163254
rect 428384 163146 428412 163254
rect 428462 163200 428518 164400
rect 429290 163200 429346 164400
rect 429396 163254 430160 163282
rect 428476 163146 428504 163200
rect 428384 163118 428504 163146
rect 429304 152794 429332 163200
rect 428004 152788 428056 152794
rect 428004 152730 428056 152736
rect 429292 152788 429344 152794
rect 429292 152730 429344 152736
rect 427820 152380 427872 152386
rect 427820 152322 427872 152328
rect 428016 150226 428044 152730
rect 429396 152658 429424 163254
rect 430132 163146 430160 163254
rect 430210 163200 430266 164400
rect 430684 163254 430988 163282
rect 430224 163146 430252 163200
rect 430132 163118 430252 163146
rect 429936 159656 429988 159662
rect 429936 159598 429988 159604
rect 429200 152652 429252 152658
rect 429200 152594 429252 152600
rect 429384 152652 429436 152658
rect 429384 152594 429436 152600
rect 428648 152176 428700 152182
rect 428648 152118 428700 152124
rect 428660 150226 428688 152118
rect 429212 151814 429240 152594
rect 429212 151786 429332 151814
rect 429304 150226 429332 151786
rect 429948 150226 429976 159598
rect 430578 152416 430634 152425
rect 430578 152351 430634 152360
rect 430592 150226 430620 152351
rect 430684 152182 430712 163254
rect 430960 163146 430988 163254
rect 431038 163200 431094 164400
rect 431236 163254 431816 163282
rect 431052 163146 431080 163200
rect 430960 163118 431080 163146
rect 431132 153060 431184 153066
rect 431132 153002 431184 153008
rect 430672 152176 430724 152182
rect 430672 152118 430724 152124
rect 431144 151814 431172 153002
rect 431236 152561 431264 163254
rect 431788 163146 431816 163254
rect 431866 163200 431922 164400
rect 431972 163254 432644 163282
rect 431880 163146 431908 163200
rect 431788 163118 431908 163146
rect 431972 153066 432000 163254
rect 432616 163146 432644 163254
rect 432694 163200 432750 164400
rect 433522 163200 433578 164400
rect 433628 163254 433932 163282
rect 432708 163146 432736 163200
rect 432616 163118 432736 163146
rect 433536 163146 433564 163200
rect 433628 163146 433656 163254
rect 433536 163118 433656 163146
rect 432512 159588 432564 159594
rect 432512 159530 432564 159536
rect 431960 153060 432012 153066
rect 431960 153002 432012 153008
rect 431222 152552 431278 152561
rect 431222 152487 431278 152496
rect 431868 151836 431920 151842
rect 431144 151786 431264 151814
rect 431236 150226 431264 151786
rect 431868 151778 431920 151784
rect 431880 150226 431908 151778
rect 432524 150226 432552 159530
rect 433156 152856 433208 152862
rect 433156 152798 433208 152804
rect 433168 150226 433196 152798
rect 433904 152114 433932 163254
rect 434350 163200 434406 164400
rect 434732 163254 435128 163282
rect 434364 152862 434392 163200
rect 434732 153134 434760 163254
rect 435100 163146 435128 163254
rect 435178 163200 435234 164400
rect 436098 163200 436154 164400
rect 436926 163200 436982 164400
rect 437492 163254 437704 163282
rect 435192 163146 435220 163200
rect 435100 163118 435220 163146
rect 435088 159384 435140 159390
rect 435088 159326 435140 159332
rect 434628 153128 434680 153134
rect 434628 153070 434680 153076
rect 434720 153128 434772 153134
rect 434720 153070 434772 153076
rect 434352 152856 434404 152862
rect 434352 152798 434404 152804
rect 433800 152108 433852 152114
rect 433800 152050 433852 152056
rect 433892 152108 433944 152114
rect 433892 152050 433944 152056
rect 433812 150226 433840 152050
rect 434640 152046 434668 153070
rect 434444 152040 434496 152046
rect 434444 151982 434496 151988
rect 434628 152040 434680 152046
rect 434628 151982 434680 151988
rect 434456 150226 434484 151982
rect 435100 150226 435128 159326
rect 435732 152516 435784 152522
rect 435732 152458 435784 152464
rect 435744 150226 435772 152458
rect 436112 151842 436140 163200
rect 436376 152924 436428 152930
rect 436376 152866 436428 152872
rect 436100 151836 436152 151842
rect 436100 151778 436152 151784
rect 436388 150226 436416 152866
rect 436940 152522 436968 163200
rect 436928 152516 436980 152522
rect 436928 152458 436980 152464
rect 437492 151910 437520 163254
rect 437676 163146 437704 163254
rect 437754 163200 437810 164400
rect 437860 163254 438532 163282
rect 437768 163146 437796 163200
rect 437676 163118 437796 163146
rect 437664 159724 437716 159730
rect 437664 159666 437716 159672
rect 437572 153196 437624 153202
rect 437572 153138 437624 153144
rect 437584 152998 437612 153138
rect 437572 152992 437624 152998
rect 437572 152934 437624 152940
rect 437020 151904 437072 151910
rect 437020 151846 437072 151852
rect 437480 151904 437532 151910
rect 437480 151846 437532 151852
rect 437032 150226 437060 151846
rect 437676 150226 437704 159666
rect 437860 153202 437888 163254
rect 438504 163146 438532 163254
rect 438582 163200 438638 164400
rect 438872 163254 439360 163282
rect 438596 163146 438624 163200
rect 438504 163118 438624 163146
rect 437848 153196 437900 153202
rect 437848 153138 437900 153144
rect 438308 152992 438360 152998
rect 438308 152934 438360 152940
rect 438320 150226 438348 152934
rect 438872 152930 438900 163254
rect 439332 163146 439360 163254
rect 439410 163200 439466 164400
rect 440238 163200 440294 164400
rect 440344 163254 441016 163282
rect 439424 163146 439452 163200
rect 439332 163118 439452 163146
rect 439044 152992 439096 152998
rect 439044 152934 439096 152940
rect 438860 152924 438912 152930
rect 438860 152866 438912 152872
rect 439056 152590 439084 152934
rect 438952 152584 439004 152590
rect 438952 152526 439004 152532
rect 439044 152584 439096 152590
rect 439044 152526 439096 152532
rect 438964 150226 438992 152526
rect 440252 151978 440280 163200
rect 440344 152998 440372 163254
rect 440988 163146 441016 163254
rect 441066 163200 441122 164400
rect 441632 163254 441936 163282
rect 441080 163146 441108 163200
rect 440988 163118 441108 163146
rect 440424 159792 440476 159798
rect 440424 159734 440476 159740
rect 440332 152992 440384 152998
rect 440332 152934 440384 152940
rect 439596 151972 439648 151978
rect 439596 151914 439648 151920
rect 440240 151972 440292 151978
rect 440240 151914 440292 151920
rect 439608 150226 439636 151914
rect 440436 151814 440464 159734
rect 440884 152584 440936 152590
rect 440884 152526 440936 152532
rect 440344 151786 440464 151814
rect 440344 150226 440372 151786
rect 427372 150198 427446 150226
rect 428016 150198 428090 150226
rect 428660 150198 428734 150226
rect 429304 150198 429378 150226
rect 429948 150198 430022 150226
rect 430592 150198 430666 150226
rect 431236 150198 431310 150226
rect 431880 150198 431954 150226
rect 432524 150198 432598 150226
rect 433168 150198 433242 150226
rect 433812 150198 433886 150226
rect 434456 150198 434530 150226
rect 435100 150198 435174 150226
rect 435744 150198 435818 150226
rect 436388 150198 436462 150226
rect 437032 150198 437106 150226
rect 437676 150198 437750 150226
rect 438320 150198 438394 150226
rect 438964 150198 439038 150226
rect 439608 150198 439682 150226
rect 426820 150062 426894 150090
rect 426866 149940 426894 150062
rect 427418 149940 427446 150198
rect 428062 149940 428090 150198
rect 428706 149940 428734 150198
rect 429350 149940 429378 150198
rect 429994 149940 430022 150198
rect 430638 149940 430666 150198
rect 431282 149940 431310 150198
rect 431926 149940 431954 150198
rect 432570 149940 432598 150198
rect 433214 149940 433242 150198
rect 433858 149940 433886 150198
rect 434502 149940 434530 150198
rect 435146 149940 435174 150198
rect 435790 149940 435818 150198
rect 436434 149940 436462 150198
rect 437078 149940 437106 150198
rect 437722 149940 437750 150198
rect 438366 149940 438394 150198
rect 439010 149940 439038 150198
rect 439654 149940 439682 150198
rect 440298 150198 440372 150226
rect 440896 150226 440924 152526
rect 441632 152318 441660 163254
rect 441908 163146 441936 163254
rect 441986 163200 442042 164400
rect 442092 163254 442764 163282
rect 442000 163146 442028 163200
rect 441908 163118 442028 163146
rect 442092 153066 442120 163254
rect 442736 163146 442764 163254
rect 442814 163200 442870 164400
rect 443012 163254 443592 163282
rect 442828 163146 442856 163200
rect 442736 163118 442856 163146
rect 442816 159860 442868 159866
rect 442816 159802 442868 159808
rect 441988 153060 442040 153066
rect 441988 153002 442040 153008
rect 442080 153060 442132 153066
rect 442080 153002 442132 153008
rect 442000 152658 442028 153002
rect 441988 152652 442040 152658
rect 441988 152594 442040 152600
rect 442172 152448 442224 152454
rect 442172 152390 442224 152396
rect 441528 152312 441580 152318
rect 441528 152254 441580 152260
rect 441620 152312 441672 152318
rect 441620 152254 441672 152260
rect 441540 150226 441568 152254
rect 442184 150226 442212 152390
rect 442828 150226 442856 159802
rect 443012 152454 443040 163254
rect 443564 163146 443592 163254
rect 443642 163200 443698 164400
rect 444470 163200 444526 164400
rect 445298 163200 445354 164400
rect 446126 163200 446182 164400
rect 446324 163254 446904 163282
rect 443656 163146 443684 163200
rect 443564 163118 443684 163146
rect 443920 153128 443972 153134
rect 443918 153096 443920 153105
rect 444012 153128 444064 153134
rect 443972 153096 443974 153105
rect 444012 153070 444064 153076
rect 443918 153031 443974 153040
rect 444024 152862 444052 153070
rect 444012 152856 444064 152862
rect 444012 152798 444064 152804
rect 444484 152794 444512 163200
rect 444930 153096 444986 153105
rect 444930 153031 444986 153040
rect 444944 152794 444972 153031
rect 444472 152788 444524 152794
rect 444472 152730 444524 152736
rect 444932 152788 444984 152794
rect 444932 152730 444984 152736
rect 444748 152720 444800 152726
rect 444748 152662 444800 152668
rect 443000 152448 443052 152454
rect 443000 152390 443052 152396
rect 444104 152244 444156 152250
rect 444104 152186 444156 152192
rect 443460 152040 443512 152046
rect 443460 151982 443512 151988
rect 443472 150226 443500 151982
rect 444116 150226 444144 152186
rect 444760 150226 444788 152662
rect 445312 152250 445340 163200
rect 446140 159866 446168 163200
rect 446128 159860 446180 159866
rect 446128 159802 446180 159808
rect 445392 159452 445444 159458
rect 445392 159394 445444 159400
rect 445300 152244 445352 152250
rect 445300 152186 445352 152192
rect 445404 150226 445432 159394
rect 446128 152652 446180 152658
rect 446128 152594 446180 152600
rect 446140 152386 446168 152594
rect 446036 152380 446088 152386
rect 446036 152322 446088 152328
rect 446128 152380 446180 152386
rect 446128 152322 446180 152328
rect 446048 150226 446076 152322
rect 446324 152046 446352 163254
rect 446876 163146 446904 163254
rect 446954 163200 447010 164400
rect 447874 163200 447930 164400
rect 448702 163200 448758 164400
rect 449530 163200 449586 164400
rect 450358 163200 450414 164400
rect 451186 163200 451242 164400
rect 452014 163200 452070 164400
rect 452842 163200 452898 164400
rect 453762 163200 453818 164400
rect 454590 163200 454646 164400
rect 455418 163200 455474 164400
rect 456246 163200 456302 164400
rect 457074 163200 457130 164400
rect 457902 163200 457958 164400
rect 458730 163200 458786 164400
rect 459650 163200 459706 164400
rect 460478 163200 460534 164400
rect 461306 163200 461362 164400
rect 462134 163200 462190 164400
rect 462962 163200 463018 164400
rect 463790 163200 463846 164400
rect 464618 163200 464674 164400
rect 465538 163200 465594 164400
rect 466366 163200 466422 164400
rect 467194 163200 467250 164400
rect 468022 163200 468078 164400
rect 468850 163200 468906 164400
rect 469678 163200 469734 164400
rect 470506 163200 470562 164400
rect 471426 163200 471482 164400
rect 472254 163200 472310 164400
rect 473082 163200 473138 164400
rect 473910 163200 473966 164400
rect 474738 163200 474794 164400
rect 475566 163200 475622 164400
rect 476394 163200 476450 164400
rect 477314 163200 477370 164400
rect 478142 163200 478198 164400
rect 478970 163200 479026 164400
rect 479798 163200 479854 164400
rect 480626 163200 480682 164400
rect 481454 163200 481510 164400
rect 482282 163200 482338 164400
rect 483202 163200 483258 164400
rect 484030 163200 484086 164400
rect 484504 163254 484808 163282
rect 446968 163146 446996 163200
rect 446876 163118 446996 163146
rect 447888 159050 447916 163200
rect 448716 159390 448744 163200
rect 449544 159730 449572 163200
rect 450372 159798 450400 163200
rect 450360 159792 450412 159798
rect 450360 159734 450412 159740
rect 449532 159724 449584 159730
rect 449532 159666 449584 159672
rect 451200 159458 451228 163200
rect 452028 159594 452056 163200
rect 452016 159588 452068 159594
rect 452016 159530 452068 159536
rect 451188 159452 451240 159458
rect 451188 159394 451240 159400
rect 448704 159384 448756 159390
rect 448704 159326 448756 159332
rect 447876 159044 447928 159050
rect 447876 158986 447928 158992
rect 452856 158778 452884 163200
rect 453776 159662 453804 163200
rect 453764 159656 453816 159662
rect 453764 159598 453816 159604
rect 454604 158914 454632 163200
rect 454592 158908 454644 158914
rect 454592 158850 454644 158856
rect 455432 158846 455460 163200
rect 456260 158982 456288 163200
rect 456800 159860 456852 159866
rect 456800 159802 456852 159808
rect 456248 158976 456300 158982
rect 456248 158918 456300 158924
rect 455420 158840 455472 158846
rect 455420 158782 455472 158788
rect 452844 158772 452896 158778
rect 452844 158714 452896 158720
rect 456812 153202 456840 159802
rect 457088 159254 457116 163200
rect 457916 159322 457944 163200
rect 458744 159866 458772 163200
rect 458732 159860 458784 159866
rect 458732 159802 458784 159808
rect 459664 159526 459692 163200
rect 459652 159520 459704 159526
rect 459652 159462 459704 159468
rect 457904 159316 457956 159322
rect 457904 159258 457956 159264
rect 457076 159248 457128 159254
rect 457076 159190 457128 159196
rect 460492 159118 460520 163200
rect 460940 159724 460992 159730
rect 460940 159666 460992 159672
rect 460480 159112 460532 159118
rect 460480 159054 460532 159060
rect 460112 159044 460164 159050
rect 460112 158986 460164 158992
rect 459560 158772 459612 158778
rect 459560 158714 459612 158720
rect 446404 153196 446456 153202
rect 446404 153138 446456 153144
rect 456800 153196 456852 153202
rect 456800 153138 456852 153144
rect 459468 153196 459520 153202
rect 459468 153138 459520 153144
rect 446416 152658 446444 153138
rect 450544 153128 450596 153134
rect 450544 153070 450596 153076
rect 447416 153060 447468 153066
rect 447416 153002 447468 153008
rect 446680 152856 446732 152862
rect 446680 152798 446732 152804
rect 446772 152856 446824 152862
rect 446772 152798 446824 152804
rect 446404 152652 446456 152658
rect 446404 152594 446456 152600
rect 446312 152040 446364 152046
rect 446312 151982 446364 151988
rect 446692 150226 446720 152798
rect 446784 152522 446812 152798
rect 447428 152590 447456 153002
rect 447324 152584 447376 152590
rect 447324 152526 447376 152532
rect 447416 152584 447468 152590
rect 447416 152526 447468 152532
rect 448610 152552 448666 152561
rect 446772 152516 446824 152522
rect 446772 152458 446824 152464
rect 447336 150226 447364 152526
rect 448610 152487 448666 152496
rect 447968 152176 448020 152182
rect 447968 152118 448020 152124
rect 447980 150226 448008 152118
rect 448624 150226 448652 152487
rect 449256 152380 449308 152386
rect 449256 152322 449308 152328
rect 449268 150226 449296 152322
rect 449900 152108 449952 152114
rect 449900 152050 449952 152056
rect 449912 150226 449940 152050
rect 450556 150226 450584 153070
rect 455696 152992 455748 152998
rect 455696 152934 455748 152940
rect 454408 152924 454460 152930
rect 454408 152866 454460 152872
rect 452476 152856 452528 152862
rect 452476 152798 452528 152804
rect 451188 152788 451240 152794
rect 451188 152730 451240 152736
rect 451200 150226 451228 152730
rect 451832 151836 451884 151842
rect 451832 151778 451884 151784
rect 451844 150226 451872 151778
rect 452488 150226 452516 152798
rect 453764 152652 453816 152658
rect 453764 152594 453816 152600
rect 453120 151904 453172 151910
rect 453120 151846 453172 151852
rect 453132 150226 453160 151846
rect 453776 150226 453804 152594
rect 454420 150226 454448 152866
rect 455052 151972 455104 151978
rect 455052 151914 455104 151920
rect 455064 150226 455092 151914
rect 455708 150226 455736 152934
rect 458180 152720 458232 152726
rect 458180 152662 458232 152668
rect 456984 152584 457036 152590
rect 456984 152526 457036 152532
rect 456340 152312 456392 152318
rect 456340 152254 456392 152260
rect 456352 150226 456380 152254
rect 456996 150226 457024 152526
rect 457628 152448 457680 152454
rect 457628 152390 457680 152396
rect 457640 150226 457668 152390
rect 458192 150226 458220 152662
rect 458824 152244 458876 152250
rect 458824 152186 458876 152192
rect 458836 150226 458864 152186
rect 459480 150226 459508 153138
rect 459572 152522 459600 158714
rect 459560 152516 459612 152522
rect 459560 152458 459612 152464
rect 460020 152040 460072 152046
rect 460020 151982 460072 151988
rect 440896 150198 440970 150226
rect 441540 150198 441614 150226
rect 442184 150198 442258 150226
rect 442828 150198 442902 150226
rect 443472 150198 443546 150226
rect 444116 150198 444190 150226
rect 444760 150198 444834 150226
rect 445404 150198 445478 150226
rect 446048 150198 446122 150226
rect 446692 150198 446766 150226
rect 447336 150198 447410 150226
rect 447980 150198 448054 150226
rect 448624 150198 448698 150226
rect 449268 150198 449342 150226
rect 449912 150198 449986 150226
rect 450556 150198 450630 150226
rect 451200 150198 451274 150226
rect 451844 150198 451918 150226
rect 452488 150198 452562 150226
rect 453132 150198 453206 150226
rect 453776 150198 453850 150226
rect 454420 150198 454494 150226
rect 455064 150198 455138 150226
rect 455708 150198 455782 150226
rect 456352 150198 456426 150226
rect 456996 150198 457070 150226
rect 457640 150198 457714 150226
rect 458192 150198 458266 150226
rect 458836 150198 458910 150226
rect 459480 150198 459554 150226
rect 440298 149940 440326 150198
rect 440942 149940 440970 150198
rect 441586 149940 441614 150198
rect 442230 149940 442258 150198
rect 442874 149940 442902 150198
rect 443518 149940 443546 150198
rect 444162 149940 444190 150198
rect 444806 149940 444834 150198
rect 445450 149940 445478 150198
rect 446094 149940 446122 150198
rect 446738 149940 446766 150198
rect 447382 149940 447410 150198
rect 448026 149940 448054 150198
rect 448670 149940 448698 150198
rect 449314 149940 449342 150198
rect 449958 149940 449986 150198
rect 450602 149940 450630 150198
rect 451246 149940 451274 150198
rect 451890 149940 451918 150198
rect 452534 149940 452562 150198
rect 453178 149940 453206 150198
rect 453822 149940 453850 150198
rect 454466 149940 454494 150198
rect 455110 149940 455138 150198
rect 455754 149940 455782 150198
rect 456398 149940 456426 150198
rect 457042 149940 457070 150198
rect 457686 149940 457714 150198
rect 458238 149940 458266 150198
rect 458882 149940 458910 150198
rect 459526 149940 459554 150198
rect 460032 150192 460060 151982
rect 460124 151814 460152 158986
rect 460124 151786 460796 151814
rect 460768 150226 460796 151786
rect 460768 150198 460842 150226
rect 460952 150210 460980 159666
rect 461320 159186 461348 163200
rect 461400 159384 461452 159390
rect 461400 159326 461452 159332
rect 461308 159180 461360 159186
rect 461308 159122 461360 159128
rect 461412 150226 461440 159326
rect 462148 159050 462176 163200
rect 462320 159792 462372 159798
rect 462320 159734 462372 159740
rect 462136 159044 462188 159050
rect 462136 158986 462188 158992
rect 461860 158908 461912 158914
rect 461860 158850 461912 158856
rect 461872 153202 461900 158850
rect 461860 153196 461912 153202
rect 461860 153138 461912 153144
rect 462332 151814 462360 159734
rect 462872 159452 462924 159458
rect 462872 159394 462924 159400
rect 462780 158840 462832 158846
rect 462780 158782 462832 158788
rect 462792 153134 462820 158782
rect 462780 153128 462832 153134
rect 462780 153070 462832 153076
rect 462884 151814 462912 159394
rect 462976 158778 463004 163200
rect 463804 159730 463832 163200
rect 463792 159724 463844 159730
rect 463792 159666 463844 159672
rect 463976 159588 464028 159594
rect 463976 159530 464028 159536
rect 463148 158976 463200 158982
rect 463148 158918 463200 158924
rect 462964 158772 463016 158778
rect 462964 158714 463016 158720
rect 463160 153066 463188 158918
rect 463148 153060 463200 153066
rect 463148 153002 463200 153008
rect 462332 151786 462728 151814
rect 462884 151786 463372 151814
rect 462700 150226 462728 151786
rect 463344 150226 463372 151786
rect 463988 150226 464016 159530
rect 464436 159316 464488 159322
rect 464436 159258 464488 159264
rect 464160 159248 464212 159254
rect 464160 159190 464212 159196
rect 464172 152998 464200 159190
rect 464160 152992 464212 152998
rect 464160 152934 464212 152940
rect 464448 152930 464476 159258
rect 464632 158846 464660 163200
rect 465080 159860 465132 159866
rect 465080 159802 465132 159808
rect 464620 158840 464672 158846
rect 464620 158782 464672 158788
rect 464436 152924 464488 152930
rect 464436 152866 464488 152872
rect 465092 152862 465120 159802
rect 465264 159656 465316 159662
rect 465264 159598 465316 159604
rect 465080 152856 465132 152862
rect 465080 152798 465132 152804
rect 464620 152516 464672 152522
rect 464620 152458 464672 152464
rect 464632 150226 464660 152458
rect 465276 150226 465304 159598
rect 465552 158914 465580 163200
rect 466380 158982 466408 163200
rect 467208 159594 467236 163200
rect 468036 159662 468064 163200
rect 468024 159656 468076 159662
rect 468024 159598 468076 159604
rect 467196 159588 467248 159594
rect 467196 159530 467248 159536
rect 468864 159526 468892 163200
rect 466644 159520 466696 159526
rect 466644 159462 466696 159468
rect 468852 159520 468904 159526
rect 468852 159462 468904 159468
rect 466460 159112 466512 159118
rect 466460 159054 466512 159060
rect 466368 158976 466420 158982
rect 466368 158918 466420 158924
rect 465540 158908 465592 158914
rect 465540 158850 465592 158856
rect 466472 153202 466500 159054
rect 465908 153196 465960 153202
rect 465908 153138 465960 153144
rect 466460 153196 466512 153202
rect 466460 153138 466512 153144
rect 465920 150226 465948 153138
rect 466656 153134 466684 159462
rect 469692 159390 469720 163200
rect 470520 159866 470548 163200
rect 471440 159866 471468 163200
rect 470508 159860 470560 159866
rect 470508 159802 470560 159808
rect 471428 159860 471480 159866
rect 471428 159802 471480 159808
rect 471428 159724 471480 159730
rect 471428 159666 471480 159672
rect 469680 159384 469732 159390
rect 469680 159326 469732 159332
rect 468024 159180 468076 159186
rect 468024 159122 468076 159128
rect 467932 159044 467984 159050
rect 467932 158986 467984 158992
rect 466552 153128 466604 153134
rect 466552 153070 466604 153076
rect 466644 153128 466696 153134
rect 466644 153070 466696 153076
rect 466564 150226 466592 153070
rect 467196 153060 467248 153066
rect 467196 153002 467248 153008
rect 467208 150226 467236 153002
rect 467840 152992 467892 152998
rect 467840 152934 467892 152940
rect 467852 150226 467880 152934
rect 467944 151842 467972 158986
rect 468036 151910 468064 159122
rect 469220 158772 469272 158778
rect 469220 158714 469272 158720
rect 468392 152924 468444 152930
rect 468392 152866 468444 152872
rect 468024 151904 468076 151910
rect 468024 151846 468076 151852
rect 467932 151836 467984 151842
rect 468404 151814 468432 152866
rect 469128 152856 469180 152862
rect 469128 152798 469180 152804
rect 468404 151786 468524 151814
rect 467932 151778 467984 151784
rect 468496 150226 468524 151786
rect 469140 150226 469168 152798
rect 469232 151978 469260 158714
rect 470416 153196 470468 153202
rect 470416 153138 470468 153144
rect 469772 153128 469824 153134
rect 469772 153070 469824 153076
rect 469220 151972 469272 151978
rect 469220 151914 469272 151920
rect 469784 150226 469812 153070
rect 470428 150226 470456 153138
rect 471440 152998 471468 159666
rect 472268 159118 472296 163200
rect 473096 159798 473124 163200
rect 473084 159792 473136 159798
rect 473084 159734 473136 159740
rect 473360 159588 473412 159594
rect 473360 159530 473412 159536
rect 472256 159112 472308 159118
rect 472256 159054 472308 159060
rect 472624 158976 472676 158982
rect 472624 158918 472676 158924
rect 472256 158908 472308 158914
rect 472256 158850 472308 158856
rect 471520 158840 471572 158846
rect 471520 158782 471572 158788
rect 471532 153202 471560 158782
rect 471520 153196 471572 153202
rect 471520 153138 471572 153144
rect 472268 153134 472296 158850
rect 472256 153128 472308 153134
rect 472256 153070 472308 153076
rect 472636 153066 472664 158918
rect 472624 153060 472676 153066
rect 472624 153002 472676 153008
rect 473372 152998 473400 159530
rect 473924 159050 473952 163200
rect 473912 159044 473964 159050
rect 473912 158986 473964 158992
rect 474752 158914 474780 163200
rect 474832 159520 474884 159526
rect 474832 159462 474884 159468
rect 474740 158908 474792 158914
rect 474740 158850 474792 158856
rect 474844 153202 474872 159462
rect 475580 158982 475608 163200
rect 476120 159928 476172 159934
rect 476120 159870 476172 159876
rect 476028 159656 476080 159662
rect 476028 159598 476080 159604
rect 475568 158976 475620 158982
rect 475568 158918 475620 158924
rect 473636 153196 473688 153202
rect 473636 153138 473688 153144
rect 474832 153196 474884 153202
rect 474832 153138 474884 153144
rect 471428 152992 471480 152998
rect 471428 152934 471480 152940
rect 472992 152992 473044 152998
rect 472992 152934 473044 152940
rect 473360 152992 473412 152998
rect 473360 152934 473412 152940
rect 472348 151972 472400 151978
rect 472348 151914 472400 151920
rect 471060 151904 471112 151910
rect 471060 151846 471112 151852
rect 471072 150226 471100 151846
rect 471704 151836 471756 151842
rect 471704 151778 471756 151784
rect 471716 150226 471744 151778
rect 472360 150226 472388 151914
rect 473004 150226 473032 152934
rect 473648 150226 473676 153138
rect 474280 153128 474332 153134
rect 474280 153070 474332 153076
rect 474292 150226 474320 153070
rect 474924 153060 474976 153066
rect 474924 153002 474976 153008
rect 474936 150226 474964 153002
rect 475568 152992 475620 152998
rect 475568 152934 475620 152940
rect 475580 150226 475608 152934
rect 476040 151814 476068 159598
rect 476132 153134 476160 159870
rect 476408 158846 476436 163200
rect 477328 159526 477356 163200
rect 477684 159860 477736 159866
rect 477684 159802 477736 159808
rect 477316 159520 477368 159526
rect 477316 159462 477368 159468
rect 477408 159384 477460 159390
rect 477408 159326 477460 159332
rect 476396 158840 476448 158846
rect 476396 158782 476448 158788
rect 476948 153196 477000 153202
rect 476948 153138 477000 153144
rect 476120 153128 476172 153134
rect 476120 153070 476172 153076
rect 476040 151786 476252 151814
rect 476224 150226 476252 151786
rect 476960 150226 476988 153138
rect 477420 151814 477448 159326
rect 477420 151786 477540 151814
rect 460032 150164 460198 150192
rect 460170 149940 460198 150164
rect 460814 149940 460842 150198
rect 460940 150204 460992 150210
rect 461412 150198 461486 150226
rect 460940 150146 460992 150152
rect 461458 149940 461486 150198
rect 462090 150204 462142 150210
rect 462700 150198 462774 150226
rect 463344 150198 463418 150226
rect 463988 150198 464062 150226
rect 464632 150198 464706 150226
rect 465276 150198 465350 150226
rect 465920 150198 465994 150226
rect 466564 150198 466638 150226
rect 467208 150198 467282 150226
rect 467852 150198 467926 150226
rect 468496 150198 468570 150226
rect 469140 150198 469214 150226
rect 469784 150198 469858 150226
rect 470428 150198 470502 150226
rect 471072 150198 471146 150226
rect 471716 150198 471790 150226
rect 472360 150198 472434 150226
rect 473004 150198 473078 150226
rect 473648 150198 473722 150226
rect 474292 150198 474366 150226
rect 474936 150198 475010 150226
rect 475580 150198 475654 150226
rect 476224 150198 476298 150226
rect 462090 150146 462142 150152
rect 462102 149940 462130 150146
rect 462746 149940 462774 150198
rect 463390 149940 463418 150198
rect 464034 149940 464062 150198
rect 464678 149940 464706 150198
rect 465322 149940 465350 150198
rect 465966 149940 465994 150198
rect 466610 149940 466638 150198
rect 467254 149940 467282 150198
rect 467898 149940 467926 150198
rect 468542 149940 468570 150198
rect 469186 149940 469214 150198
rect 469830 149940 469858 150198
rect 470474 149940 470502 150198
rect 471118 149940 471146 150198
rect 471762 149940 471790 150198
rect 472406 149940 472434 150198
rect 473050 149940 473078 150198
rect 473694 149940 473722 150198
rect 474338 149940 474366 150198
rect 474982 149940 475010 150198
rect 475626 149940 475654 150198
rect 476270 149940 476298 150198
rect 476914 150198 476988 150226
rect 477512 150226 477540 151786
rect 477512 150198 477586 150226
rect 477696 150210 477724 159802
rect 478156 159390 478184 163200
rect 478984 159730 479012 163200
rect 478972 159724 479024 159730
rect 478972 159666 479024 159672
rect 479812 159662 479840 163200
rect 480640 159934 480668 163200
rect 480628 159928 480680 159934
rect 480628 159870 480680 159876
rect 480076 159792 480128 159798
rect 480076 159734 480128 159740
rect 479800 159656 479852 159662
rect 479800 159598 479852 159604
rect 478144 159384 478196 159390
rect 478144 159326 478196 159332
rect 479156 159112 479208 159118
rect 479156 159054 479208 159060
rect 478144 153128 478196 153134
rect 478144 153070 478196 153076
rect 478156 150226 478184 153070
rect 479168 151814 479196 159054
rect 479168 151786 479472 151814
rect 479444 150226 479472 151786
rect 480088 150226 480116 159734
rect 480260 159044 480312 159050
rect 480260 158986 480312 158992
rect 480272 151814 480300 158986
rect 481364 158908 481416 158914
rect 481364 158850 481416 158856
rect 480272 151786 480760 151814
rect 480732 150226 480760 151786
rect 481376 150226 481404 158850
rect 481468 158778 481496 163200
rect 481640 158976 481692 158982
rect 481640 158918 481692 158924
rect 481456 158772 481508 158778
rect 481456 158714 481508 158720
rect 481652 151814 481680 158918
rect 482296 158914 482324 163200
rect 483216 161474 483244 163200
rect 483124 161446 483244 161474
rect 482284 158908 482336 158914
rect 482284 158850 482336 158856
rect 482652 158840 482704 158846
rect 482652 158782 482704 158788
rect 481652 151786 482048 151814
rect 482020 150226 482048 151786
rect 482664 150226 482692 158782
rect 483124 152998 483152 161446
rect 483296 159520 483348 159526
rect 483296 159462 483348 159468
rect 483204 159384 483256 159390
rect 483204 159326 483256 159332
rect 483112 152992 483164 152998
rect 483112 152934 483164 152940
rect 476914 149940 476942 150198
rect 477558 149940 477586 150198
rect 477684 150204 477736 150210
rect 478156 150198 478230 150226
rect 477684 150146 477736 150152
rect 478202 149940 478230 150198
rect 478834 150204 478886 150210
rect 479444 150198 479518 150226
rect 480088 150198 480162 150226
rect 480732 150198 480806 150226
rect 481376 150198 481450 150226
rect 482020 150198 482094 150226
rect 482664 150198 482738 150226
rect 483216 150210 483244 159326
rect 483308 150226 483336 159462
rect 484044 153134 484072 163200
rect 484032 153128 484084 153134
rect 484032 153070 484084 153076
rect 484504 153066 484532 163254
rect 484780 163146 484808 163254
rect 484858 163200 484914 164400
rect 485686 163200 485742 164400
rect 485792 163254 486464 163282
rect 484872 163146 484900 163200
rect 484780 163118 484900 163146
rect 484676 159724 484728 159730
rect 484676 159666 484728 159672
rect 484492 153060 484544 153066
rect 484492 153002 484544 153008
rect 484688 150226 484716 159666
rect 485228 159656 485280 159662
rect 485228 159598 485280 159604
rect 478834 150146 478886 150152
rect 478846 149940 478874 150146
rect 479490 149940 479518 150198
rect 480134 149940 480162 150198
rect 480778 149940 480806 150198
rect 481422 149940 481450 150198
rect 482066 149940 482094 150198
rect 482710 149940 482738 150198
rect 483204 150204 483256 150210
rect 483308 150198 483382 150226
rect 483204 150146 483256 150152
rect 483354 149940 483382 150198
rect 483986 150204 484038 150210
rect 483986 150146 484038 150152
rect 484642 150198 484716 150226
rect 485240 150226 485268 159598
rect 485700 153202 485728 163200
rect 485688 153196 485740 153202
rect 485688 153138 485740 153144
rect 485792 152046 485820 163254
rect 486436 163146 486464 163254
rect 486514 163200 486570 164400
rect 487342 163200 487398 164400
rect 488170 163200 488226 164400
rect 488552 163254 489040 163282
rect 486528 163146 486556 163200
rect 486436 163118 486556 163146
rect 485964 159928 486016 159934
rect 485964 159870 486016 159876
rect 485780 152040 485832 152046
rect 485780 151982 485832 151988
rect 485976 150226 486004 159870
rect 487252 158908 487304 158914
rect 487252 158850 487304 158856
rect 486516 158772 486568 158778
rect 486516 158714 486568 158720
rect 485240 150198 485314 150226
rect 483998 149940 484026 150146
rect 484642 149940 484670 150198
rect 485286 149940 485314 150198
rect 485930 150198 486004 150226
rect 486528 150226 486556 158714
rect 487264 150226 487292 158850
rect 487356 151910 487384 163200
rect 487804 152992 487856 152998
rect 487804 152934 487856 152940
rect 487344 151904 487396 151910
rect 487344 151846 487396 151852
rect 486528 150198 486602 150226
rect 485930 149940 485958 150198
rect 486574 149940 486602 150198
rect 487218 150198 487292 150226
rect 487816 150226 487844 152934
rect 488184 151842 488212 163200
rect 488448 153128 488500 153134
rect 488448 153070 488500 153076
rect 488172 151836 488224 151842
rect 488172 151778 488224 151784
rect 488460 150226 488488 153070
rect 488552 151978 488580 163254
rect 489012 163146 489040 163254
rect 489090 163200 489146 164400
rect 489918 163200 489974 164400
rect 490746 163200 490802 164400
rect 491574 163200 491630 164400
rect 492402 163200 492458 164400
rect 492692 163254 493180 163282
rect 489104 163146 489132 163200
rect 489012 163118 489132 163146
rect 489644 153196 489696 153202
rect 489644 153138 489696 153144
rect 489000 153060 489052 153066
rect 489000 153002 489052 153008
rect 488540 151972 488592 151978
rect 488540 151914 488592 151920
rect 489012 150226 489040 153002
rect 489656 150226 489684 153138
rect 489932 152930 489960 163200
rect 490760 153202 490788 163200
rect 490748 153196 490800 153202
rect 490748 153138 490800 153144
rect 491588 152998 491616 163200
rect 492416 153134 492444 163200
rect 492404 153128 492456 153134
rect 492404 153070 492456 153076
rect 492692 153066 492720 163254
rect 493152 163146 493180 163254
rect 493230 163200 493286 164400
rect 494058 163200 494114 164400
rect 494978 163200 495034 164400
rect 495544 163254 495756 163282
rect 493244 163146 493272 163200
rect 493152 163118 493272 163146
rect 494072 153202 494100 163200
rect 493508 153196 493560 153202
rect 493508 153138 493560 153144
rect 494060 153196 494112 153202
rect 494060 153138 494112 153144
rect 492680 153060 492732 153066
rect 492680 153002 492732 153008
rect 491576 152992 491628 152998
rect 491576 152934 491628 152940
rect 489920 152924 489972 152930
rect 489920 152866 489972 152872
rect 492864 152924 492916 152930
rect 492864 152866 492916 152872
rect 490288 152040 490340 152046
rect 490288 151982 490340 151988
rect 490300 150226 490328 151982
rect 492220 151972 492272 151978
rect 492220 151914 492272 151920
rect 490932 151904 490984 151910
rect 490932 151846 490984 151852
rect 490944 150226 490972 151846
rect 491576 151836 491628 151842
rect 491576 151778 491628 151784
rect 491588 150226 491616 151778
rect 492232 150226 492260 151914
rect 492876 150226 492904 152866
rect 493520 150226 493548 153138
rect 494992 153134 495020 163200
rect 494796 153128 494848 153134
rect 494796 153070 494848 153076
rect 494980 153128 495032 153134
rect 494980 153070 495032 153076
rect 494152 152992 494204 152998
rect 494152 152934 494204 152940
rect 494164 150226 494192 152934
rect 494808 150226 494836 153070
rect 495544 153066 495572 163254
rect 495728 163146 495756 163254
rect 495806 163200 495862 164400
rect 496634 163200 496690 164400
rect 496832 163254 497412 163282
rect 495820 163146 495848 163200
rect 495728 163118 495848 163146
rect 496648 153202 496676 163200
rect 496084 153196 496136 153202
rect 496084 153138 496136 153144
rect 496636 153196 496688 153202
rect 496636 153138 496688 153144
rect 495440 153060 495492 153066
rect 495440 153002 495492 153008
rect 495532 153060 495584 153066
rect 495532 153002 495584 153008
rect 495452 150226 495480 153002
rect 496096 150226 496124 153138
rect 496832 153134 496860 163254
rect 497384 163146 497412 163254
rect 497462 163200 497518 164400
rect 498290 163200 498346 164400
rect 499118 163200 499174 164400
rect 499946 163200 500002 164400
rect 500052 163254 500632 163282
rect 497476 163146 497504 163200
rect 497384 163118 497504 163146
rect 498304 156670 498332 163200
rect 498292 156664 498344 156670
rect 498292 156606 498344 156612
rect 498016 153196 498068 153202
rect 498016 153138 498068 153144
rect 496728 153128 496780 153134
rect 496728 153070 496780 153076
rect 496820 153128 496872 153134
rect 496820 153070 496872 153076
rect 496740 150226 496768 153070
rect 497372 153060 497424 153066
rect 497372 153002 497424 153008
rect 497384 150226 497412 153002
rect 498028 150226 498056 153138
rect 498660 153128 498712 153134
rect 498660 153070 498712 153076
rect 498672 150226 498700 153070
rect 499132 151842 499160 163200
rect 499960 163146 499988 163200
rect 500052 163146 500080 163254
rect 499960 163118 500080 163146
rect 499304 156664 499356 156670
rect 499304 156606 499356 156612
rect 499120 151836 499172 151842
rect 499120 151778 499172 151784
rect 499316 150226 499344 156606
rect 499948 151836 500000 151842
rect 499948 151778 500000 151784
rect 499960 150226 499988 151778
rect 500604 150226 500632 163254
rect 500866 163200 500922 164400
rect 501694 163200 501750 164400
rect 502522 163200 502578 164400
rect 503350 163200 503406 164400
rect 503824 163254 504128 163282
rect 500880 151814 500908 163200
rect 501708 161474 501736 163200
rect 501708 161446 501920 161474
rect 500880 151786 501276 151814
rect 501248 150226 501276 151786
rect 501892 150226 501920 161446
rect 502340 156664 502392 156670
rect 502340 156606 502392 156612
rect 487816 150198 487890 150226
rect 488460 150198 488534 150226
rect 489012 150198 489086 150226
rect 489656 150198 489730 150226
rect 490300 150198 490374 150226
rect 490944 150198 491018 150226
rect 491588 150198 491662 150226
rect 492232 150198 492306 150226
rect 492876 150198 492950 150226
rect 493520 150198 493594 150226
rect 494164 150198 494238 150226
rect 494808 150198 494882 150226
rect 495452 150198 495526 150226
rect 496096 150198 496170 150226
rect 496740 150198 496814 150226
rect 497384 150198 497458 150226
rect 498028 150198 498102 150226
rect 498672 150198 498746 150226
rect 499316 150198 499390 150226
rect 499960 150198 500034 150226
rect 500604 150198 500678 150226
rect 501248 150198 501322 150226
rect 501892 150198 501966 150226
rect 502352 150210 502380 156606
rect 502536 150226 502564 163200
rect 503364 156670 503392 163200
rect 503352 156664 503404 156670
rect 503352 156606 503404 156612
rect 503720 156664 503772 156670
rect 503720 156606 503772 156612
rect 487218 149940 487246 150198
rect 487862 149940 487890 150198
rect 488506 149940 488534 150198
rect 489058 149940 489086 150198
rect 489702 149940 489730 150198
rect 490346 149940 490374 150198
rect 490990 149940 491018 150198
rect 491634 149940 491662 150198
rect 492278 149940 492306 150198
rect 492922 149940 492950 150198
rect 493566 149940 493594 150198
rect 494210 149940 494238 150198
rect 494854 149940 494882 150198
rect 495498 149940 495526 150198
rect 496142 149940 496170 150198
rect 496786 149940 496814 150198
rect 497430 149940 497458 150198
rect 498074 149940 498102 150198
rect 498718 149940 498746 150198
rect 499362 149940 499390 150198
rect 500006 149940 500034 150198
rect 500650 149940 500678 150198
rect 501294 149940 501322 150198
rect 501938 149940 501966 150198
rect 502340 150204 502392 150210
rect 502536 150198 502610 150226
rect 503732 150210 503760 156606
rect 503824 150226 503852 163254
rect 504100 163146 504128 163254
rect 504178 163200 504234 164400
rect 505006 163200 505062 164400
rect 505112 163254 505784 163282
rect 504192 163146 504220 163200
rect 504100 163118 504220 163146
rect 505020 156670 505048 163200
rect 505008 156664 505060 156670
rect 505008 156606 505060 156612
rect 505112 150226 505140 163254
rect 505756 163146 505784 163254
rect 505834 163200 505890 164400
rect 506754 163200 506810 164400
rect 507582 163200 507638 164400
rect 508410 163200 508466 164400
rect 509238 163200 509294 164400
rect 509344 163254 509556 163282
rect 505848 163146 505876 163200
rect 505756 163118 505876 163146
rect 505284 158840 505336 158846
rect 505284 158782 505336 158788
rect 502340 150146 502392 150152
rect 502582 149940 502610 150198
rect 503214 150204 503266 150210
rect 503214 150146 503266 150152
rect 503720 150204 503772 150210
rect 503824 150198 503898 150226
rect 503720 150146 503772 150152
rect 503226 149940 503254 150146
rect 503870 149940 503898 150198
rect 504502 150204 504554 150210
rect 505112 150198 505186 150226
rect 505296 150210 505324 158782
rect 506768 158778 506796 163200
rect 507596 158846 507624 163200
rect 508320 158908 508372 158914
rect 508320 158850 508372 158856
rect 507584 158840 507636 158846
rect 507584 158782 507636 158788
rect 505744 158772 505796 158778
rect 505744 158714 505796 158720
rect 506756 158772 506808 158778
rect 506756 158714 506808 158720
rect 507032 158772 507084 158778
rect 507032 158714 507084 158720
rect 505756 150226 505784 158714
rect 507044 150226 507072 158714
rect 507768 151904 507820 151910
rect 507768 151846 507820 151852
rect 507780 150226 507808 151846
rect 504502 150146 504554 150152
rect 504514 149940 504542 150146
rect 505158 149940 505186 150198
rect 505284 150204 505336 150210
rect 505756 150198 505830 150226
rect 505284 150146 505336 150152
rect 505802 149940 505830 150198
rect 506434 150204 506486 150210
rect 507044 150198 507118 150226
rect 506434 150146 506486 150152
rect 506446 149940 506474 150146
rect 507090 149940 507118 150198
rect 507734 150198 507808 150226
rect 508332 150226 508360 158850
rect 508424 158778 508452 163200
rect 509252 163146 509280 163200
rect 509344 163146 509372 163254
rect 509252 163118 509372 163146
rect 508412 158772 508464 158778
rect 508412 158714 508464 158720
rect 509424 158772 509476 158778
rect 509424 158714 509476 158720
rect 509056 151972 509108 151978
rect 509056 151914 509108 151920
rect 509068 150226 509096 151914
rect 509436 151814 509464 158714
rect 509528 151910 509556 163254
rect 510066 163200 510122 164400
rect 510894 163200 510950 164400
rect 511722 163200 511778 164400
rect 512012 163254 512592 163282
rect 510080 158914 510108 163200
rect 510068 158908 510120 158914
rect 510068 158850 510120 158856
rect 510344 152856 510396 152862
rect 510344 152798 510396 152804
rect 509516 151904 509568 151910
rect 509516 151846 509568 151852
rect 509436 151786 509648 151814
rect 508332 150198 508406 150226
rect 507734 149940 507762 150198
rect 508378 149940 508406 150198
rect 509022 150198 509096 150226
rect 509620 150226 509648 151786
rect 510356 150226 510384 152798
rect 510908 151978 510936 163200
rect 511736 158778 511764 163200
rect 511724 158772 511776 158778
rect 511724 158714 511776 158720
rect 510988 153128 511040 153134
rect 510988 153070 511040 153076
rect 510896 151972 510948 151978
rect 510896 151914 510948 151920
rect 511000 150226 511028 153070
rect 511632 153060 511684 153066
rect 511632 153002 511684 153008
rect 511644 150226 511672 153002
rect 512012 152862 512040 163254
rect 512564 163146 512592 163254
rect 512642 163200 512698 164400
rect 513470 163200 513526 164400
rect 514298 163200 514354 164400
rect 514864 163254 515076 163282
rect 512656 163146 512684 163200
rect 512564 163118 512684 163146
rect 512276 153196 512328 153202
rect 512276 153138 512328 153144
rect 512000 152856 512052 152862
rect 512000 152798 512052 152804
rect 512288 150226 512316 153138
rect 513484 153134 513512 163200
rect 513472 153128 513524 153134
rect 513472 153070 513524 153076
rect 513564 153128 513616 153134
rect 513564 153070 513616 153076
rect 512920 152992 512972 152998
rect 512920 152934 512972 152940
rect 512932 150226 512960 152934
rect 513576 150226 513604 153070
rect 514312 153066 514340 163200
rect 514864 153202 514892 163254
rect 515048 163146 515076 163254
rect 515126 163200 515182 164400
rect 515954 163200 516010 164400
rect 516152 163254 516732 163282
rect 515140 163146 515168 163200
rect 515048 163118 515168 163146
rect 514944 158772 514996 158778
rect 514944 158714 514996 158720
rect 514852 153196 514904 153202
rect 514852 153138 514904 153144
rect 514300 153060 514352 153066
rect 514300 153002 514352 153008
rect 514208 152924 514260 152930
rect 514208 152866 514260 152872
rect 514220 150226 514248 152866
rect 514956 151814 514984 158714
rect 515968 152998 515996 163200
rect 516152 153134 516180 163254
rect 516704 163146 516732 163254
rect 516782 163200 516838 164400
rect 517610 163200 517666 164400
rect 518530 163200 518586 164400
rect 519004 163254 519308 163282
rect 516796 163146 516824 163200
rect 516704 163118 516824 163146
rect 517624 161474 517652 163200
rect 517532 161446 517652 161474
rect 517532 158794 517560 161446
rect 517440 158766 517560 158794
rect 518544 158778 518572 163200
rect 518808 159452 518860 159458
rect 518808 159394 518860 159400
rect 518716 159384 518768 159390
rect 518716 159326 518768 159332
rect 518532 158772 518584 158778
rect 516140 153128 516192 153134
rect 516140 153070 516192 153076
rect 515956 152992 516008 152998
rect 515956 152934 516008 152940
rect 517440 152930 517468 158766
rect 518532 158714 518584 158720
rect 517428 152924 517480 152930
rect 517428 152866 517480 152872
rect 516692 152108 516744 152114
rect 516692 152050 516744 152056
rect 516048 151904 516100 151910
rect 516048 151846 516100 151852
rect 514864 151786 514984 151814
rect 515496 151836 515548 151842
rect 514864 150226 514892 151786
rect 515496 151778 515548 151784
rect 515508 150226 515536 151778
rect 509620 150198 509694 150226
rect 509022 149940 509050 150198
rect 509666 149940 509694 150198
rect 510310 150198 510384 150226
rect 510954 150198 511028 150226
rect 511598 150198 511672 150226
rect 512242 150198 512316 150226
rect 512886 150198 512960 150226
rect 513530 150198 513604 150226
rect 514174 150198 514248 150226
rect 514818 150198 514892 150226
rect 515462 150198 515536 150226
rect 516060 150226 516088 151846
rect 516704 150226 516732 152050
rect 517428 151972 517480 151978
rect 517428 151914 517480 151920
rect 517440 150226 517468 151914
rect 518728 150226 518756 159326
rect 516060 150198 516134 150226
rect 516704 150198 516778 150226
rect 510310 149940 510338 150198
rect 510954 149940 510982 150198
rect 511598 149940 511626 150198
rect 512242 149940 512270 150198
rect 512886 149940 512914 150198
rect 513530 149940 513558 150198
rect 514174 149940 514202 150198
rect 514818 149940 514846 150198
rect 515462 149940 515490 150198
rect 516106 149940 516134 150198
rect 516750 149940 516778 150198
rect 517394 150198 517468 150226
rect 518026 150204 518078 150210
rect 517394 149940 517422 150198
rect 518026 150146 518078 150152
rect 518682 150198 518756 150226
rect 518820 150210 518848 159394
rect 519004 151842 519032 163254
rect 519280 163146 519308 163254
rect 519358 163200 519414 164400
rect 519924 163254 520136 163282
rect 519372 163146 519400 163200
rect 519280 163118 519400 163146
rect 519726 163160 519782 163169
rect 519726 163095 519782 163104
rect 519542 161664 519598 161673
rect 519542 161599 519598 161608
rect 518992 151836 519044 151842
rect 518992 151778 519044 151784
rect 519450 151192 519506 151201
rect 519450 151127 519506 151136
rect 518808 150204 518860 150210
rect 518038 149940 518066 150146
rect 518682 149940 518710 150198
rect 518808 150146 518860 150152
rect 519358 140584 519414 140593
rect 519358 140519 519414 140528
rect 117240 132518 117360 132546
rect 117332 132410 117360 132518
rect 117240 132382 117360 132410
rect 117240 127945 117268 132382
rect 519372 128897 519400 140519
rect 519464 138417 519492 151127
rect 519556 147937 519584 161599
rect 519634 160168 519690 160177
rect 519634 160103 519690 160112
rect 519542 147928 519598 147937
rect 519542 147863 519598 147872
rect 519648 146577 519676 160103
rect 519740 149297 519768 163095
rect 519818 157176 519874 157185
rect 519818 157111 519874 157120
rect 519726 149288 519782 149297
rect 519726 149223 519782 149232
rect 519726 148200 519782 148209
rect 519726 148135 519782 148144
rect 519634 146568 519690 146577
rect 519634 146503 519690 146512
rect 519634 145208 519690 145217
rect 519634 145143 519690 145152
rect 519542 142216 519598 142225
rect 519542 142151 519598 142160
rect 519450 138408 519506 138417
rect 519450 138343 519506 138352
rect 519450 136096 519506 136105
rect 519450 136031 519506 136040
rect 519358 128888 519414 128897
rect 519358 128823 519414 128832
rect 117226 127936 117282 127945
rect 117226 127871 117282 127880
rect 519464 124817 519492 136031
rect 519556 130257 519584 142151
rect 519648 132977 519676 145143
rect 519740 135697 519768 148135
rect 519832 143857 519860 157111
rect 519924 151910 519952 163254
rect 520108 163146 520136 163254
rect 520186 163200 520242 164400
rect 520292 163254 520964 163282
rect 520200 163146 520228 163200
rect 520108 163118 520228 163146
rect 520186 158672 520242 158681
rect 520186 158607 520242 158616
rect 520094 155680 520150 155689
rect 520094 155615 520150 155624
rect 520002 154184 520058 154193
rect 520002 154119 520058 154128
rect 519912 151904 519964 151910
rect 519912 151846 519964 151852
rect 519910 149696 519966 149705
rect 519910 149631 519966 149640
rect 519818 143848 519874 143857
rect 519818 143783 519874 143792
rect 519924 137057 519952 149631
rect 520016 141137 520044 154119
rect 520108 142497 520136 155615
rect 520200 145353 520228 158607
rect 520292 152114 520320 163254
rect 520936 163146 520964 163254
rect 521014 163200 521070 164400
rect 521842 163200 521898 164400
rect 522670 163200 522726 164400
rect 523498 163200 523554 164400
rect 521028 163146 521056 163200
rect 520936 163118 521056 163146
rect 521856 161474 521884 163200
rect 521672 161446 521884 161474
rect 521672 158794 521700 161446
rect 522684 159458 522712 163200
rect 522672 159452 522724 159458
rect 522672 159394 522724 159400
rect 523512 159390 523540 163200
rect 523500 159384 523552 159390
rect 523500 159326 523552 159332
rect 521580 158766 521700 158794
rect 521014 152688 521070 152697
rect 521014 152623 521070 152632
rect 520280 152108 520332 152114
rect 520280 152050 520332 152056
rect 520186 145344 520242 145353
rect 520186 145279 520242 145288
rect 520922 143712 520978 143721
rect 520922 143647 520978 143656
rect 520094 142488 520150 142497
rect 520094 142423 520150 142432
rect 520002 141128 520058 141137
rect 520002 141063 520058 141072
rect 520002 139088 520058 139097
rect 520002 139023 520058 139032
rect 519910 137048 519966 137057
rect 519910 136983 519966 136992
rect 519726 135688 519782 135697
rect 519726 135623 519782 135632
rect 519818 133104 519874 133113
rect 519818 133039 519874 133048
rect 519634 132968 519690 132977
rect 519634 132903 519690 132912
rect 519542 130248 519598 130257
rect 519542 130183 519598 130192
rect 519726 130112 519782 130121
rect 519726 130047 519782 130056
rect 519634 128616 519690 128625
rect 519634 128551 519690 128560
rect 519542 127120 519598 127129
rect 519542 127055 519598 127064
rect 519450 124808 519506 124817
rect 519450 124743 519506 124752
rect 519266 124128 519322 124137
rect 519266 124063 519322 124072
rect 519280 113937 519308 124063
rect 519358 122632 519414 122641
rect 519358 122567 519414 122576
rect 519266 113928 519322 113937
rect 519266 113863 519322 113872
rect 519372 112577 519400 122567
rect 519450 119640 519506 119649
rect 519450 119575 519506 119584
rect 519358 112568 519414 112577
rect 519358 112503 519414 112512
rect 519464 109857 519492 119575
rect 519556 116657 519584 127055
rect 519648 118017 519676 128551
rect 519740 119377 519768 130047
rect 519832 122097 519860 133039
rect 519910 131608 519966 131617
rect 519910 131543 519966 131552
rect 519818 122088 519874 122097
rect 519818 122023 519874 122032
rect 519924 120737 519952 131543
rect 520016 127537 520044 139023
rect 520186 137592 520242 137601
rect 520186 137527 520242 137536
rect 520094 134600 520150 134609
rect 520094 134535 520150 134544
rect 520002 127528 520058 127537
rect 520002 127463 520058 127472
rect 520002 125624 520058 125633
rect 520002 125559 520058 125568
rect 519910 120728 519966 120737
rect 519910 120663 519966 120672
rect 519726 119368 519782 119377
rect 519726 119303 519782 119312
rect 519818 118144 519874 118153
rect 519818 118079 519874 118088
rect 519634 118008 519690 118017
rect 519634 117943 519690 117952
rect 519542 116648 519598 116657
rect 519542 116583 519598 116592
rect 519726 113520 519782 113529
rect 519726 113455 519782 113464
rect 519634 112024 519690 112033
rect 519634 111959 519690 111968
rect 519542 110528 519598 110537
rect 519542 110463 519598 110472
rect 519450 109848 519506 109857
rect 519450 109783 519506 109792
rect 117134 104816 117190 104825
rect 117134 104751 117190 104760
rect 519556 101697 519584 110463
rect 519648 103057 519676 111959
rect 519740 104417 519768 113455
rect 519832 108497 519860 118079
rect 519910 116512 519966 116521
rect 519910 116447 519966 116456
rect 519818 108488 519874 108497
rect 519818 108423 519874 108432
rect 519924 107137 519952 116447
rect 520016 115297 520044 125559
rect 520108 123457 520136 134535
rect 520200 126177 520228 137527
rect 520936 131753 520964 143647
rect 521028 139777 521056 152623
rect 521580 151978 521608 158766
rect 521568 151972 521620 151978
rect 521568 151914 521620 151920
rect 521106 146704 521162 146713
rect 521106 146639 521162 146648
rect 521014 139768 521070 139777
rect 521014 139703 521070 139712
rect 521120 134337 521148 146639
rect 521106 134328 521162 134337
rect 521106 134263 521162 134272
rect 520922 131744 520978 131753
rect 520922 131679 520978 131688
rect 520186 126168 520242 126177
rect 520186 126103 520242 126112
rect 520094 123448 520150 123457
rect 520094 123383 520150 123392
rect 520094 121136 520150 121145
rect 520094 121071 520150 121080
rect 520002 115288 520058 115297
rect 520002 115223 520058 115232
rect 520108 111217 520136 121071
rect 520186 115016 520242 115025
rect 520186 114951 520242 114960
rect 520094 111208 520150 111217
rect 520094 111143 520150 111152
rect 519910 107128 519966 107137
rect 519910 107063 519966 107072
rect 520200 105777 520228 114951
rect 521290 109032 521346 109041
rect 521290 108967 521346 108976
rect 521106 107536 521162 107545
rect 521106 107471 521162 107480
rect 520278 106040 520334 106049
rect 520278 105975 520334 105984
rect 520186 105768 520242 105777
rect 520186 105703 520242 105712
rect 519726 104408 519782 104417
rect 519726 104343 519782 104352
rect 519634 103048 519690 103057
rect 519634 102983 519690 102992
rect 519542 101688 519598 101697
rect 519542 101623 519598 101632
rect 117042 101008 117098 101017
rect 117042 100943 117098 100952
rect 116858 99104 116914 99113
rect 116858 99039 116914 99048
rect 520292 97617 520320 105975
rect 521014 104544 521070 104553
rect 521014 104479 521070 104488
rect 520922 101552 520978 101561
rect 520922 101487 520978 101496
rect 520278 97608 520334 97617
rect 520278 97543 520334 97552
rect 116766 97200 116822 97209
rect 116766 97135 116822 97144
rect 520278 95568 520334 95577
rect 520278 95503 520334 95512
rect 116674 95296 116730 95305
rect 116674 95231 116730 95240
rect 116582 93392 116638 93401
rect 116582 93327 116638 93336
rect 116124 92472 116176 92478
rect 116124 92414 116176 92420
rect 519634 92440 519690 92449
rect 116136 91361 116164 92414
rect 519634 92375 519690 92384
rect 116122 91352 116178 91361
rect 116122 91287 116178 91296
rect 116124 89684 116176 89690
rect 116124 89626 116176 89632
rect 116136 89457 116164 89626
rect 116122 89448 116178 89457
rect 116122 89383 116178 89392
rect 116032 88324 116084 88330
rect 116032 88266 116084 88272
rect 116044 87553 116072 88266
rect 116030 87544 116086 87553
rect 116030 87479 116086 87488
rect 115202 85640 115258 85649
rect 115202 85575 115258 85584
rect 519648 85377 519676 92375
rect 520002 90944 520058 90953
rect 520002 90879 520058 90888
rect 519726 89448 519782 89457
rect 519726 89383 519782 89392
rect 519634 85368 519690 85377
rect 519634 85303 519690 85312
rect 519082 84960 519138 84969
rect 519082 84895 519138 84904
rect 116584 83972 116636 83978
rect 116584 83914 116636 83920
rect 116596 83745 116624 83914
rect 116582 83736 116638 83745
rect 116582 83671 116638 83680
rect 116216 82816 116268 82822
rect 116216 82758 116268 82764
rect 116228 81841 116256 82758
rect 116214 81832 116270 81841
rect 116214 81767 116270 81776
rect 115940 80028 115992 80034
rect 115940 79970 115992 79976
rect 115952 79937 115980 79970
rect 115938 79928 115994 79937
rect 115938 79863 115994 79872
rect 114192 78668 114244 78674
rect 114192 78610 114244 78616
rect 116124 78668 116176 78674
rect 116124 78610 116176 78616
rect 116136 78033 116164 78610
rect 519096 78577 519124 84895
rect 519740 82657 519768 89383
rect 519910 87952 519966 87961
rect 519910 87887 519966 87896
rect 519818 86456 519874 86465
rect 519818 86391 519874 86400
rect 519726 82648 519782 82657
rect 519726 82583 519782 82592
rect 519450 81968 519506 81977
rect 519450 81903 519506 81912
rect 519082 78568 519138 78577
rect 519082 78503 519138 78512
rect 116122 78024 116178 78033
rect 116122 77959 116178 77968
rect 519464 75993 519492 81903
rect 519832 79937 519860 86391
rect 519924 81297 519952 87887
rect 520016 84017 520044 90879
rect 520292 88097 520320 95503
rect 520936 93537 520964 101487
rect 521028 96257 521056 104479
rect 521120 98977 521148 107471
rect 521198 103048 521254 103057
rect 521198 102983 521254 102992
rect 521106 98968 521162 98977
rect 521106 98903 521162 98912
rect 521014 96248 521070 96257
rect 521014 96183 521070 96192
rect 521212 94897 521240 102983
rect 521304 100337 521332 108967
rect 521290 100328 521346 100337
rect 521290 100263 521346 100272
rect 521474 100056 521530 100065
rect 521474 99991 521530 100000
rect 521290 98560 521346 98569
rect 521290 98495 521346 98504
rect 521198 94888 521254 94897
rect 521198 94823 521254 94832
rect 521014 93936 521070 93945
rect 521014 93871 521070 93880
rect 520922 93528 520978 93537
rect 520922 93463 520978 93472
rect 520278 88088 520334 88097
rect 520278 88023 520334 88032
rect 521028 86737 521056 93871
rect 521304 90817 521332 98495
rect 521382 97064 521438 97073
rect 521382 96999 521438 97008
rect 521290 90808 521346 90817
rect 521290 90743 521346 90752
rect 521396 89593 521424 96999
rect 521488 92177 521516 99991
rect 521474 92168 521530 92177
rect 521474 92103 521530 92112
rect 521382 89584 521438 89593
rect 521382 89519 521438 89528
rect 521014 86728 521070 86737
rect 521014 86663 521070 86672
rect 520002 84008 520058 84017
rect 520002 83943 520058 83952
rect 520094 83464 520150 83473
rect 520094 83399 520150 83408
rect 519910 81288 519966 81297
rect 519910 81223 519966 81232
rect 519818 79928 519874 79937
rect 519818 79863 519874 79872
rect 520002 78976 520058 78985
rect 520002 78911 520058 78920
rect 519818 77480 519874 77489
rect 519818 77415 519874 77424
rect 519450 75984 519506 75993
rect 519450 75919 519506 75928
rect 116674 74080 116730 74089
rect 116674 74015 116730 74024
rect 116582 72176 116638 72185
rect 116582 72111 116638 72120
rect 116596 71806 116624 72111
rect 114192 71800 114244 71806
rect 114192 71742 114244 71748
rect 116584 71800 116636 71806
rect 116584 71742 116636 71748
rect 114100 69080 114152 69086
rect 114100 69022 114152 69028
rect 114008 67652 114060 67658
rect 114008 67594 114060 67600
rect 113916 66292 113968 66298
rect 113916 66234 113968 66240
rect 113364 64728 113416 64734
rect 113364 64670 113416 64676
rect 113376 64569 113404 64670
rect 113362 64560 113418 64569
rect 113362 64495 113418 64504
rect 113824 63572 113876 63578
rect 113824 63514 113876 63520
rect 112444 62144 112496 62150
rect 112444 62086 112496 62092
rect 110326 53952 110382 53961
rect 109696 53910 110326 53938
rect 109696 12434 109724 53910
rect 110326 53887 110382 53896
rect 110326 52592 110382 52601
rect 110326 52527 110382 52536
rect 110340 51218 110368 52527
rect 110340 51190 110460 51218
rect 110326 51096 110382 51105
rect 109512 12406 109724 12434
rect 109788 51054 110326 51082
rect 109512 3913 109540 12406
rect 109788 8242 109816 51054
rect 110326 51031 110382 51040
rect 110432 50946 110460 51190
rect 109604 8214 109816 8242
rect 109880 50918 110460 50946
rect 109498 3904 109554 3913
rect 109498 3839 109554 3848
rect 109498 3496 109554 3505
rect 109498 3431 109554 3440
rect 32402 2680 32458 2689
rect 36358 2680 36414 2689
rect 36018 2638 36358 2666
rect 32402 2615 32458 2624
rect 36358 2615 36414 2624
rect 62394 2680 62450 2689
rect 62394 2615 62450 2624
rect 64142 2680 64198 2689
rect 64142 2615 64198 2624
rect 65338 2680 65394 2689
rect 65338 2615 65394 2624
rect 68006 2680 68062 2689
rect 68006 2615 68062 2624
rect 68282 2680 68338 2689
rect 68282 2615 68338 2624
rect 68466 2680 68522 2689
rect 68466 2615 68522 2624
rect 69386 2680 69442 2689
rect 69386 2615 69442 2624
rect 75642 2680 75698 2689
rect 77482 2680 77538 2689
rect 75642 2615 75698 2624
rect 77220 2638 77482 2666
rect 29550 2408 29606 2417
rect 29302 2366 29550 2394
rect 29550 2343 29606 2352
rect 26054 2272 26110 2281
rect 25990 2230 26054 2258
rect 26054 2207 26110 2216
rect 22926 2136 22982 2145
rect 2700 1290 2728 2108
rect 6012 1737 6040 2108
rect 5998 1728 6054 1737
rect 5998 1663 6054 1672
rect 9324 1465 9352 2108
rect 12636 1601 12664 2108
rect 15948 1873 15976 2108
rect 19366 2094 19656 2122
rect 22678 2094 22926 2122
rect 19628 2009 19656 2094
rect 22926 2071 22982 2080
rect 19614 2000 19670 2009
rect 19614 1935 19670 1944
rect 15934 1864 15990 1873
rect 15934 1799 15990 1808
rect 12622 1592 12678 1601
rect 12622 1527 12678 1536
rect 9310 1456 9366 1465
rect 9310 1391 9366 1400
rect 2688 1284 2740 1290
rect 2688 1226 2740 1232
rect 32416 762 32444 2615
rect 33046 2544 33102 2553
rect 32706 2502 33046 2530
rect 33046 2479 33102 2488
rect 39316 1222 39344 2108
rect 42628 1494 42656 2108
rect 42616 1488 42668 1494
rect 42616 1430 42668 1436
rect 46032 1426 46060 2108
rect 46020 1420 46072 1426
rect 46020 1362 46072 1368
rect 39304 1216 39356 1222
rect 39304 1158 39356 1164
rect 49344 1154 49372 2108
rect 49332 1148 49384 1154
rect 49332 1090 49384 1096
rect 52656 1086 52684 2108
rect 55968 1358 55996 2108
rect 59372 1630 59400 2108
rect 62408 1902 62436 2615
rect 62396 1896 62448 1902
rect 62396 1838 62448 1844
rect 62684 1766 62712 2108
rect 64156 1834 64184 2615
rect 65352 1902 65380 2615
rect 65340 1896 65392 1902
rect 65340 1838 65392 1844
rect 64144 1828 64196 1834
rect 64144 1770 64196 1776
rect 62672 1760 62724 1766
rect 62672 1702 62724 1708
rect 59360 1624 59412 1630
rect 59360 1566 59412 1572
rect 55956 1352 56008 1358
rect 55956 1294 56008 1300
rect 52644 1080 52696 1086
rect 52644 1022 52696 1028
rect 65996 1018 66024 2108
rect 68020 1902 68048 2615
rect 68008 1896 68060 1902
rect 68008 1838 68060 1844
rect 68296 1494 68324 2615
rect 68480 1630 68508 2615
rect 69308 1698 69336 2108
rect 69400 1834 69428 2615
rect 69388 1828 69440 1834
rect 69388 1770 69440 1776
rect 69296 1692 69348 1698
rect 69296 1634 69348 1640
rect 68468 1624 68520 1630
rect 68468 1566 68520 1572
rect 72712 1562 72740 2108
rect 75656 1834 75684 2615
rect 75644 1828 75696 1834
rect 75644 1770 75696 1776
rect 72700 1556 72752 1562
rect 72700 1498 72752 1504
rect 68284 1488 68336 1494
rect 68284 1430 68336 1436
rect 65984 1012 66036 1018
rect 65984 954 66036 960
rect 76024 950 76052 2108
rect 77220 1766 77248 2638
rect 77482 2615 77538 2624
rect 85394 2680 85450 2689
rect 85394 2615 85450 2624
rect 86682 2680 86738 2689
rect 86682 2615 86738 2624
rect 91742 2680 91798 2689
rect 93030 2680 93086 2689
rect 92690 2638 93030 2666
rect 91742 2615 91798 2624
rect 93030 2615 93086 2624
rect 98918 2680 98974 2689
rect 99194 2680 99250 2689
rect 98974 2638 99194 2666
rect 98918 2615 98974 2624
rect 99194 2615 99250 2624
rect 99562 2680 99618 2689
rect 99562 2615 99618 2624
rect 99746 2680 99802 2689
rect 103426 2680 103482 2689
rect 99746 2615 99802 2624
rect 102796 2638 103426 2666
rect 77208 1760 77260 1766
rect 77208 1702 77260 1708
rect 79336 1630 79364 2108
rect 82648 1766 82676 2108
rect 85408 1834 85436 2615
rect 86052 1834 86080 2108
rect 85396 1828 85448 1834
rect 85396 1770 85448 1776
rect 86040 1828 86092 1834
rect 86040 1770 86092 1776
rect 82636 1760 82688 1766
rect 82636 1702 82688 1708
rect 79324 1624 79376 1630
rect 79324 1566 79376 1572
rect 86696 1329 86724 2615
rect 91650 2544 91706 2553
rect 91650 2479 91706 2488
rect 91664 2145 91692 2479
rect 87970 2136 88026 2145
rect 91650 2136 91706 2145
rect 87970 2071 88026 2080
rect 87984 1494 88012 2071
rect 89364 1902 89392 2108
rect 91650 2071 91706 2080
rect 89260 1896 89312 1902
rect 89260 1838 89312 1844
rect 89352 1896 89404 1902
rect 89352 1838 89404 1844
rect 87972 1488 88024 1494
rect 87972 1430 88024 1436
rect 86682 1320 86738 1329
rect 86682 1255 86738 1264
rect 89272 1193 89300 1838
rect 89258 1184 89314 1193
rect 89258 1119 89314 1128
rect 76012 944 76064 950
rect 32692 870 32812 898
rect 76012 886 76064 892
rect 91756 882 91784 2615
rect 95698 2544 95754 2553
rect 96342 2544 96398 2553
rect 96002 2502 96342 2530
rect 95698 2479 95754 2488
rect 96342 2479 96398 2488
rect 32692 762 32720 870
rect 32784 800 32812 870
rect 91744 876 91796 882
rect 91744 818 91796 824
rect 95712 814 95740 2479
rect 97172 1896 97224 1902
rect 97172 1838 97224 1844
rect 97184 1494 97212 1838
rect 99392 1630 99420 2108
rect 97264 1624 97316 1630
rect 97264 1566 97316 1572
rect 99380 1624 99432 1630
rect 99380 1566 99432 1572
rect 97276 1494 97304 1566
rect 97172 1488 97224 1494
rect 97172 1430 97224 1436
rect 97264 1488 97316 1494
rect 97264 1430 97316 1436
rect 98274 1184 98330 1193
rect 98274 1119 98330 1128
rect 95700 808 95752 814
rect 32416 734 32720 762
rect 32770 -400 32826 800
rect 98288 800 98316 1119
rect 99576 814 99604 2615
rect 99760 882 99788 2615
rect 99838 2544 99894 2553
rect 99838 2479 99894 2488
rect 99852 1057 99880 2479
rect 102704 1698 102732 2108
rect 102600 1692 102652 1698
rect 102600 1634 102652 1640
rect 102692 1692 102744 1698
rect 102692 1634 102744 1640
rect 102612 1578 102640 1634
rect 102796 1578 102824 2638
rect 103426 2615 103482 2624
rect 104162 2544 104218 2553
rect 104162 2479 104218 2488
rect 104176 2145 104204 2479
rect 104162 2136 104218 2145
rect 104162 2071 104218 2080
rect 104346 2136 104402 2145
rect 106030 2094 106228 2122
rect 104346 2071 104402 2080
rect 104360 1902 104388 2071
rect 104348 1896 104400 1902
rect 104532 1896 104584 1902
rect 104348 1838 104400 1844
rect 104452 1856 104532 1884
rect 104072 1760 104124 1766
rect 104452 1714 104480 1856
rect 104532 1838 104584 1844
rect 105728 1896 105780 1902
rect 105728 1838 105780 1844
rect 105820 1896 105872 1902
rect 105820 1838 105872 1844
rect 105912 1896 105964 1902
rect 105912 1838 105964 1844
rect 104124 1708 104480 1714
rect 104072 1702 104480 1708
rect 104084 1686 104480 1702
rect 102612 1550 102824 1578
rect 105740 1476 105768 1838
rect 105832 1698 105860 1838
rect 105820 1692 105872 1698
rect 105820 1634 105872 1640
rect 105924 1630 105952 1838
rect 106200 1698 106228 2094
rect 109328 1902 109356 2108
rect 109224 1896 109276 1902
rect 109224 1838 109276 1844
rect 109316 1896 109368 1902
rect 109316 1838 109368 1844
rect 106188 1692 106240 1698
rect 106188 1634 106240 1640
rect 105912 1624 105964 1630
rect 105912 1566 105964 1572
rect 106004 1624 106056 1630
rect 106004 1566 106056 1572
rect 106016 1476 106044 1566
rect 105740 1448 106044 1476
rect 108212 1488 108264 1494
rect 108212 1430 108264 1436
rect 108304 1488 108356 1494
rect 108304 1430 108356 1436
rect 103486 1366 103928 1394
rect 103334 1320 103390 1329
rect 103486 1306 103514 1366
rect 103390 1278 103514 1306
rect 103334 1255 103390 1264
rect 99838 1048 99894 1057
rect 99838 983 99894 992
rect 103900 882 103928 1366
rect 108224 1329 108252 1430
rect 108210 1320 108266 1329
rect 108210 1255 108266 1264
rect 108316 882 108344 1430
rect 109236 1170 109264 1838
rect 109512 1737 109540 3431
rect 109604 1834 109632 8214
rect 109880 3641 109908 50918
rect 110326 48376 110382 48385
rect 109972 48334 110326 48362
rect 109866 3632 109922 3641
rect 109866 3567 109922 3576
rect 109866 2816 109922 2825
rect 109866 2751 109922 2760
rect 109592 1828 109644 1834
rect 109592 1770 109644 1776
rect 109498 1728 109554 1737
rect 109498 1663 109554 1672
rect 109880 1442 109908 2751
rect 109972 1766 110000 48334
rect 110326 48311 110382 48320
rect 110326 47152 110382 47161
rect 110326 47087 110382 47096
rect 110340 45554 110368 47087
rect 110064 45526 110368 45554
rect 110064 7290 110092 45526
rect 110326 44296 110382 44305
rect 110156 44254 110326 44282
rect 110156 8106 110184 44254
rect 110326 44231 110382 44240
rect 110326 41440 110382 41449
rect 110326 41375 110382 41384
rect 110340 35894 110368 41375
rect 110248 35866 110368 35894
rect 110248 8242 110276 35866
rect 110326 34640 110382 34649
rect 110326 34575 110382 34584
rect 110340 8378 110368 34575
rect 110340 8350 110736 8378
rect 110326 8256 110382 8265
rect 110248 8214 110326 8242
rect 110326 8191 110382 8200
rect 110510 8256 110566 8265
rect 110510 8191 110566 8200
rect 110156 8078 110276 8106
rect 110064 7262 110184 7290
rect 110156 3074 110184 7262
rect 110248 4026 110276 8078
rect 110248 3998 110368 4026
rect 110234 3904 110290 3913
rect 110234 3839 110290 3848
rect 110248 3505 110276 3839
rect 110234 3496 110290 3505
rect 110234 3431 110290 3440
rect 110064 3046 110184 3074
rect 109960 1760 110012 1766
rect 109960 1702 110012 1708
rect 110064 1630 110092 3046
rect 110142 2952 110198 2961
rect 110142 2887 110198 2896
rect 110052 1624 110104 1630
rect 110052 1566 110104 1572
rect 109788 1414 109908 1442
rect 109788 1306 109816 1414
rect 109604 1278 109816 1306
rect 109604 1170 109632 1278
rect 110156 1193 110184 2887
rect 110340 2836 110368 3998
rect 110248 2808 110368 2836
rect 110248 1329 110276 2808
rect 110524 1562 110552 8191
rect 110602 5672 110658 5681
rect 110602 5607 110658 5616
rect 110616 2825 110644 5607
rect 110708 3233 110736 8350
rect 111062 7984 111118 7993
rect 111062 7919 111118 7928
rect 110694 3224 110750 3233
rect 110694 3159 110750 3168
rect 110602 2816 110658 2825
rect 110602 2751 110658 2760
rect 111076 1970 111104 7919
rect 111706 2952 111762 2961
rect 111706 2887 111762 2896
rect 111720 2854 111748 2887
rect 111708 2848 111760 2854
rect 111708 2790 111760 2796
rect 111064 1964 111116 1970
rect 111064 1906 111116 1912
rect 112456 1766 112484 62086
rect 112536 42832 112588 42838
rect 112536 42774 112588 42780
rect 112444 1760 112496 1766
rect 112444 1702 112496 1708
rect 110512 1556 110564 1562
rect 110512 1498 110564 1504
rect 110234 1320 110290 1329
rect 110234 1255 110290 1264
rect 109236 1142 109632 1170
rect 110142 1184 110198 1193
rect 110142 1119 110198 1128
rect 112548 950 112576 42774
rect 113836 7721 113864 63514
rect 113928 19009 113956 66234
rect 114020 30433 114048 67594
rect 114112 41857 114140 69022
rect 114204 53145 114232 71742
rect 116306 70272 116362 70281
rect 116306 70207 116362 70216
rect 116320 69086 116348 70207
rect 116308 69080 116360 69086
rect 116308 69022 116360 69028
rect 116122 68368 116178 68377
rect 116122 68303 116178 68312
rect 116136 67658 116164 68303
rect 116124 67652 116176 67658
rect 116124 67594 116176 67600
rect 116582 66464 116638 66473
rect 116582 66399 116638 66408
rect 116596 66298 116624 66399
rect 116584 66292 116636 66298
rect 116584 66234 116636 66240
rect 116688 64874 116716 74015
rect 519832 71913 519860 77415
rect 519910 75984 519966 75993
rect 519910 75919 519966 75928
rect 519818 71904 519874 71913
rect 519818 71839 519874 71848
rect 519924 70553 519952 75919
rect 520016 73273 520044 78911
rect 520108 77217 520136 83399
rect 520186 80472 520242 80481
rect 520186 80407 520242 80416
rect 520094 77208 520150 77217
rect 520094 77143 520150 77152
rect 520200 74633 520228 80407
rect 520186 74624 520242 74633
rect 520186 74559 520242 74568
rect 521106 74488 521162 74497
rect 521106 74423 521162 74432
rect 520002 73264 520058 73273
rect 520002 73199 520058 73208
rect 520922 72992 520978 73001
rect 520922 72927 520978 72936
rect 519910 70544 519966 70553
rect 519910 70479 519966 70488
rect 520936 67833 520964 72927
rect 521014 69864 521070 69873
rect 521014 69799 521070 69808
rect 520922 67824 520978 67833
rect 520922 67759 520978 67768
rect 520462 66872 520518 66881
rect 520462 66807 520518 66816
rect 520370 65376 520426 65385
rect 520370 65311 520426 65320
rect 116596 64846 116716 64874
rect 116596 64734 116624 64846
rect 116584 64728 116636 64734
rect 116584 64670 116636 64676
rect 116214 64560 116270 64569
rect 116214 64495 116270 64504
rect 116228 63578 116256 64495
rect 116216 63572 116268 63578
rect 116216 63514 116268 63520
rect 116122 62656 116178 62665
rect 116122 62591 116178 62600
rect 116136 62150 116164 62591
rect 116124 62144 116176 62150
rect 116124 62086 116176 62092
rect 520384 61033 520412 65311
rect 520476 62393 520504 66807
rect 521028 65113 521056 69799
rect 521120 69193 521148 74423
rect 521198 71496 521254 71505
rect 521198 71431 521254 71440
rect 521106 69184 521162 69193
rect 521106 69119 521162 69128
rect 521106 68368 521162 68377
rect 521106 68303 521162 68312
rect 521014 65104 521070 65113
rect 521014 65039 521070 65048
rect 521120 63753 521148 68303
rect 521212 66473 521240 71431
rect 521198 66464 521254 66473
rect 521198 66399 521254 66408
rect 521198 63880 521254 63889
rect 521198 63815 521254 63824
rect 521106 63744 521162 63753
rect 521106 63679 521162 63688
rect 520462 62384 520518 62393
rect 520462 62319 520518 62328
rect 521014 62384 521070 62393
rect 521014 62319 521070 62328
rect 520370 61024 520426 61033
rect 520370 60959 520426 60968
rect 520738 60888 520794 60897
rect 520738 60823 520794 60832
rect 116582 60616 116638 60625
rect 116582 60551 116638 60560
rect 114190 53136 114246 53145
rect 114190 53071 114246 53080
rect 116122 43344 116178 43353
rect 116122 43279 116178 43288
rect 116136 42838 116164 43279
rect 116124 42832 116176 42838
rect 116124 42774 116176 42780
rect 114098 41848 114154 41857
rect 114098 41783 114154 41792
rect 114006 30424 114062 30433
rect 114006 30359 114062 30368
rect 116490 27976 116546 27985
rect 116490 27911 116546 27920
rect 116306 26072 116362 26081
rect 116306 26007 116362 26016
rect 116214 22264 116270 22273
rect 116214 22199 116270 22208
rect 116030 20360 116086 20369
rect 116030 20295 116086 20304
rect 113914 19000 113970 19009
rect 113914 18935 113970 18944
rect 115938 16416 115994 16425
rect 115938 16351 115994 16360
rect 113822 7712 113878 7721
rect 113822 7647 113878 7656
rect 115952 2281 115980 16351
rect 116044 2553 116072 20295
rect 116122 18456 116178 18465
rect 116122 18391 116178 18400
rect 116030 2544 116086 2553
rect 116030 2479 116086 2488
rect 116136 2417 116164 18391
rect 116228 2689 116256 22199
rect 116320 3641 116348 26007
rect 116398 24168 116454 24177
rect 116398 24103 116454 24112
rect 116306 3632 116362 3641
rect 116306 3567 116362 3576
rect 116306 3088 116362 3097
rect 116306 3023 116362 3032
rect 116214 2680 116270 2689
rect 116214 2615 116270 2624
rect 116122 2408 116178 2417
rect 116122 2343 116178 2352
rect 115938 2272 115994 2281
rect 115938 2207 115994 2216
rect 116320 1290 116348 3023
rect 116308 1284 116360 1290
rect 116308 1226 116360 1232
rect 116412 1222 116440 24103
rect 116504 1426 116532 27911
rect 116596 1698 116624 60551
rect 116766 58712 116822 58721
rect 116766 58647 116822 58656
rect 116674 56808 116730 56817
rect 116674 56743 116730 56752
rect 116688 7954 116716 56743
rect 116780 7993 116808 58647
rect 519910 57896 519966 57905
rect 519910 57831 519966 57840
rect 519818 56400 519874 56409
rect 519818 56335 519874 56344
rect 519082 53408 519138 53417
rect 519082 53343 519138 53352
rect 519096 50153 519124 53343
rect 519832 52873 519860 56335
rect 519924 54233 519952 57831
rect 520752 56953 520780 60823
rect 521028 58313 521056 62319
rect 521212 59673 521240 63815
rect 521198 59664 521254 59673
rect 521198 59599 521254 59608
rect 521106 59392 521162 59401
rect 521106 59327 521162 59336
rect 521014 58304 521070 58313
rect 521014 58239 521070 58248
rect 520738 56944 520794 56953
rect 520738 56879 520794 56888
rect 521120 55593 521148 59327
rect 521106 55584 521162 55593
rect 521106 55519 521162 55528
rect 520186 54904 520242 54913
rect 520186 54839 520242 54848
rect 519910 54224 519966 54233
rect 519910 54159 519966 54168
rect 519818 52864 519874 52873
rect 519818 52799 519874 52808
rect 520094 51912 520150 51921
rect 520094 51847 520150 51856
rect 519082 50144 519138 50153
rect 519082 50079 519138 50088
rect 519082 48920 519138 48929
rect 519082 48855 519138 48864
rect 519096 46073 519124 48855
rect 520108 48793 520136 51847
rect 520200 51513 520228 54839
rect 520186 51504 520242 51513
rect 520186 51439 520242 51448
rect 520186 50416 520242 50425
rect 520186 50351 520242 50360
rect 520094 48784 520150 48793
rect 520094 48719 520150 48728
rect 520200 47433 520228 50351
rect 520186 47424 520242 47433
rect 520186 47359 520242 47368
rect 519910 47288 519966 47297
rect 519910 47223 519966 47232
rect 519082 46064 519138 46073
rect 519082 45999 519138 46008
rect 519726 45792 519782 45801
rect 519726 45727 519782 45736
rect 519740 43353 519768 45727
rect 519924 44713 519952 47223
rect 519910 44704 519966 44713
rect 519910 44639 519966 44648
rect 520186 44296 520242 44305
rect 520186 44231 520242 44240
rect 519726 43344 519782 43353
rect 519726 43279 519782 43288
rect 520200 41993 520228 44231
rect 520738 42800 520794 42809
rect 520738 42735 520794 42744
rect 520186 41984 520242 41993
rect 520186 41919 520242 41928
rect 520752 41313 520780 42735
rect 520738 41304 520794 41313
rect 520738 41239 520794 41248
rect 520922 41304 520978 41313
rect 520922 41239 520978 41248
rect 520936 39953 520964 41239
rect 520922 39944 520978 39953
rect 520922 39879 520978 39888
rect 520922 39808 520978 39817
rect 520922 39743 520978 39752
rect 116950 39536 117006 39545
rect 116950 39471 117006 39480
rect 116858 37632 116914 37641
rect 116858 37567 116914 37576
rect 116766 7984 116822 7993
rect 116676 7948 116728 7954
rect 116872 7954 116900 37567
rect 116766 7919 116822 7928
rect 116860 7948 116912 7954
rect 116676 7890 116728 7896
rect 116860 7890 116912 7896
rect 116964 7834 116992 39471
rect 520936 37913 520964 39743
rect 521106 38312 521162 38321
rect 521106 38247 521162 38256
rect 520922 37904 520978 37913
rect 520922 37839 520978 37848
rect 521120 37233 521148 38247
rect 521106 37224 521162 37233
rect 521106 37159 521162 37168
rect 521566 36816 521622 36825
rect 521566 36751 521622 36760
rect 521580 36009 521608 36751
rect 521566 36000 521622 36009
rect 521566 35935 521622 35944
rect 520922 35320 520978 35329
rect 520922 35255 520978 35264
rect 520936 34513 520964 35255
rect 520922 34504 520978 34513
rect 520922 34439 520978 34448
rect 117134 33824 117190 33833
rect 117134 33759 117190 33768
rect 521106 33824 521162 33833
rect 521106 33759 521162 33768
rect 117042 31784 117098 31793
rect 117042 31719 117098 31728
rect 116688 7806 116992 7834
rect 117056 7818 117084 31719
rect 117044 7812 117096 7818
rect 116688 3233 116716 7806
rect 117044 7754 117096 7760
rect 116860 7744 116912 7750
rect 117148 7698 117176 33759
rect 521120 33153 521148 33759
rect 521106 33144 521162 33153
rect 521106 33079 521162 33088
rect 521106 32328 521162 32337
rect 521106 32263 521162 32272
rect 521120 31657 521148 32263
rect 521106 31648 521162 31657
rect 521106 31583 521162 31592
rect 117226 29880 117282 29889
rect 117226 29815 117282 29824
rect 116860 7686 116912 7692
rect 116768 7676 116820 7682
rect 116768 7618 116820 7624
rect 116674 3224 116730 3233
rect 116674 3159 116730 3168
rect 116584 1692 116636 1698
rect 116584 1634 116636 1640
rect 116492 1420 116544 1426
rect 116492 1362 116544 1368
rect 116400 1216 116452 1222
rect 116400 1158 116452 1164
rect 116780 1154 116808 7618
rect 116768 1148 116820 1154
rect 116768 1090 116820 1096
rect 116872 1018 116900 7686
rect 116964 7670 117176 7698
rect 117240 7682 117268 29815
rect 520922 29336 520978 29345
rect 520922 29271 520978 29280
rect 520936 28393 520964 29271
rect 520922 28384 520978 28393
rect 520922 28319 520978 28328
rect 521106 24848 521162 24857
rect 521106 24783 521162 24792
rect 521120 23633 521148 24783
rect 521106 23624 521162 23633
rect 521106 23559 521162 23568
rect 520370 23216 520426 23225
rect 520370 23151 520426 23160
rect 520384 22273 520412 23151
rect 520370 22264 520426 22273
rect 520370 22199 520426 22208
rect 520922 21720 520978 21729
rect 520922 21655 520978 21664
rect 520936 20913 520964 21655
rect 520922 20904 520978 20913
rect 520922 20839 520978 20848
rect 521106 20224 521162 20233
rect 521106 20159 521162 20168
rect 521120 19553 521148 20159
rect 521106 19544 521162 19553
rect 521106 19479 521162 19488
rect 521106 9344 521162 9353
rect 521106 9279 521162 9288
rect 521120 8265 521148 9279
rect 521106 8256 521162 8265
rect 521106 8191 521162 8200
rect 520370 7984 520426 7993
rect 520370 7919 520426 7928
rect 117320 7812 117372 7818
rect 117320 7754 117372 7760
rect 117228 7676 117280 7682
rect 116964 3369 116992 7670
rect 117228 7618 117280 7624
rect 117332 7562 117360 7754
rect 117240 7534 117360 7562
rect 117044 7472 117096 7478
rect 117044 7414 117096 7420
rect 117056 5681 117084 7414
rect 117134 6896 117190 6905
rect 117134 6831 117190 6840
rect 117042 5672 117098 5681
rect 117042 5607 117098 5616
rect 116950 3360 117006 3369
rect 116950 3295 117006 3304
rect 117148 1465 117176 6831
rect 117134 1456 117190 1465
rect 117134 1391 117190 1400
rect 117240 1086 117268 7534
rect 520384 6769 520412 7919
rect 520370 6760 520426 6769
rect 520370 6695 520426 6704
rect 521106 6624 521162 6633
rect 521106 6559 521162 6568
rect 521120 5273 521148 6559
rect 520922 5264 520978 5273
rect 520922 5199 520978 5208
rect 521106 5264 521162 5273
rect 521106 5199 521162 5208
rect 520936 3777 520964 5199
rect 521014 3904 521070 3913
rect 521014 3839 521070 3848
rect 520922 3768 520978 3777
rect 520922 3703 520978 3712
rect 193600 2514 193936 2530
rect 443656 2514 443992 2530
rect 193588 2508 193936 2514
rect 193640 2502 193936 2508
rect 425796 2508 425848 2514
rect 193588 2450 193640 2456
rect 425796 2450 425848 2456
rect 443644 2508 443992 2514
rect 443696 2502 443992 2508
rect 443644 2450 443696 2456
rect 143644 2094 143980 2122
rect 243648 2094 243984 2122
rect 293604 2094 293940 2122
rect 343652 2094 343988 2122
rect 393608 2094 393944 2122
rect 143644 1494 143672 2094
rect 229282 1592 229338 1601
rect 229282 1527 229338 1536
rect 143632 1488 143684 1494
rect 143632 1430 143684 1436
rect 163778 1456 163834 1465
rect 163778 1391 163834 1400
rect 117228 1080 117280 1086
rect 117228 1022 117280 1028
rect 116860 1012 116912 1018
rect 116860 954 116912 960
rect 112536 944 112588 950
rect 112536 886 112588 892
rect 99748 876 99800 882
rect 99748 818 99800 824
rect 103888 876 103940 882
rect 103888 818 103940 824
rect 108304 876 108356 882
rect 108304 818 108356 824
rect 99564 808 99616 814
rect 95700 750 95752 756
rect 98274 -400 98330 800
rect 163792 800 163820 1391
rect 229296 800 229324 1527
rect 243648 1465 243676 2094
rect 293604 1601 293632 2094
rect 293590 1592 293646 1601
rect 293590 1527 293646 1536
rect 243634 1456 243690 1465
rect 343652 1426 343680 2094
rect 393608 1465 393636 2094
rect 360290 1456 360346 1465
rect 243634 1391 243690 1400
rect 294788 1420 294840 1426
rect 294788 1362 294840 1368
rect 343640 1420 343692 1426
rect 360290 1391 360346 1400
rect 393594 1456 393650 1465
rect 393594 1391 393650 1400
rect 343640 1362 343692 1368
rect 294800 800 294828 1362
rect 360304 800 360332 1391
rect 425808 800 425836 2450
rect 521028 2281 521056 3839
rect 521106 2680 521162 2689
rect 521106 2615 521162 2624
rect 521014 2272 521070 2281
rect 521014 2207 521070 2216
rect 493612 2094 493948 2122
rect 493612 1426 493640 2094
rect 491300 1420 491352 1426
rect 491300 1362 491352 1368
rect 493600 1420 493652 1426
rect 493600 1362 493652 1368
rect 491312 800 491340 1362
rect 99564 750 99616 756
rect 163778 -400 163834 800
rect 229282 -400 229338 800
rect 294786 -400 294842 800
rect 360290 -400 360346 800
rect 425794 -400 425850 800
rect 491298 -400 491354 800
rect 521120 785 521148 2615
rect 521106 776 521162 785
rect 521106 711 521162 720
<< via2 >>
rect 2962 153720 3018 153776
rect 16302 159296 16358 159352
rect 16578 153856 16634 153912
rect 19890 153992 19946 154048
rect 23018 159432 23074 159488
rect 12438 152496 12494 152552
rect 8850 152360 8906 152416
rect 6090 150592 6146 150648
rect 2686 150456 2742 150512
rect 28078 156576 28134 156632
rect 29826 159568 29882 159624
rect 31482 156712 31538 156768
rect 30378 154128 30434 154184
rect 33966 157936 34022 157992
rect 40682 158208 40738 158264
rect 44086 158072 44142 158128
rect 57518 158344 57574 158400
rect 55862 156848 55918 156904
rect 54298 154264 54354 154320
rect 62578 155488 62634 155544
rect 65982 155216 66038 155272
rect 72698 156984 72754 157040
rect 68466 155352 68522 155408
rect 76010 155760 76066 155816
rect 78586 155624 78642 155680
rect 85302 155896 85358 155952
rect 85578 154400 85634 154456
rect 104622 158480 104678 158536
rect 82818 149640 82874 149696
rect 109590 148008 109646 148064
rect 115570 157120 115626 157176
rect 110878 150456 110934 150512
rect 111246 150592 111302 150648
rect 110326 146376 110382 146432
rect 110326 106256 110382 106312
rect 113822 144200 113878 144256
rect 116122 145152 116178 145208
rect 116030 143248 116086 143304
rect 115294 141344 115350 141400
rect 116122 139440 116178 139496
rect 116122 137536 116178 137592
rect 115202 135496 115258 135552
rect 116030 133592 116086 133648
rect 114190 132776 114246 132832
rect 113914 121352 113970 121408
rect 114006 110064 114062 110120
rect 114098 98640 114154 98696
rect 114190 87216 114246 87272
rect 116122 131688 116178 131744
rect 116582 149640 116638 149696
rect 116490 129784 116546 129840
rect 116122 125976 116178 126032
rect 116122 124108 116124 124128
rect 116124 124108 116176 124128
rect 116176 124108 116178 124128
rect 116122 124072 116178 124108
rect 115938 122168 115994 122224
rect 116122 120128 116178 120184
rect 116122 118224 116178 118280
rect 116122 116320 116178 116376
rect 116122 114452 116124 114472
rect 116124 114452 116176 114472
rect 116176 114452 116178 114472
rect 116122 114416 116178 114452
rect 115938 112512 115994 112568
rect 116122 110608 116178 110664
rect 116122 108704 116178 108760
rect 116950 102856 117006 102912
rect 121734 153720 121790 153776
rect 121918 153720 121974 153776
rect 126242 152360 126298 152416
rect 126794 152360 126850 152416
rect 131026 159296 131082 159352
rect 128818 152496 128874 152552
rect 133602 159432 133658 159488
rect 132038 153856 132094 153912
rect 133602 153040 133658 153096
rect 134614 153992 134670 154048
rect 136546 153040 136602 153096
rect 138018 159568 138074 159624
rect 140410 156576 140466 156632
rect 143078 156712 143134 156768
rect 142250 153992 142306 154048
rect 142434 154028 142436 154048
rect 142436 154028 142488 154048
rect 142488 154028 142490 154048
rect 142434 153992 142490 154028
rect 142986 153992 143042 154048
rect 145102 157936 145158 157992
rect 143630 152360 143686 152416
rect 147586 154164 147588 154184
rect 147588 154164 147640 154184
rect 147640 154164 147642 154184
rect 147586 154128 147642 154164
rect 148138 154128 148194 154184
rect 149610 158208 149666 158264
rect 152554 158072 152610 158128
rect 161662 156848 161718 156904
rect 160926 154264 160982 154320
rect 162858 158344 162914 158400
rect 166722 155488 166778 155544
rect 168378 155216 168434 155272
rect 171230 155352 171286 155408
rect 174450 156984 174506 157040
rect 177026 155760 177082 155816
rect 178958 155624 179014 155680
rect 184018 155896 184074 155952
rect 184662 154400 184718 154456
rect 190918 154436 190920 154456
rect 190920 154436 190972 154456
rect 190972 154436 190974 154456
rect 190918 154400 190974 154436
rect 191286 154400 191342 154456
rect 192390 153720 192446 153776
rect 195886 153448 195942 153504
rect 196070 153448 196126 153504
rect 198738 158480 198794 158536
rect 204718 159296 204774 159352
rect 207202 157120 207258 157176
rect 211526 153720 211582 153776
rect 227442 152360 227498 152416
rect 274546 159432 274602 159488
rect 275190 159296 275246 159352
rect 280986 153720 281042 153776
rect 292578 152360 292634 152416
rect 313370 152360 313426 152416
rect 328550 159432 328606 159488
rect 357438 152360 357494 152416
rect 407670 152360 407726 152416
rect 421930 152516 421986 152552
rect 421930 152496 421932 152516
rect 421932 152496 421984 152516
rect 421984 152496 421986 152516
rect 424506 152496 424562 152552
rect 430578 152360 430634 152416
rect 431222 152496 431278 152552
rect 443918 153076 443920 153096
rect 443920 153076 443972 153096
rect 443972 153076 443974 153096
rect 443918 153040 443974 153076
rect 444930 153040 444986 153096
rect 448610 152496 448666 152552
rect 519726 163104 519782 163160
rect 519542 161608 519598 161664
rect 519450 151136 519506 151192
rect 519358 140528 519414 140584
rect 519634 160112 519690 160168
rect 519542 147872 519598 147928
rect 519818 157120 519874 157176
rect 519726 149232 519782 149288
rect 519726 148144 519782 148200
rect 519634 146512 519690 146568
rect 519634 145152 519690 145208
rect 519542 142160 519598 142216
rect 519450 138352 519506 138408
rect 519450 136040 519506 136096
rect 519358 128832 519414 128888
rect 117226 127880 117282 127936
rect 520186 158616 520242 158672
rect 520094 155624 520150 155680
rect 520002 154128 520058 154184
rect 519910 149640 519966 149696
rect 519818 143792 519874 143848
rect 521014 152632 521070 152688
rect 520186 145288 520242 145344
rect 520922 143656 520978 143712
rect 520094 142432 520150 142488
rect 520002 141072 520058 141128
rect 520002 139032 520058 139088
rect 519910 136992 519966 137048
rect 519726 135632 519782 135688
rect 519818 133048 519874 133104
rect 519634 132912 519690 132968
rect 519542 130192 519598 130248
rect 519726 130056 519782 130112
rect 519634 128560 519690 128616
rect 519542 127064 519598 127120
rect 519450 124752 519506 124808
rect 519266 124072 519322 124128
rect 519358 122576 519414 122632
rect 519266 113872 519322 113928
rect 519450 119584 519506 119640
rect 519358 112512 519414 112568
rect 519910 131552 519966 131608
rect 519818 122032 519874 122088
rect 520186 137536 520242 137592
rect 520094 134544 520150 134600
rect 520002 127472 520058 127528
rect 520002 125568 520058 125624
rect 519910 120672 519966 120728
rect 519726 119312 519782 119368
rect 519818 118088 519874 118144
rect 519634 117952 519690 118008
rect 519542 116592 519598 116648
rect 519726 113464 519782 113520
rect 519634 111968 519690 112024
rect 519542 110472 519598 110528
rect 519450 109792 519506 109848
rect 117134 104760 117190 104816
rect 519910 116456 519966 116512
rect 519818 108432 519874 108488
rect 521106 146648 521162 146704
rect 521014 139712 521070 139768
rect 521106 134272 521162 134328
rect 520922 131688 520978 131744
rect 520186 126112 520242 126168
rect 520094 123392 520150 123448
rect 520094 121080 520150 121136
rect 520002 115232 520058 115288
rect 520186 114960 520242 115016
rect 520094 111152 520150 111208
rect 519910 107072 519966 107128
rect 521290 108976 521346 109032
rect 521106 107480 521162 107536
rect 520278 105984 520334 106040
rect 520186 105712 520242 105768
rect 519726 104352 519782 104408
rect 519634 102992 519690 103048
rect 519542 101632 519598 101688
rect 117042 100952 117098 101008
rect 116858 99048 116914 99104
rect 521014 104488 521070 104544
rect 520922 101496 520978 101552
rect 520278 97552 520334 97608
rect 116766 97144 116822 97200
rect 520278 95512 520334 95568
rect 116674 95240 116730 95296
rect 116582 93336 116638 93392
rect 519634 92384 519690 92440
rect 116122 91296 116178 91352
rect 116122 89392 116178 89448
rect 116030 87488 116086 87544
rect 115202 85584 115258 85640
rect 520002 90888 520058 90944
rect 519726 89392 519782 89448
rect 519634 85312 519690 85368
rect 519082 84904 519138 84960
rect 116582 83680 116638 83736
rect 116214 81776 116270 81832
rect 115938 79872 115994 79928
rect 519910 87896 519966 87952
rect 519818 86400 519874 86456
rect 519726 82592 519782 82648
rect 519450 81912 519506 81968
rect 519082 78512 519138 78568
rect 116122 77968 116178 78024
rect 521198 102992 521254 103048
rect 521106 98912 521162 98968
rect 521014 96192 521070 96248
rect 521290 100272 521346 100328
rect 521474 100000 521530 100056
rect 521290 98504 521346 98560
rect 521198 94832 521254 94888
rect 521014 93880 521070 93936
rect 520922 93472 520978 93528
rect 520278 88032 520334 88088
rect 521382 97008 521438 97064
rect 521290 90752 521346 90808
rect 521474 92112 521530 92168
rect 521382 89528 521438 89584
rect 521014 86672 521070 86728
rect 520002 83952 520058 84008
rect 520094 83408 520150 83464
rect 519910 81232 519966 81288
rect 519818 79872 519874 79928
rect 520002 78920 520058 78976
rect 519818 77424 519874 77480
rect 519450 75928 519506 75984
rect 116674 74024 116730 74080
rect 116582 72120 116638 72176
rect 113362 64504 113418 64560
rect 110326 53896 110382 53952
rect 110326 52536 110382 52592
rect 110326 51040 110382 51096
rect 109498 3848 109554 3904
rect 109498 3440 109554 3496
rect 32402 2624 32458 2680
rect 36358 2624 36414 2680
rect 62394 2624 62450 2680
rect 64142 2624 64198 2680
rect 65338 2624 65394 2680
rect 68006 2624 68062 2680
rect 68282 2624 68338 2680
rect 68466 2624 68522 2680
rect 69386 2624 69442 2680
rect 75642 2624 75698 2680
rect 29550 2352 29606 2408
rect 26054 2216 26110 2272
rect 5998 1672 6054 1728
rect 22926 2080 22982 2136
rect 19614 1944 19670 2000
rect 15934 1808 15990 1864
rect 12622 1536 12678 1592
rect 9310 1400 9366 1456
rect 33046 2488 33102 2544
rect 77482 2624 77538 2680
rect 85394 2624 85450 2680
rect 86682 2624 86738 2680
rect 91742 2624 91798 2680
rect 93030 2624 93086 2680
rect 98918 2624 98974 2680
rect 99194 2624 99250 2680
rect 99562 2624 99618 2680
rect 99746 2624 99802 2680
rect 91650 2488 91706 2544
rect 87970 2080 88026 2136
rect 91650 2080 91706 2136
rect 86682 1264 86738 1320
rect 89258 1128 89314 1184
rect 95698 2488 95754 2544
rect 96342 2488 96398 2544
rect 98274 1128 98330 1184
rect 99838 2488 99894 2544
rect 103426 2624 103482 2680
rect 104162 2488 104218 2544
rect 104162 2080 104218 2136
rect 104346 2080 104402 2136
rect 103334 1264 103390 1320
rect 99838 992 99894 1048
rect 108210 1264 108266 1320
rect 109866 3576 109922 3632
rect 109866 2760 109922 2816
rect 109498 1672 109554 1728
rect 110326 48320 110382 48376
rect 110326 47096 110382 47152
rect 110326 44240 110382 44296
rect 110326 41384 110382 41440
rect 110326 34584 110382 34640
rect 110326 8200 110382 8256
rect 110510 8200 110566 8256
rect 110234 3848 110290 3904
rect 110234 3440 110290 3496
rect 110142 2896 110198 2952
rect 110602 5616 110658 5672
rect 111062 7928 111118 7984
rect 110694 3168 110750 3224
rect 110602 2760 110658 2816
rect 111706 2896 111762 2952
rect 110234 1264 110290 1320
rect 110142 1128 110198 1184
rect 116306 70216 116362 70272
rect 116122 68312 116178 68368
rect 116582 66408 116638 66464
rect 519910 75928 519966 75984
rect 519818 71848 519874 71904
rect 520186 80416 520242 80472
rect 520094 77152 520150 77208
rect 520186 74568 520242 74624
rect 521106 74432 521162 74488
rect 520002 73208 520058 73264
rect 520922 72936 520978 72992
rect 519910 70488 519966 70544
rect 521014 69808 521070 69864
rect 520922 67768 520978 67824
rect 520462 66816 520518 66872
rect 520370 65320 520426 65376
rect 116214 64504 116270 64560
rect 116122 62600 116178 62656
rect 521198 71440 521254 71496
rect 521106 69128 521162 69184
rect 521106 68312 521162 68368
rect 521014 65048 521070 65104
rect 521198 66408 521254 66464
rect 521198 63824 521254 63880
rect 521106 63688 521162 63744
rect 520462 62328 520518 62384
rect 521014 62328 521070 62384
rect 520370 60968 520426 61024
rect 520738 60832 520794 60888
rect 116582 60560 116638 60616
rect 114190 53080 114246 53136
rect 116122 43288 116178 43344
rect 114098 41792 114154 41848
rect 114006 30368 114062 30424
rect 116490 27920 116546 27976
rect 116306 26016 116362 26072
rect 116214 22208 116270 22264
rect 116030 20304 116086 20360
rect 113914 18944 113970 19000
rect 115938 16360 115994 16416
rect 113822 7656 113878 7712
rect 116122 18400 116178 18456
rect 116030 2488 116086 2544
rect 116398 24112 116454 24168
rect 116306 3576 116362 3632
rect 116306 3032 116362 3088
rect 116214 2624 116270 2680
rect 116122 2352 116178 2408
rect 115938 2216 115994 2272
rect 116766 58656 116822 58712
rect 116674 56752 116730 56808
rect 519910 57840 519966 57896
rect 519818 56344 519874 56400
rect 519082 53352 519138 53408
rect 521198 59608 521254 59664
rect 521106 59336 521162 59392
rect 521014 58248 521070 58304
rect 520738 56888 520794 56944
rect 521106 55528 521162 55584
rect 520186 54848 520242 54904
rect 519910 54168 519966 54224
rect 519818 52808 519874 52864
rect 520094 51856 520150 51912
rect 519082 50088 519138 50144
rect 519082 48864 519138 48920
rect 520186 51448 520242 51504
rect 520186 50360 520242 50416
rect 520094 48728 520150 48784
rect 520186 47368 520242 47424
rect 519910 47232 519966 47288
rect 519082 46008 519138 46064
rect 519726 45736 519782 45792
rect 519910 44648 519966 44704
rect 520186 44240 520242 44296
rect 519726 43288 519782 43344
rect 520738 42744 520794 42800
rect 520186 41928 520242 41984
rect 520738 41248 520794 41304
rect 520922 41248 520978 41304
rect 520922 39888 520978 39944
rect 520922 39752 520978 39808
rect 116950 39480 117006 39536
rect 116858 37576 116914 37632
rect 116766 7928 116822 7984
rect 521106 38256 521162 38312
rect 520922 37848 520978 37904
rect 521106 37168 521162 37224
rect 521566 36760 521622 36816
rect 521566 35944 521622 36000
rect 520922 35264 520978 35320
rect 520922 34448 520978 34504
rect 117134 33768 117190 33824
rect 521106 33768 521162 33824
rect 117042 31728 117098 31784
rect 521106 33088 521162 33144
rect 521106 32272 521162 32328
rect 521106 31592 521162 31648
rect 117226 29824 117282 29880
rect 116674 3168 116730 3224
rect 520922 29280 520978 29336
rect 520922 28328 520978 28384
rect 521106 24792 521162 24848
rect 521106 23568 521162 23624
rect 520370 23160 520426 23216
rect 520370 22208 520426 22264
rect 520922 21664 520978 21720
rect 520922 20848 520978 20904
rect 521106 20168 521162 20224
rect 521106 19488 521162 19544
rect 521106 9288 521162 9344
rect 521106 8200 521162 8256
rect 520370 7928 520426 7984
rect 117134 6840 117190 6896
rect 117042 5616 117098 5672
rect 116950 3304 117006 3360
rect 117134 1400 117190 1456
rect 520370 6704 520426 6760
rect 521106 6568 521162 6624
rect 520922 5208 520978 5264
rect 521106 5208 521162 5264
rect 521014 3848 521070 3904
rect 520922 3712 520978 3768
rect 229282 1536 229338 1592
rect 163778 1400 163834 1456
rect 293590 1536 293646 1592
rect 243634 1400 243690 1456
rect 360290 1400 360346 1456
rect 393594 1400 393650 1456
rect 521106 2624 521162 2680
rect 521014 2216 521070 2272
rect 521106 720 521162 776
<< metal3 >>
rect 519721 163162 519787 163165
rect 523200 163162 524400 163192
rect 519721 163160 524400 163162
rect 519721 163104 519726 163160
rect 519782 163104 524400 163160
rect 519721 163102 524400 163104
rect 519721 163099 519787 163102
rect 523200 163072 524400 163102
rect 519537 161666 519603 161669
rect 523200 161666 524400 161696
rect 519537 161664 524400 161666
rect 519537 161608 519542 161664
rect 519598 161608 524400 161664
rect 519537 161606 524400 161608
rect 519537 161603 519603 161606
rect 523200 161576 524400 161606
rect 519629 160170 519695 160173
rect 523200 160170 524400 160200
rect 519629 160168 524400 160170
rect 519629 160112 519634 160168
rect 519690 160112 524400 160168
rect 519629 160110 524400 160112
rect 519629 160107 519695 160110
rect 523200 160080 524400 160110
rect 29821 159626 29887 159629
rect 138013 159626 138079 159629
rect 29821 159624 138079 159626
rect 29821 159568 29826 159624
rect 29882 159568 138018 159624
rect 138074 159568 138079 159624
rect 29821 159566 138079 159568
rect 29821 159563 29887 159566
rect 138013 159563 138079 159566
rect 23013 159490 23079 159493
rect 133597 159490 133663 159493
rect 23013 159488 133663 159490
rect 23013 159432 23018 159488
rect 23074 159432 133602 159488
rect 133658 159432 133663 159488
rect 23013 159430 133663 159432
rect 23013 159427 23079 159430
rect 133597 159427 133663 159430
rect 274541 159490 274607 159493
rect 328545 159490 328611 159493
rect 274541 159488 328611 159490
rect 274541 159432 274546 159488
rect 274602 159432 328550 159488
rect 328606 159432 328611 159488
rect 274541 159430 328611 159432
rect 274541 159427 274607 159430
rect 328545 159427 328611 159430
rect 16297 159354 16363 159357
rect 131021 159354 131087 159357
rect 16297 159352 131087 159354
rect 16297 159296 16302 159352
rect 16358 159296 131026 159352
rect 131082 159296 131087 159352
rect 16297 159294 131087 159296
rect 16297 159291 16363 159294
rect 131021 159291 131087 159294
rect 204713 159354 204779 159357
rect 275185 159354 275251 159357
rect 204713 159352 275251 159354
rect 204713 159296 204718 159352
rect 204774 159296 275190 159352
rect 275246 159296 275251 159352
rect 204713 159294 275251 159296
rect 204713 159291 204779 159294
rect 275185 159291 275251 159294
rect 520181 158674 520247 158677
rect 523200 158674 524400 158704
rect 520181 158672 524400 158674
rect 520181 158616 520186 158672
rect 520242 158616 524400 158672
rect 520181 158614 524400 158616
rect 520181 158611 520247 158614
rect 523200 158584 524400 158614
rect 104617 158538 104683 158541
rect 198733 158538 198799 158541
rect 104617 158536 198799 158538
rect 104617 158480 104622 158536
rect 104678 158480 198738 158536
rect 198794 158480 198799 158536
rect 104617 158478 198799 158480
rect 104617 158475 104683 158478
rect 198733 158475 198799 158478
rect 57513 158402 57579 158405
rect 162853 158402 162919 158405
rect 57513 158400 162919 158402
rect 57513 158344 57518 158400
rect 57574 158344 162858 158400
rect 162914 158344 162919 158400
rect 57513 158342 162919 158344
rect 57513 158339 57579 158342
rect 162853 158339 162919 158342
rect 40677 158266 40743 158269
rect 149605 158266 149671 158269
rect 40677 158264 149671 158266
rect 40677 158208 40682 158264
rect 40738 158208 149610 158264
rect 149666 158208 149671 158264
rect 40677 158206 149671 158208
rect 40677 158203 40743 158206
rect 149605 158203 149671 158206
rect 44081 158130 44147 158133
rect 152549 158130 152615 158133
rect 44081 158128 152615 158130
rect 44081 158072 44086 158128
rect 44142 158072 152554 158128
rect 152610 158072 152615 158128
rect 44081 158070 152615 158072
rect 44081 158067 44147 158070
rect 152549 158067 152615 158070
rect 33961 157994 34027 157997
rect 145097 157994 145163 157997
rect 33961 157992 145163 157994
rect 33961 157936 33966 157992
rect 34022 157936 145102 157992
rect 145158 157936 145163 157992
rect 33961 157934 145163 157936
rect 33961 157931 34027 157934
rect 145097 157931 145163 157934
rect 115565 157178 115631 157181
rect 207197 157178 207263 157181
rect 115565 157176 207263 157178
rect 115565 157120 115570 157176
rect 115626 157120 207202 157176
rect 207258 157120 207263 157176
rect 115565 157118 207263 157120
rect 115565 157115 115631 157118
rect 207197 157115 207263 157118
rect 519813 157178 519879 157181
rect 523200 157178 524400 157208
rect 519813 157176 524400 157178
rect 519813 157120 519818 157176
rect 519874 157120 524400 157176
rect 519813 157118 524400 157120
rect 519813 157115 519879 157118
rect 523200 157088 524400 157118
rect 72693 157042 72759 157045
rect 174445 157042 174511 157045
rect 72693 157040 174511 157042
rect 72693 156984 72698 157040
rect 72754 156984 174450 157040
rect 174506 156984 174511 157040
rect 72693 156982 174511 156984
rect 72693 156979 72759 156982
rect 174445 156979 174511 156982
rect 55857 156906 55923 156909
rect 161657 156906 161723 156909
rect 55857 156904 161723 156906
rect 55857 156848 55862 156904
rect 55918 156848 161662 156904
rect 161718 156848 161723 156904
rect 55857 156846 161723 156848
rect 55857 156843 55923 156846
rect 161657 156843 161723 156846
rect 31477 156770 31543 156773
rect 143073 156770 143139 156773
rect 31477 156768 143139 156770
rect 31477 156712 31482 156768
rect 31538 156712 143078 156768
rect 143134 156712 143139 156768
rect 31477 156710 143139 156712
rect 31477 156707 31543 156710
rect 143073 156707 143139 156710
rect 28073 156634 28139 156637
rect 140405 156634 140471 156637
rect 28073 156632 140471 156634
rect 28073 156576 28078 156632
rect 28134 156576 140410 156632
rect 140466 156576 140471 156632
rect 28073 156574 140471 156576
rect 28073 156571 28139 156574
rect 140405 156571 140471 156574
rect 85297 155954 85363 155957
rect 184013 155954 184079 155957
rect 85297 155952 184079 155954
rect 85297 155896 85302 155952
rect 85358 155896 184018 155952
rect 184074 155896 184079 155952
rect 85297 155894 184079 155896
rect 85297 155891 85363 155894
rect 184013 155891 184079 155894
rect 76005 155818 76071 155821
rect 177021 155818 177087 155821
rect 76005 155816 177087 155818
rect 76005 155760 76010 155816
rect 76066 155760 177026 155816
rect 177082 155760 177087 155816
rect 76005 155758 177087 155760
rect 76005 155755 76071 155758
rect 177021 155755 177087 155758
rect 78581 155682 78647 155685
rect 178953 155682 179019 155685
rect 78581 155680 179019 155682
rect 78581 155624 78586 155680
rect 78642 155624 178958 155680
rect 179014 155624 179019 155680
rect 78581 155622 179019 155624
rect 78581 155619 78647 155622
rect 178953 155619 179019 155622
rect 520089 155682 520155 155685
rect 523200 155682 524400 155712
rect 520089 155680 524400 155682
rect 520089 155624 520094 155680
rect 520150 155624 524400 155680
rect 520089 155622 524400 155624
rect 520089 155619 520155 155622
rect 523200 155592 524400 155622
rect 62573 155546 62639 155549
rect 166717 155546 166783 155549
rect 62573 155544 166783 155546
rect 62573 155488 62578 155544
rect 62634 155488 166722 155544
rect 166778 155488 166783 155544
rect 62573 155486 166783 155488
rect 62573 155483 62639 155486
rect 166717 155483 166783 155486
rect 68461 155410 68527 155413
rect 171225 155410 171291 155413
rect 68461 155408 171291 155410
rect 68461 155352 68466 155408
rect 68522 155352 171230 155408
rect 171286 155352 171291 155408
rect 68461 155350 171291 155352
rect 68461 155347 68527 155350
rect 171225 155347 171291 155350
rect 65977 155274 66043 155277
rect 168373 155274 168439 155277
rect 65977 155272 168439 155274
rect 65977 155216 65982 155272
rect 66038 155216 168378 155272
rect 168434 155216 168439 155272
rect 65977 155214 168439 155216
rect 65977 155211 66043 155214
rect 168373 155211 168439 155214
rect 85573 154458 85639 154461
rect 184657 154458 184723 154461
rect 85573 154456 184723 154458
rect 85573 154400 85578 154456
rect 85634 154400 184662 154456
rect 184718 154400 184723 154456
rect 85573 154398 184723 154400
rect 85573 154395 85639 154398
rect 184657 154395 184723 154398
rect 190913 154458 190979 154461
rect 191281 154458 191347 154461
rect 190913 154456 191347 154458
rect 190913 154400 190918 154456
rect 190974 154400 191286 154456
rect 191342 154400 191347 154456
rect 190913 154398 191347 154400
rect 190913 154395 190979 154398
rect 191281 154395 191347 154398
rect 54293 154322 54359 154325
rect 160921 154322 160987 154325
rect 54293 154320 160987 154322
rect 54293 154264 54298 154320
rect 54354 154264 160926 154320
rect 160982 154264 160987 154320
rect 54293 154262 160987 154264
rect 54293 154259 54359 154262
rect 160921 154259 160987 154262
rect 30373 154186 30439 154189
rect 147581 154186 147647 154189
rect 148133 154186 148199 154189
rect 30373 154184 138030 154186
rect 30373 154128 30378 154184
rect 30434 154128 138030 154184
rect 30373 154126 138030 154128
rect 30373 154123 30439 154126
rect 19885 154050 19951 154053
rect 134609 154050 134675 154053
rect 19885 154048 134675 154050
rect 19885 153992 19890 154048
rect 19946 153992 134614 154048
rect 134670 153992 134675 154048
rect 19885 153990 134675 153992
rect 137970 154050 138030 154126
rect 147581 154184 148199 154186
rect 147581 154128 147586 154184
rect 147642 154128 148138 154184
rect 148194 154128 148199 154184
rect 147581 154126 148199 154128
rect 147581 154123 147647 154126
rect 148133 154123 148199 154126
rect 519997 154186 520063 154189
rect 523200 154186 524400 154216
rect 519997 154184 524400 154186
rect 519997 154128 520002 154184
rect 520058 154128 524400 154184
rect 519997 154126 524400 154128
rect 519997 154123 520063 154126
rect 523200 154096 524400 154126
rect 142245 154050 142311 154053
rect 137970 154048 142311 154050
rect 137970 153992 142250 154048
rect 142306 153992 142311 154048
rect 137970 153990 142311 153992
rect 19885 153987 19951 153990
rect 134609 153987 134675 153990
rect 142245 153987 142311 153990
rect 142429 154050 142495 154053
rect 142981 154050 143047 154053
rect 142429 154048 143047 154050
rect 142429 153992 142434 154048
rect 142490 153992 142986 154048
rect 143042 153992 143047 154048
rect 142429 153990 143047 153992
rect 142429 153987 142495 153990
rect 142981 153987 143047 153990
rect 16573 153914 16639 153917
rect 132033 153914 132099 153917
rect 16573 153912 132099 153914
rect 16573 153856 16578 153912
rect 16634 153856 132038 153912
rect 132094 153856 132099 153912
rect 16573 153854 132099 153856
rect 16573 153851 16639 153854
rect 132033 153851 132099 153854
rect 2957 153778 3023 153781
rect 121729 153778 121795 153781
rect 2957 153776 121795 153778
rect 2957 153720 2962 153776
rect 3018 153720 121734 153776
rect 121790 153720 121795 153776
rect 2957 153718 121795 153720
rect 2957 153715 3023 153718
rect 121729 153715 121795 153718
rect 121913 153778 121979 153781
rect 192385 153778 192451 153781
rect 121913 153776 192451 153778
rect 121913 153720 121918 153776
rect 121974 153720 192390 153776
rect 192446 153720 192451 153776
rect 121913 153718 192451 153720
rect 121913 153715 121979 153718
rect 192385 153715 192451 153718
rect 211521 153778 211587 153781
rect 280981 153778 281047 153781
rect 211521 153776 281047 153778
rect 211521 153720 211526 153776
rect 211582 153720 280986 153776
rect 281042 153720 281047 153776
rect 211521 153718 281047 153720
rect 211521 153715 211587 153718
rect 280981 153715 281047 153718
rect 195881 153506 195947 153509
rect 196065 153506 196131 153509
rect 195881 153504 196131 153506
rect 195881 153448 195886 153504
rect 195942 153448 196070 153504
rect 196126 153448 196131 153504
rect 195881 153446 196131 153448
rect 195881 153443 195947 153446
rect 196065 153443 196131 153446
rect 133597 153098 133663 153101
rect 136541 153098 136607 153101
rect 133597 153096 136607 153098
rect 133597 153040 133602 153096
rect 133658 153040 136546 153096
rect 136602 153040 136607 153096
rect 133597 153038 136607 153040
rect 133597 153035 133663 153038
rect 136541 153035 136607 153038
rect 443913 153098 443979 153101
rect 444925 153098 444991 153101
rect 443913 153096 444991 153098
rect 443913 153040 443918 153096
rect 443974 153040 444930 153096
rect 444986 153040 444991 153096
rect 443913 153038 444991 153040
rect 443913 153035 443979 153038
rect 444925 153035 444991 153038
rect 521009 152690 521075 152693
rect 523200 152690 524400 152720
rect 521009 152688 524400 152690
rect 521009 152632 521014 152688
rect 521070 152632 524400 152688
rect 521009 152630 524400 152632
rect 521009 152627 521075 152630
rect 523200 152600 524400 152630
rect 12433 152554 12499 152557
rect 128813 152554 128879 152557
rect 12433 152552 128879 152554
rect 12433 152496 12438 152552
rect 12494 152496 128818 152552
rect 128874 152496 128879 152552
rect 12433 152494 128879 152496
rect 12433 152491 12499 152494
rect 128813 152491 128879 152494
rect 421925 152554 421991 152557
rect 424501 152554 424567 152557
rect 421925 152552 424567 152554
rect 421925 152496 421930 152552
rect 421986 152496 424506 152552
rect 424562 152496 424567 152552
rect 421925 152494 424567 152496
rect 421925 152491 421991 152494
rect 424501 152491 424567 152494
rect 431217 152554 431283 152557
rect 448605 152554 448671 152557
rect 431217 152552 448671 152554
rect 431217 152496 431222 152552
rect 431278 152496 448610 152552
rect 448666 152496 448671 152552
rect 431217 152494 448671 152496
rect 431217 152491 431283 152494
rect 448605 152491 448671 152494
rect 8845 152418 8911 152421
rect 126237 152418 126303 152421
rect 8845 152416 126303 152418
rect 8845 152360 8850 152416
rect 8906 152360 126242 152416
rect 126298 152360 126303 152416
rect 8845 152358 126303 152360
rect 8845 152355 8911 152358
rect 126237 152355 126303 152358
rect 126789 152418 126855 152421
rect 143625 152418 143691 152421
rect 126789 152416 143691 152418
rect 126789 152360 126794 152416
rect 126850 152360 143630 152416
rect 143686 152360 143691 152416
rect 126789 152358 143691 152360
rect 126789 152355 126855 152358
rect 143625 152355 143691 152358
rect 227437 152418 227503 152421
rect 292573 152418 292639 152421
rect 227437 152416 292639 152418
rect 227437 152360 227442 152416
rect 227498 152360 292578 152416
rect 292634 152360 292639 152416
rect 227437 152358 292639 152360
rect 227437 152355 227503 152358
rect 292573 152355 292639 152358
rect 313365 152418 313431 152421
rect 357433 152418 357499 152421
rect 313365 152416 357499 152418
rect 313365 152360 313370 152416
rect 313426 152360 357438 152416
rect 357494 152360 357499 152416
rect 313365 152358 357499 152360
rect 313365 152355 313431 152358
rect 357433 152355 357499 152358
rect 407665 152418 407731 152421
rect 430573 152418 430639 152421
rect 407665 152416 430639 152418
rect 407665 152360 407670 152416
rect 407726 152360 430578 152416
rect 430634 152360 430639 152416
rect 407665 152358 430639 152360
rect 407665 152355 407731 152358
rect 430573 152355 430639 152358
rect 519445 151194 519511 151197
rect 523200 151194 524400 151224
rect 519445 151192 524400 151194
rect 519445 151136 519450 151192
rect 519506 151136 524400 151192
rect 519445 151134 524400 151136
rect 519445 151131 519511 151134
rect 523200 151104 524400 151134
rect 6085 150650 6151 150653
rect 111241 150650 111307 150653
rect 6085 150648 111307 150650
rect 6085 150592 6090 150648
rect 6146 150592 111246 150648
rect 111302 150592 111307 150648
rect 6085 150590 111307 150592
rect 6085 150587 6151 150590
rect 111241 150587 111307 150590
rect 2681 150514 2747 150517
rect 110873 150514 110939 150517
rect 2681 150512 110939 150514
rect 2681 150456 2686 150512
rect 2742 150456 110878 150512
rect 110934 150456 110939 150512
rect 2681 150454 110939 150456
rect 2681 150451 2747 150454
rect 110873 150451 110939 150454
rect 82813 149698 82879 149701
rect 116577 149698 116643 149701
rect 82813 149696 116643 149698
rect 82813 149640 82818 149696
rect 82874 149640 116582 149696
rect 116638 149640 116643 149696
rect 82813 149638 116643 149640
rect 82813 149635 82879 149638
rect 116577 149635 116643 149638
rect 519905 149698 519971 149701
rect 523200 149698 524400 149728
rect 519905 149696 524400 149698
rect 519905 149640 519910 149696
rect 519966 149640 524400 149696
rect 519905 149638 524400 149640
rect 519905 149635 519971 149638
rect 523200 149608 524400 149638
rect 519721 149290 519787 149293
rect 518788 149288 519787 149290
rect 518788 149232 519726 149288
rect 519782 149232 519787 149288
rect 518788 149230 519787 149232
rect 519721 149227 519787 149230
rect 109585 148066 109651 148069
rect 119110 148066 119170 148988
rect 519721 148202 519787 148205
rect 523200 148202 524400 148232
rect 519721 148200 524400 148202
rect 519721 148144 519726 148200
rect 519782 148144 524400 148200
rect 519721 148142 524400 148144
rect 519721 148139 519787 148142
rect 523200 148112 524400 148142
rect 109585 148064 119170 148066
rect 109585 148008 109590 148064
rect 109646 148008 119170 148064
rect 109585 148006 119170 148008
rect 109585 148003 109651 148006
rect 519537 147930 519603 147933
rect 518788 147928 519603 147930
rect 518788 147872 519542 147928
rect 519598 147872 519603 147928
rect 518788 147870 519603 147872
rect 519537 147867 519603 147870
rect 110321 146434 110387 146437
rect 119110 146434 119170 147084
rect 521101 146706 521167 146709
rect 523200 146706 524400 146736
rect 521101 146704 524400 146706
rect 521101 146648 521106 146704
rect 521162 146648 524400 146704
rect 521101 146646 524400 146648
rect 521101 146643 521167 146646
rect 523200 146616 524400 146646
rect 519629 146570 519695 146573
rect 518788 146568 519695 146570
rect 518788 146512 519634 146568
rect 519690 146512 519695 146568
rect 518788 146510 519695 146512
rect 519629 146507 519695 146510
rect 110321 146432 119170 146434
rect 110321 146376 110326 146432
rect 110382 146376 119170 146432
rect 110321 146374 119170 146376
rect 110321 146371 110387 146374
rect 520181 145346 520247 145349
rect 518758 145344 520247 145346
rect 518758 145288 520186 145344
rect 520242 145288 520247 145344
rect 518758 145286 520247 145288
rect 116117 145210 116183 145213
rect 116117 145208 119140 145210
rect 116117 145152 116122 145208
rect 116178 145152 119140 145208
rect 518758 145180 518818 145286
rect 520181 145283 520247 145286
rect 519629 145210 519695 145213
rect 523200 145210 524400 145240
rect 519629 145208 524400 145210
rect 116117 145150 119140 145152
rect 519629 145152 519634 145208
rect 519690 145152 524400 145208
rect 519629 145150 524400 145152
rect 116117 145147 116183 145150
rect 519629 145147 519695 145150
rect 523200 145120 524400 145150
rect 113817 144258 113883 144261
rect 110860 144256 113883 144258
rect 110860 144200 113822 144256
rect 113878 144200 113883 144256
rect 110860 144198 113883 144200
rect 113817 144195 113883 144198
rect 519813 143850 519879 143853
rect 518788 143848 519879 143850
rect 518788 143792 519818 143848
rect 519874 143792 519879 143848
rect 518788 143790 519879 143792
rect 519813 143787 519879 143790
rect 520917 143714 520983 143717
rect 523200 143714 524400 143744
rect 520917 143712 524400 143714
rect 520917 143656 520922 143712
rect 520978 143656 524400 143712
rect 520917 143654 524400 143656
rect 520917 143651 520983 143654
rect 523200 143624 524400 143654
rect 116025 143306 116091 143309
rect 116025 143304 119140 143306
rect 116025 143248 116030 143304
rect 116086 143248 119140 143304
rect 116025 143246 119140 143248
rect 116025 143243 116091 143246
rect 520089 142490 520155 142493
rect 518788 142488 520155 142490
rect 518788 142432 520094 142488
rect 520150 142432 520155 142488
rect 518788 142430 520155 142432
rect 520089 142427 520155 142430
rect 519537 142218 519603 142221
rect 523200 142218 524400 142248
rect 519537 142216 524400 142218
rect 519537 142160 519542 142216
rect 519598 142160 524400 142216
rect 519537 142158 524400 142160
rect 519537 142155 519603 142158
rect 523200 142128 524400 142158
rect 115289 141402 115355 141405
rect 115289 141400 119140 141402
rect 115289 141344 115294 141400
rect 115350 141344 119140 141400
rect 115289 141342 119140 141344
rect 115289 141339 115355 141342
rect 519997 141130 520063 141133
rect 518788 141128 520063 141130
rect 518788 141072 520002 141128
rect 520058 141072 520063 141128
rect 518788 141070 520063 141072
rect 519997 141067 520063 141070
rect 519353 140586 519419 140589
rect 523200 140586 524400 140616
rect 519353 140584 524400 140586
rect 519353 140528 519358 140584
rect 519414 140528 524400 140584
rect 519353 140526 524400 140528
rect 519353 140523 519419 140526
rect 523200 140496 524400 140526
rect 521009 139770 521075 139773
rect 518788 139768 521075 139770
rect 518788 139712 521014 139768
rect 521070 139712 521075 139768
rect 518788 139710 521075 139712
rect 521009 139707 521075 139710
rect 116117 139498 116183 139501
rect 116117 139496 119140 139498
rect 116117 139440 116122 139496
rect 116178 139440 119140 139496
rect 116117 139438 119140 139440
rect 116117 139435 116183 139438
rect 519997 139090 520063 139093
rect 523200 139090 524400 139120
rect 519997 139088 524400 139090
rect 519997 139032 520002 139088
rect 520058 139032 524400 139088
rect 519997 139030 524400 139032
rect 519997 139027 520063 139030
rect 523200 139000 524400 139030
rect 519445 138410 519511 138413
rect 518788 138408 519511 138410
rect 518788 138352 519450 138408
rect 519506 138352 519511 138408
rect 518788 138350 519511 138352
rect 519445 138347 519511 138350
rect 116117 137594 116183 137597
rect 520181 137594 520247 137597
rect 523200 137594 524400 137624
rect 116117 137592 119140 137594
rect 116117 137536 116122 137592
rect 116178 137536 119140 137592
rect 116117 137534 119140 137536
rect 520181 137592 524400 137594
rect 520181 137536 520186 137592
rect 520242 137536 524400 137592
rect 520181 137534 524400 137536
rect 116117 137531 116183 137534
rect 520181 137531 520247 137534
rect 523200 137504 524400 137534
rect 519905 137050 519971 137053
rect 518788 137048 519971 137050
rect 518788 136992 519910 137048
rect 519966 136992 519971 137048
rect 518788 136990 519971 136992
rect 519905 136987 519971 136990
rect 519445 136098 519511 136101
rect 523200 136098 524400 136128
rect 519445 136096 524400 136098
rect 519445 136040 519450 136096
rect 519506 136040 524400 136096
rect 519445 136038 524400 136040
rect 519445 136035 519511 136038
rect 523200 136008 524400 136038
rect 519721 135690 519787 135693
rect 518788 135688 519787 135690
rect 518788 135632 519726 135688
rect 519782 135632 519787 135688
rect 518788 135630 519787 135632
rect 519721 135627 519787 135630
rect 115197 135554 115263 135557
rect 115197 135552 119140 135554
rect 115197 135496 115202 135552
rect 115258 135496 119140 135552
rect 115197 135494 119140 135496
rect 115197 135491 115263 135494
rect 520089 134602 520155 134605
rect 523200 134602 524400 134632
rect 520089 134600 524400 134602
rect 520089 134544 520094 134600
rect 520150 134544 524400 134600
rect 520089 134542 524400 134544
rect 520089 134539 520155 134542
rect 523200 134512 524400 134542
rect 521101 134330 521167 134333
rect 518788 134328 521167 134330
rect 518788 134272 521106 134328
rect 521162 134272 521167 134328
rect 518788 134270 521167 134272
rect 521101 134267 521167 134270
rect 116025 133650 116091 133653
rect 116025 133648 119140 133650
rect 116025 133592 116030 133648
rect 116086 133592 119140 133648
rect 116025 133590 119140 133592
rect 116025 133587 116091 133590
rect 519813 133106 519879 133109
rect 523200 133106 524400 133136
rect 519813 133104 524400 133106
rect 519813 133048 519818 133104
rect 519874 133048 524400 133104
rect 519813 133046 524400 133048
rect 519813 133043 519879 133046
rect 523200 133016 524400 133046
rect 519629 132970 519695 132973
rect 518788 132968 519695 132970
rect 518788 132912 519634 132968
rect 519690 132912 519695 132968
rect 518788 132910 519695 132912
rect 519629 132907 519695 132910
rect 114185 132834 114251 132837
rect 110860 132832 114251 132834
rect 110860 132776 114190 132832
rect 114246 132776 114251 132832
rect 110860 132774 114251 132776
rect 114185 132771 114251 132774
rect 116117 131746 116183 131749
rect 520917 131746 520983 131749
rect 116117 131744 119140 131746
rect 116117 131688 116122 131744
rect 116178 131688 119140 131744
rect 116117 131686 119140 131688
rect 518758 131744 520983 131746
rect 518758 131688 520922 131744
rect 520978 131688 520983 131744
rect 518758 131686 520983 131688
rect 116117 131683 116183 131686
rect 518758 131580 518818 131686
rect 520917 131683 520983 131686
rect 519905 131610 519971 131613
rect 523200 131610 524400 131640
rect 519905 131608 524400 131610
rect 519905 131552 519910 131608
rect 519966 131552 524400 131608
rect 519905 131550 524400 131552
rect 519905 131547 519971 131550
rect 523200 131520 524400 131550
rect 519537 130250 519603 130253
rect 518788 130248 519603 130250
rect 518788 130192 519542 130248
rect 519598 130192 519603 130248
rect 518788 130190 519603 130192
rect 519537 130187 519603 130190
rect 519721 130114 519787 130117
rect 523200 130114 524400 130144
rect 519721 130112 524400 130114
rect 519721 130056 519726 130112
rect 519782 130056 524400 130112
rect 519721 130054 524400 130056
rect 519721 130051 519787 130054
rect 523200 130024 524400 130054
rect 116485 129842 116551 129845
rect 116485 129840 119140 129842
rect 116485 129784 116490 129840
rect 116546 129784 119140 129840
rect 116485 129782 119140 129784
rect 116485 129779 116551 129782
rect 519353 128890 519419 128893
rect 518788 128888 519419 128890
rect 518788 128832 519358 128888
rect 519414 128832 519419 128888
rect 518788 128830 519419 128832
rect 519353 128827 519419 128830
rect 519629 128618 519695 128621
rect 523200 128618 524400 128648
rect 519629 128616 524400 128618
rect 519629 128560 519634 128616
rect 519690 128560 524400 128616
rect 519629 128558 524400 128560
rect 519629 128555 519695 128558
rect 523200 128528 524400 128558
rect 117221 127938 117287 127941
rect 117221 127936 119140 127938
rect 117221 127880 117226 127936
rect 117282 127880 119140 127936
rect 117221 127878 119140 127880
rect 117221 127875 117287 127878
rect 519997 127530 520063 127533
rect 518788 127528 520063 127530
rect 518788 127472 520002 127528
rect 520058 127472 520063 127528
rect 518788 127470 520063 127472
rect 519997 127467 520063 127470
rect 519537 127122 519603 127125
rect 523200 127122 524400 127152
rect 519537 127120 524400 127122
rect 519537 127064 519542 127120
rect 519598 127064 524400 127120
rect 519537 127062 524400 127064
rect 519537 127059 519603 127062
rect 523200 127032 524400 127062
rect 520181 126170 520247 126173
rect 518788 126168 520247 126170
rect 518788 126112 520186 126168
rect 520242 126112 520247 126168
rect 518788 126110 520247 126112
rect 520181 126107 520247 126110
rect 116117 126034 116183 126037
rect 116117 126032 119140 126034
rect 116117 125976 116122 126032
rect 116178 125976 119140 126032
rect 116117 125974 119140 125976
rect 116117 125971 116183 125974
rect 519997 125626 520063 125629
rect 523200 125626 524400 125656
rect 519997 125624 524400 125626
rect 519997 125568 520002 125624
rect 520058 125568 524400 125624
rect 519997 125566 524400 125568
rect 519997 125563 520063 125566
rect 523200 125536 524400 125566
rect 519445 124810 519511 124813
rect 518788 124808 519511 124810
rect 518788 124752 519450 124808
rect 519506 124752 519511 124808
rect 518788 124750 519511 124752
rect 519445 124747 519511 124750
rect 116117 124130 116183 124133
rect 519261 124130 519327 124133
rect 523200 124130 524400 124160
rect 116117 124128 119140 124130
rect 116117 124072 116122 124128
rect 116178 124072 119140 124128
rect 116117 124070 119140 124072
rect 519261 124128 524400 124130
rect 519261 124072 519266 124128
rect 519322 124072 524400 124128
rect 519261 124070 524400 124072
rect 116117 124067 116183 124070
rect 519261 124067 519327 124070
rect 523200 124040 524400 124070
rect 520089 123450 520155 123453
rect 518788 123448 520155 123450
rect 518788 123392 520094 123448
rect 520150 123392 520155 123448
rect 518788 123390 520155 123392
rect 520089 123387 520155 123390
rect 519353 122634 519419 122637
rect 523200 122634 524400 122664
rect 519353 122632 524400 122634
rect 519353 122576 519358 122632
rect 519414 122576 524400 122632
rect 519353 122574 524400 122576
rect 519353 122571 519419 122574
rect 523200 122544 524400 122574
rect 115933 122226 115999 122229
rect 115933 122224 119140 122226
rect 115933 122168 115938 122224
rect 115994 122168 119140 122224
rect 115933 122166 119140 122168
rect 115933 122163 115999 122166
rect 519813 122090 519879 122093
rect 518788 122088 519879 122090
rect 518788 122032 519818 122088
rect 519874 122032 519879 122088
rect 518788 122030 519879 122032
rect 519813 122027 519879 122030
rect 113909 121410 113975 121413
rect 110860 121408 113975 121410
rect 110860 121352 113914 121408
rect 113970 121352 113975 121408
rect 110860 121350 113975 121352
rect 113909 121347 113975 121350
rect 520089 121138 520155 121141
rect 523200 121138 524400 121168
rect 520089 121136 524400 121138
rect 520089 121080 520094 121136
rect 520150 121080 524400 121136
rect 520089 121078 524400 121080
rect 520089 121075 520155 121078
rect 523200 121048 524400 121078
rect 519905 120730 519971 120733
rect 518788 120728 519971 120730
rect 518788 120672 519910 120728
rect 519966 120672 519971 120728
rect 518788 120670 519971 120672
rect 519905 120667 519971 120670
rect 116117 120186 116183 120189
rect 116117 120184 119140 120186
rect 116117 120128 116122 120184
rect 116178 120128 119140 120184
rect 116117 120126 119140 120128
rect 116117 120123 116183 120126
rect 519445 119642 519511 119645
rect 523200 119642 524400 119672
rect 519445 119640 524400 119642
rect 519445 119584 519450 119640
rect 519506 119584 524400 119640
rect 519445 119582 524400 119584
rect 519445 119579 519511 119582
rect 523200 119552 524400 119582
rect 519721 119370 519787 119373
rect 518788 119368 519787 119370
rect 518788 119312 519726 119368
rect 519782 119312 519787 119368
rect 518788 119310 519787 119312
rect 519721 119307 519787 119310
rect 116117 118282 116183 118285
rect 116117 118280 119140 118282
rect 116117 118224 116122 118280
rect 116178 118224 119140 118280
rect 116117 118222 119140 118224
rect 116117 118219 116183 118222
rect 519813 118146 519879 118149
rect 523200 118146 524400 118176
rect 519813 118144 524400 118146
rect 519813 118088 519818 118144
rect 519874 118088 524400 118144
rect 519813 118086 524400 118088
rect 519813 118083 519879 118086
rect 523200 118056 524400 118086
rect 519629 118010 519695 118013
rect 518788 118008 519695 118010
rect 518788 117952 519634 118008
rect 519690 117952 519695 118008
rect 518788 117950 519695 117952
rect 519629 117947 519695 117950
rect 519537 116650 519603 116653
rect 518788 116648 519603 116650
rect 518788 116592 519542 116648
rect 519598 116592 519603 116648
rect 518788 116590 519603 116592
rect 519537 116587 519603 116590
rect 519905 116514 519971 116517
rect 523200 116514 524400 116544
rect 519905 116512 524400 116514
rect 519905 116456 519910 116512
rect 519966 116456 524400 116512
rect 519905 116454 524400 116456
rect 519905 116451 519971 116454
rect 523200 116424 524400 116454
rect 116117 116378 116183 116381
rect 116117 116376 119140 116378
rect 116117 116320 116122 116376
rect 116178 116320 119140 116376
rect 116117 116318 119140 116320
rect 116117 116315 116183 116318
rect 519997 115290 520063 115293
rect 518788 115288 520063 115290
rect 518788 115232 520002 115288
rect 520058 115232 520063 115288
rect 518788 115230 520063 115232
rect 519997 115227 520063 115230
rect 520181 115018 520247 115021
rect 523200 115018 524400 115048
rect 520181 115016 524400 115018
rect 520181 114960 520186 115016
rect 520242 114960 524400 115016
rect 520181 114958 524400 114960
rect 520181 114955 520247 114958
rect 523200 114928 524400 114958
rect 116117 114474 116183 114477
rect 116117 114472 119140 114474
rect 116117 114416 116122 114472
rect 116178 114416 119140 114472
rect 116117 114414 119140 114416
rect 116117 114411 116183 114414
rect 519261 113930 519327 113933
rect 518788 113928 519327 113930
rect 518788 113872 519266 113928
rect 519322 113872 519327 113928
rect 518788 113870 519327 113872
rect 519261 113867 519327 113870
rect 519721 113522 519787 113525
rect 523200 113522 524400 113552
rect 519721 113520 524400 113522
rect 519721 113464 519726 113520
rect 519782 113464 524400 113520
rect 519721 113462 524400 113464
rect 519721 113459 519787 113462
rect 523200 113432 524400 113462
rect 115933 112570 115999 112573
rect 519353 112570 519419 112573
rect 115933 112568 119140 112570
rect 115933 112512 115938 112568
rect 115994 112512 119140 112568
rect 115933 112510 119140 112512
rect 518788 112568 519419 112570
rect 518788 112512 519358 112568
rect 519414 112512 519419 112568
rect 518788 112510 519419 112512
rect 115933 112507 115999 112510
rect 519353 112507 519419 112510
rect 519629 112026 519695 112029
rect 523200 112026 524400 112056
rect 519629 112024 524400 112026
rect 519629 111968 519634 112024
rect 519690 111968 524400 112024
rect 519629 111966 524400 111968
rect 519629 111963 519695 111966
rect 523200 111936 524400 111966
rect 520089 111210 520155 111213
rect 518788 111208 520155 111210
rect 518788 111152 520094 111208
rect 520150 111152 520155 111208
rect 518788 111150 520155 111152
rect 520089 111147 520155 111150
rect 116117 110666 116183 110669
rect 116117 110664 119140 110666
rect 116117 110608 116122 110664
rect 116178 110608 119140 110664
rect 116117 110606 119140 110608
rect 116117 110603 116183 110606
rect 519537 110530 519603 110533
rect 523200 110530 524400 110560
rect 519537 110528 524400 110530
rect 519537 110472 519542 110528
rect 519598 110472 524400 110528
rect 519537 110470 524400 110472
rect 519537 110467 519603 110470
rect 523200 110440 524400 110470
rect 114001 110122 114067 110125
rect 110860 110120 114067 110122
rect 110860 110064 114006 110120
rect 114062 110064 114067 110120
rect 110860 110062 114067 110064
rect 114001 110059 114067 110062
rect 519445 109850 519511 109853
rect 518788 109848 519511 109850
rect 518788 109792 519450 109848
rect 519506 109792 519511 109848
rect 518788 109790 519511 109792
rect 519445 109787 519511 109790
rect 521285 109034 521351 109037
rect 523200 109034 524400 109064
rect 521285 109032 524400 109034
rect 521285 108976 521290 109032
rect 521346 108976 524400 109032
rect 521285 108974 524400 108976
rect 521285 108971 521351 108974
rect 523200 108944 524400 108974
rect 116117 108762 116183 108765
rect 116117 108760 119140 108762
rect 116117 108704 116122 108760
rect 116178 108704 119140 108760
rect 116117 108702 119140 108704
rect 116117 108699 116183 108702
rect 519813 108490 519879 108493
rect 518788 108488 519879 108490
rect 518788 108432 519818 108488
rect 519874 108432 519879 108488
rect 518788 108430 519879 108432
rect 519813 108427 519879 108430
rect 521101 107538 521167 107541
rect 523200 107538 524400 107568
rect 521101 107536 524400 107538
rect 521101 107480 521106 107536
rect 521162 107480 524400 107536
rect 521101 107478 524400 107480
rect 521101 107475 521167 107478
rect 523200 107448 524400 107478
rect 519905 107130 519971 107133
rect 518788 107128 519971 107130
rect 518788 107072 519910 107128
rect 519966 107072 519971 107128
rect 518788 107070 519971 107072
rect 519905 107067 519971 107070
rect 110321 106314 110387 106317
rect 119110 106314 119170 106828
rect 110321 106312 119170 106314
rect 110321 106256 110326 106312
rect 110382 106256 119170 106312
rect 110321 106254 119170 106256
rect 110321 106251 110387 106254
rect 520273 106042 520339 106045
rect 523200 106042 524400 106072
rect 520273 106040 524400 106042
rect 520273 105984 520278 106040
rect 520334 105984 524400 106040
rect 520273 105982 524400 105984
rect 520273 105979 520339 105982
rect 523200 105952 524400 105982
rect 520181 105770 520247 105773
rect 518788 105768 520247 105770
rect 518788 105712 520186 105768
rect 520242 105712 520247 105768
rect 518788 105710 520247 105712
rect 520181 105707 520247 105710
rect 117129 104818 117195 104821
rect 117129 104816 119140 104818
rect 117129 104760 117134 104816
rect 117190 104760 119140 104816
rect 117129 104758 119140 104760
rect 117129 104755 117195 104758
rect 521009 104546 521075 104549
rect 523200 104546 524400 104576
rect 521009 104544 524400 104546
rect 521009 104488 521014 104544
rect 521070 104488 524400 104544
rect 521009 104486 524400 104488
rect 521009 104483 521075 104486
rect 523200 104456 524400 104486
rect 519721 104410 519787 104413
rect 518788 104408 519787 104410
rect 518788 104352 519726 104408
rect 519782 104352 519787 104408
rect 518788 104350 519787 104352
rect 519721 104347 519787 104350
rect 519629 103050 519695 103053
rect 518788 103048 519695 103050
rect 518788 102992 519634 103048
rect 519690 102992 519695 103048
rect 518788 102990 519695 102992
rect 519629 102987 519695 102990
rect 521193 103050 521259 103053
rect 523200 103050 524400 103080
rect 521193 103048 524400 103050
rect 521193 102992 521198 103048
rect 521254 102992 524400 103048
rect 521193 102990 524400 102992
rect 521193 102987 521259 102990
rect 523200 102960 524400 102990
rect 116945 102914 117011 102917
rect 116945 102912 119140 102914
rect 116945 102856 116950 102912
rect 117006 102856 119140 102912
rect 116945 102854 119140 102856
rect 116945 102851 117011 102854
rect 519537 101690 519603 101693
rect 518788 101688 519603 101690
rect 518788 101632 519542 101688
rect 519598 101632 519603 101688
rect 518788 101630 519603 101632
rect 519537 101627 519603 101630
rect 520917 101554 520983 101557
rect 523200 101554 524400 101584
rect 520917 101552 524400 101554
rect 520917 101496 520922 101552
rect 520978 101496 524400 101552
rect 520917 101494 524400 101496
rect 520917 101491 520983 101494
rect 523200 101464 524400 101494
rect 117037 101010 117103 101013
rect 117037 101008 119140 101010
rect 117037 100952 117042 101008
rect 117098 100952 119140 101008
rect 117037 100950 119140 100952
rect 117037 100947 117103 100950
rect 521285 100330 521351 100333
rect 518788 100328 521351 100330
rect 518788 100272 521290 100328
rect 521346 100272 521351 100328
rect 518788 100270 521351 100272
rect 521285 100267 521351 100270
rect 521469 100058 521535 100061
rect 523200 100058 524400 100088
rect 521469 100056 524400 100058
rect 521469 100000 521474 100056
rect 521530 100000 524400 100056
rect 521469 99998 524400 100000
rect 521469 99995 521535 99998
rect 523200 99968 524400 99998
rect 116853 99106 116919 99109
rect 116853 99104 119140 99106
rect 116853 99048 116858 99104
rect 116914 99048 119140 99104
rect 116853 99046 119140 99048
rect 116853 99043 116919 99046
rect 521101 98970 521167 98973
rect 518788 98968 521167 98970
rect 518788 98912 521106 98968
rect 521162 98912 521167 98968
rect 518788 98910 521167 98912
rect 521101 98907 521167 98910
rect 114093 98698 114159 98701
rect 110860 98696 114159 98698
rect 110860 98640 114098 98696
rect 114154 98640 114159 98696
rect 110860 98638 114159 98640
rect 114093 98635 114159 98638
rect 521285 98562 521351 98565
rect 523200 98562 524400 98592
rect 521285 98560 524400 98562
rect 521285 98504 521290 98560
rect 521346 98504 524400 98560
rect 521285 98502 524400 98504
rect 521285 98499 521351 98502
rect 523200 98472 524400 98502
rect 520273 97610 520339 97613
rect 518788 97608 520339 97610
rect 518788 97552 520278 97608
rect 520334 97552 520339 97608
rect 518788 97550 520339 97552
rect 520273 97547 520339 97550
rect 116761 97202 116827 97205
rect 116761 97200 119140 97202
rect 116761 97144 116766 97200
rect 116822 97144 119140 97200
rect 116761 97142 119140 97144
rect 116761 97139 116827 97142
rect 521377 97066 521443 97069
rect 523200 97066 524400 97096
rect 521377 97064 524400 97066
rect 521377 97008 521382 97064
rect 521438 97008 524400 97064
rect 521377 97006 524400 97008
rect 521377 97003 521443 97006
rect 523200 96976 524400 97006
rect 521009 96250 521075 96253
rect 518788 96248 521075 96250
rect 518788 96192 521014 96248
rect 521070 96192 521075 96248
rect 518788 96190 521075 96192
rect 521009 96187 521075 96190
rect 520273 95570 520339 95573
rect 523200 95570 524400 95600
rect 520273 95568 524400 95570
rect 520273 95512 520278 95568
rect 520334 95512 524400 95568
rect 520273 95510 524400 95512
rect 520273 95507 520339 95510
rect 523200 95480 524400 95510
rect 116669 95298 116735 95301
rect 116669 95296 119140 95298
rect 116669 95240 116674 95296
rect 116730 95240 119140 95296
rect 116669 95238 119140 95240
rect 116669 95235 116735 95238
rect 521193 94890 521259 94893
rect 518788 94888 521259 94890
rect 518788 94832 521198 94888
rect 521254 94832 521259 94888
rect 518788 94830 521259 94832
rect 521193 94827 521259 94830
rect 521009 93938 521075 93941
rect 523200 93938 524400 93968
rect 521009 93936 524400 93938
rect 521009 93880 521014 93936
rect 521070 93880 524400 93936
rect 521009 93878 524400 93880
rect 521009 93875 521075 93878
rect 523200 93848 524400 93878
rect 520917 93530 520983 93533
rect 518788 93528 520983 93530
rect 518788 93472 520922 93528
rect 520978 93472 520983 93528
rect 518788 93470 520983 93472
rect 520917 93467 520983 93470
rect 116577 93394 116643 93397
rect 116577 93392 119140 93394
rect 116577 93336 116582 93392
rect 116638 93336 119140 93392
rect 116577 93334 119140 93336
rect 116577 93331 116643 93334
rect 519629 92442 519695 92445
rect 523200 92442 524400 92472
rect 519629 92440 524400 92442
rect 519629 92384 519634 92440
rect 519690 92384 524400 92440
rect 519629 92382 524400 92384
rect 519629 92379 519695 92382
rect 523200 92352 524400 92382
rect 521469 92170 521535 92173
rect 518788 92168 521535 92170
rect 518788 92112 521474 92168
rect 521530 92112 521535 92168
rect 518788 92110 521535 92112
rect 521469 92107 521535 92110
rect 116117 91354 116183 91357
rect 116117 91352 119140 91354
rect 116117 91296 116122 91352
rect 116178 91296 119140 91352
rect 116117 91294 119140 91296
rect 116117 91291 116183 91294
rect 519997 90946 520063 90949
rect 523200 90946 524400 90976
rect 519997 90944 524400 90946
rect 519997 90888 520002 90944
rect 520058 90888 524400 90944
rect 519997 90886 524400 90888
rect 519997 90883 520063 90886
rect 523200 90856 524400 90886
rect 521285 90810 521351 90813
rect 518788 90808 521351 90810
rect 518788 90752 521290 90808
rect 521346 90752 521351 90808
rect 518788 90750 521351 90752
rect 521285 90747 521351 90750
rect 521377 89586 521443 89589
rect 518758 89584 521443 89586
rect 518758 89528 521382 89584
rect 521438 89528 521443 89584
rect 518758 89526 521443 89528
rect 116117 89450 116183 89453
rect 116117 89448 119140 89450
rect 116117 89392 116122 89448
rect 116178 89392 119140 89448
rect 518758 89420 518818 89526
rect 521377 89523 521443 89526
rect 519721 89450 519787 89453
rect 523200 89450 524400 89480
rect 519721 89448 524400 89450
rect 116117 89390 119140 89392
rect 519721 89392 519726 89448
rect 519782 89392 524400 89448
rect 519721 89390 524400 89392
rect 116117 89387 116183 89390
rect 519721 89387 519787 89390
rect 523200 89360 524400 89390
rect 520273 88090 520339 88093
rect 518788 88088 520339 88090
rect 518788 88032 520278 88088
rect 520334 88032 520339 88088
rect 518788 88030 520339 88032
rect 520273 88027 520339 88030
rect 519905 87954 519971 87957
rect 523200 87954 524400 87984
rect 519905 87952 524400 87954
rect 519905 87896 519910 87952
rect 519966 87896 524400 87952
rect 519905 87894 524400 87896
rect 519905 87891 519971 87894
rect 523200 87864 524400 87894
rect 116025 87546 116091 87549
rect 116025 87544 119140 87546
rect 116025 87488 116030 87544
rect 116086 87488 119140 87544
rect 116025 87486 119140 87488
rect 116025 87483 116091 87486
rect 114185 87274 114251 87277
rect 110860 87272 114251 87274
rect 110860 87216 114190 87272
rect 114246 87216 114251 87272
rect 110860 87214 114251 87216
rect 114185 87211 114251 87214
rect 521009 86730 521075 86733
rect 518788 86728 521075 86730
rect 518788 86672 521014 86728
rect 521070 86672 521075 86728
rect 518788 86670 521075 86672
rect 521009 86667 521075 86670
rect 519813 86458 519879 86461
rect 523200 86458 524400 86488
rect 519813 86456 524400 86458
rect 519813 86400 519818 86456
rect 519874 86400 524400 86456
rect 519813 86398 524400 86400
rect 519813 86395 519879 86398
rect 523200 86368 524400 86398
rect 115197 85642 115263 85645
rect 115197 85640 119140 85642
rect 115197 85584 115202 85640
rect 115258 85584 119140 85640
rect 115197 85582 119140 85584
rect 115197 85579 115263 85582
rect 519629 85370 519695 85373
rect 518788 85368 519695 85370
rect 518788 85312 519634 85368
rect 519690 85312 519695 85368
rect 518788 85310 519695 85312
rect 519629 85307 519695 85310
rect 519077 84962 519143 84965
rect 523200 84962 524400 84992
rect 519077 84960 524400 84962
rect 519077 84904 519082 84960
rect 519138 84904 524400 84960
rect 519077 84902 524400 84904
rect 519077 84899 519143 84902
rect 523200 84872 524400 84902
rect 519997 84010 520063 84013
rect 518788 84008 520063 84010
rect 518788 83952 520002 84008
rect 520058 83952 520063 84008
rect 518788 83950 520063 83952
rect 519997 83947 520063 83950
rect 116577 83738 116643 83741
rect 116577 83736 119140 83738
rect 116577 83680 116582 83736
rect 116638 83680 119140 83736
rect 116577 83678 119140 83680
rect 116577 83675 116643 83678
rect 520089 83466 520155 83469
rect 523200 83466 524400 83496
rect 520089 83464 524400 83466
rect 520089 83408 520094 83464
rect 520150 83408 524400 83464
rect 520089 83406 524400 83408
rect 520089 83403 520155 83406
rect 523200 83376 524400 83406
rect 519721 82650 519787 82653
rect 518788 82648 519787 82650
rect 518788 82592 519726 82648
rect 519782 82592 519787 82648
rect 518788 82590 519787 82592
rect 519721 82587 519787 82590
rect 519445 81970 519511 81973
rect 523200 81970 524400 82000
rect 519445 81968 524400 81970
rect 519445 81912 519450 81968
rect 519506 81912 524400 81968
rect 519445 81910 524400 81912
rect 519445 81907 519511 81910
rect 523200 81880 524400 81910
rect 116209 81834 116275 81837
rect 116209 81832 119140 81834
rect 116209 81776 116214 81832
rect 116270 81776 119140 81832
rect 116209 81774 119140 81776
rect 116209 81771 116275 81774
rect 519905 81290 519971 81293
rect 518788 81288 519971 81290
rect 518788 81232 519910 81288
rect 519966 81232 519971 81288
rect 518788 81230 519971 81232
rect 519905 81227 519971 81230
rect 520181 80474 520247 80477
rect 523200 80474 524400 80504
rect 520181 80472 524400 80474
rect 520181 80416 520186 80472
rect 520242 80416 524400 80472
rect 520181 80414 524400 80416
rect 520181 80411 520247 80414
rect 523200 80384 524400 80414
rect 115933 79930 115999 79933
rect 519813 79930 519879 79933
rect 115933 79928 119140 79930
rect 115933 79872 115938 79928
rect 115994 79872 119140 79928
rect 115933 79870 119140 79872
rect 518788 79928 519879 79930
rect 518788 79872 519818 79928
rect 519874 79872 519879 79928
rect 518788 79870 519879 79872
rect 115933 79867 115999 79870
rect 519813 79867 519879 79870
rect 519997 78978 520063 78981
rect 523200 78978 524400 79008
rect 519997 78976 524400 78978
rect 519997 78920 520002 78976
rect 520058 78920 524400 78976
rect 519997 78918 524400 78920
rect 519997 78915 520063 78918
rect 523200 78888 524400 78918
rect 519077 78570 519143 78573
rect 518788 78568 519143 78570
rect 518788 78512 519082 78568
rect 519138 78512 519143 78568
rect 518788 78510 519143 78512
rect 519077 78507 519143 78510
rect 116117 78026 116183 78029
rect 116117 78024 119140 78026
rect 116117 77968 116122 78024
rect 116178 77968 119140 78024
rect 116117 77966 119140 77968
rect 116117 77963 116183 77966
rect 519813 77482 519879 77485
rect 523200 77482 524400 77512
rect 519813 77480 524400 77482
rect 519813 77424 519818 77480
rect 519874 77424 524400 77480
rect 519813 77422 524400 77424
rect 519813 77419 519879 77422
rect 523200 77392 524400 77422
rect 520089 77210 520155 77213
rect 518788 77208 520155 77210
rect 518788 77152 520094 77208
rect 520150 77152 520155 77208
rect 518788 77150 520155 77152
rect 520089 77147 520155 77150
rect 519445 75986 519511 75989
rect 110860 75926 119140 75986
rect 518788 75984 519511 75986
rect 518788 75928 519450 75984
rect 519506 75928 519511 75984
rect 518788 75926 519511 75928
rect 519445 75923 519511 75926
rect 519905 75986 519971 75989
rect 523200 75986 524400 76016
rect 519905 75984 524400 75986
rect 519905 75928 519910 75984
rect 519966 75928 524400 75984
rect 519905 75926 524400 75928
rect 519905 75923 519971 75926
rect 523200 75896 524400 75926
rect 520181 74626 520247 74629
rect 518788 74624 520247 74626
rect 518788 74568 520186 74624
rect 520242 74568 520247 74624
rect 518788 74566 520247 74568
rect 520181 74563 520247 74566
rect 521101 74490 521167 74493
rect 523200 74490 524400 74520
rect 521101 74488 524400 74490
rect 521101 74432 521106 74488
rect 521162 74432 524400 74488
rect 521101 74430 524400 74432
rect 521101 74427 521167 74430
rect 523200 74400 524400 74430
rect 116669 74082 116735 74085
rect 116669 74080 119140 74082
rect 116669 74024 116674 74080
rect 116730 74024 119140 74080
rect 116669 74022 119140 74024
rect 116669 74019 116735 74022
rect 519997 73266 520063 73269
rect 518788 73264 520063 73266
rect 518788 73208 520002 73264
rect 520058 73208 520063 73264
rect 518788 73206 520063 73208
rect 519997 73203 520063 73206
rect 520917 72994 520983 72997
rect 523200 72994 524400 73024
rect 520917 72992 524400 72994
rect 520917 72936 520922 72992
rect 520978 72936 524400 72992
rect 520917 72934 524400 72936
rect 520917 72931 520983 72934
rect 523200 72904 524400 72934
rect 116577 72178 116643 72181
rect 116577 72176 119140 72178
rect 116577 72120 116582 72176
rect 116638 72120 119140 72176
rect 116577 72118 119140 72120
rect 116577 72115 116643 72118
rect 519813 71906 519879 71909
rect 518788 71904 519879 71906
rect 518788 71848 519818 71904
rect 519874 71848 519879 71904
rect 518788 71846 519879 71848
rect 519813 71843 519879 71846
rect 521193 71498 521259 71501
rect 523200 71498 524400 71528
rect 521193 71496 524400 71498
rect 521193 71440 521198 71496
rect 521254 71440 524400 71496
rect 521193 71438 524400 71440
rect 521193 71435 521259 71438
rect 523200 71408 524400 71438
rect 519905 70546 519971 70549
rect 518788 70544 519971 70546
rect 518788 70488 519910 70544
rect 519966 70488 519971 70544
rect 518788 70486 519971 70488
rect 519905 70483 519971 70486
rect 116301 70274 116367 70277
rect 116301 70272 119140 70274
rect 116301 70216 116306 70272
rect 116362 70216 119140 70272
rect 116301 70214 119140 70216
rect 116301 70211 116367 70214
rect 521009 69866 521075 69869
rect 523200 69866 524400 69896
rect 521009 69864 524400 69866
rect 521009 69808 521014 69864
rect 521070 69808 524400 69864
rect 521009 69806 524400 69808
rect 521009 69803 521075 69806
rect 523200 69776 524400 69806
rect 521101 69186 521167 69189
rect 518788 69184 521167 69186
rect 518788 69128 521106 69184
rect 521162 69128 521167 69184
rect 518788 69126 521167 69128
rect 521101 69123 521167 69126
rect 116117 68370 116183 68373
rect 521101 68370 521167 68373
rect 523200 68370 524400 68400
rect 116117 68368 119140 68370
rect 116117 68312 116122 68368
rect 116178 68312 119140 68368
rect 116117 68310 119140 68312
rect 521101 68368 524400 68370
rect 521101 68312 521106 68368
rect 521162 68312 524400 68368
rect 521101 68310 524400 68312
rect 116117 68307 116183 68310
rect 521101 68307 521167 68310
rect 523200 68280 524400 68310
rect 520917 67826 520983 67829
rect 518788 67824 520983 67826
rect 518788 67768 520922 67824
rect 520978 67768 520983 67824
rect 518788 67766 520983 67768
rect 520917 67763 520983 67766
rect 520457 66874 520523 66877
rect 523200 66874 524400 66904
rect 520457 66872 524400 66874
rect 520457 66816 520462 66872
rect 520518 66816 524400 66872
rect 520457 66814 524400 66816
rect 520457 66811 520523 66814
rect 523200 66784 524400 66814
rect 116577 66466 116643 66469
rect 521193 66466 521259 66469
rect 116577 66464 119140 66466
rect 116577 66408 116582 66464
rect 116638 66408 119140 66464
rect 116577 66406 119140 66408
rect 518788 66464 521259 66466
rect 518788 66408 521198 66464
rect 521254 66408 521259 66464
rect 518788 66406 521259 66408
rect 116577 66403 116643 66406
rect 521193 66403 521259 66406
rect 520365 65378 520431 65381
rect 523200 65378 524400 65408
rect 520365 65376 524400 65378
rect 520365 65320 520370 65376
rect 520426 65320 524400 65376
rect 520365 65318 524400 65320
rect 520365 65315 520431 65318
rect 523200 65288 524400 65318
rect 521009 65106 521075 65109
rect 518788 65104 521075 65106
rect 518788 65048 521014 65104
rect 521070 65048 521075 65104
rect 518788 65046 521075 65048
rect 521009 65043 521075 65046
rect 113357 64562 113423 64565
rect 110860 64560 113423 64562
rect 110860 64504 113362 64560
rect 113418 64504 113423 64560
rect 110860 64502 113423 64504
rect 113357 64499 113423 64502
rect 116209 64562 116275 64565
rect 116209 64560 119140 64562
rect 116209 64504 116214 64560
rect 116270 64504 119140 64560
rect 116209 64502 119140 64504
rect 116209 64499 116275 64502
rect 521193 63882 521259 63885
rect 523200 63882 524400 63912
rect 521193 63880 524400 63882
rect 521193 63824 521198 63880
rect 521254 63824 524400 63880
rect 521193 63822 524400 63824
rect 521193 63819 521259 63822
rect 523200 63792 524400 63822
rect 521101 63746 521167 63749
rect 518788 63744 521167 63746
rect 518788 63688 521106 63744
rect 521162 63688 521167 63744
rect 518788 63686 521167 63688
rect 521101 63683 521167 63686
rect 116117 62658 116183 62661
rect 116117 62656 119140 62658
rect 116117 62600 116122 62656
rect 116178 62600 119140 62656
rect 116117 62598 119140 62600
rect 116117 62595 116183 62598
rect 520457 62386 520523 62389
rect 518788 62384 520523 62386
rect 518788 62328 520462 62384
rect 520518 62328 520523 62384
rect 518788 62326 520523 62328
rect 520457 62323 520523 62326
rect 521009 62386 521075 62389
rect 523200 62386 524400 62416
rect 521009 62384 524400 62386
rect 521009 62328 521014 62384
rect 521070 62328 524400 62384
rect 521009 62326 524400 62328
rect 521009 62323 521075 62326
rect 523200 62296 524400 62326
rect 520365 61026 520431 61029
rect 518788 61024 520431 61026
rect 518788 60968 520370 61024
rect 520426 60968 520431 61024
rect 518788 60966 520431 60968
rect 520365 60963 520431 60966
rect 520733 60890 520799 60893
rect 523200 60890 524400 60920
rect 520733 60888 524400 60890
rect 520733 60832 520738 60888
rect 520794 60832 524400 60888
rect 520733 60830 524400 60832
rect 520733 60827 520799 60830
rect 523200 60800 524400 60830
rect 116577 60618 116643 60621
rect 116577 60616 119140 60618
rect 116577 60560 116582 60616
rect 116638 60560 119140 60616
rect 116577 60558 119140 60560
rect 116577 60555 116643 60558
rect 521193 59666 521259 59669
rect 518788 59664 521259 59666
rect 518788 59608 521198 59664
rect 521254 59608 521259 59664
rect 518788 59606 521259 59608
rect 521193 59603 521259 59606
rect 521101 59394 521167 59397
rect 523200 59394 524400 59424
rect 521101 59392 524400 59394
rect 521101 59336 521106 59392
rect 521162 59336 524400 59392
rect 521101 59334 524400 59336
rect 521101 59331 521167 59334
rect 523200 59304 524400 59334
rect 116761 58714 116827 58717
rect 116761 58712 119140 58714
rect 116761 58656 116766 58712
rect 116822 58656 119140 58712
rect 116761 58654 119140 58656
rect 116761 58651 116827 58654
rect 521009 58306 521075 58309
rect 518788 58304 521075 58306
rect 518788 58248 521014 58304
rect 521070 58248 521075 58304
rect 518788 58246 521075 58248
rect 521009 58243 521075 58246
rect 519905 57898 519971 57901
rect 523200 57898 524400 57928
rect 519905 57896 524400 57898
rect 519905 57840 519910 57896
rect 519966 57840 524400 57896
rect 519905 57838 524400 57840
rect 519905 57835 519971 57838
rect 523200 57808 524400 57838
rect 520733 56946 520799 56949
rect 518788 56944 520799 56946
rect 518788 56888 520738 56944
rect 520794 56888 520799 56944
rect 518788 56886 520799 56888
rect 520733 56883 520799 56886
rect 116669 56810 116735 56813
rect 116669 56808 119140 56810
rect 116669 56752 116674 56808
rect 116730 56752 119140 56808
rect 116669 56750 119140 56752
rect 116669 56747 116735 56750
rect 519813 56402 519879 56405
rect 523200 56402 524400 56432
rect 519813 56400 524400 56402
rect 519813 56344 519818 56400
rect 519874 56344 524400 56400
rect 519813 56342 524400 56344
rect 519813 56339 519879 56342
rect 523200 56312 524400 56342
rect 521101 55586 521167 55589
rect 518788 55584 521167 55586
rect 518788 55528 521106 55584
rect 521162 55528 521167 55584
rect 518788 55526 521167 55528
rect 521101 55523 521167 55526
rect 520181 54906 520247 54909
rect 523200 54906 524400 54936
rect 520181 54904 524400 54906
rect 110321 53954 110387 53957
rect 119110 53954 119170 54876
rect 520181 54848 520186 54904
rect 520242 54848 524400 54904
rect 520181 54846 524400 54848
rect 520181 54843 520247 54846
rect 523200 54816 524400 54846
rect 519905 54226 519971 54229
rect 518788 54224 519971 54226
rect 518788 54168 519910 54224
rect 519966 54168 519971 54224
rect 518788 54166 519971 54168
rect 519905 54163 519971 54166
rect 110321 53952 119170 53954
rect 110321 53896 110326 53952
rect 110382 53896 119170 53952
rect 110321 53894 119170 53896
rect 110321 53891 110387 53894
rect 519077 53410 519143 53413
rect 523200 53410 524400 53440
rect 519077 53408 524400 53410
rect 519077 53352 519082 53408
rect 519138 53352 524400 53408
rect 519077 53350 524400 53352
rect 519077 53347 519143 53350
rect 523200 53320 524400 53350
rect 114185 53138 114251 53141
rect 110860 53136 114251 53138
rect 110860 53080 114190 53136
rect 114246 53080 114251 53136
rect 110860 53078 114251 53080
rect 114185 53075 114251 53078
rect 110321 52594 110387 52597
rect 119110 52594 119170 52972
rect 519813 52866 519879 52869
rect 518788 52864 519879 52866
rect 518788 52808 519818 52864
rect 519874 52808 519879 52864
rect 518788 52806 519879 52808
rect 519813 52803 519879 52806
rect 110321 52592 119170 52594
rect 110321 52536 110326 52592
rect 110382 52536 119170 52592
rect 110321 52534 119170 52536
rect 110321 52531 110387 52534
rect 520089 51914 520155 51917
rect 523200 51914 524400 51944
rect 520089 51912 524400 51914
rect 520089 51856 520094 51912
rect 520150 51856 524400 51912
rect 520089 51854 524400 51856
rect 520089 51851 520155 51854
rect 523200 51824 524400 51854
rect 520181 51506 520247 51509
rect 518788 51504 520247 51506
rect 518788 51448 520186 51504
rect 520242 51448 520247 51504
rect 518788 51446 520247 51448
rect 520181 51443 520247 51446
rect 110321 51098 110387 51101
rect 110321 51096 119140 51098
rect 110321 51040 110326 51096
rect 110382 51040 119140 51096
rect 110321 51038 119140 51040
rect 110321 51035 110387 51038
rect 520181 50418 520247 50421
rect 523200 50418 524400 50448
rect 520181 50416 524400 50418
rect 520181 50360 520186 50416
rect 520242 50360 524400 50416
rect 520181 50358 524400 50360
rect 520181 50355 520247 50358
rect 523200 50328 524400 50358
rect 519077 50146 519143 50149
rect 518788 50144 519143 50146
rect 518788 50088 519082 50144
rect 519138 50088 519143 50144
rect 518788 50086 519143 50088
rect 519077 50083 519143 50086
rect 110321 48378 110387 48381
rect 119110 48378 119170 49164
rect 519077 48922 519143 48925
rect 523200 48922 524400 48952
rect 519077 48920 524400 48922
rect 519077 48864 519082 48920
rect 519138 48864 524400 48920
rect 519077 48862 524400 48864
rect 519077 48859 519143 48862
rect 523200 48832 524400 48862
rect 520089 48786 520155 48789
rect 518788 48784 520155 48786
rect 518788 48728 520094 48784
rect 520150 48728 520155 48784
rect 518788 48726 520155 48728
rect 520089 48723 520155 48726
rect 110321 48376 119170 48378
rect 110321 48320 110326 48376
rect 110382 48320 119170 48376
rect 110321 48318 119170 48320
rect 110321 48315 110387 48318
rect 520181 47426 520247 47429
rect 518788 47424 520247 47426
rect 518788 47368 520186 47424
rect 520242 47368 520247 47424
rect 518788 47366 520247 47368
rect 520181 47363 520247 47366
rect 519905 47290 519971 47293
rect 523200 47290 524400 47320
rect 519905 47288 524400 47290
rect 519905 47232 519910 47288
rect 519966 47232 524400 47288
rect 519905 47230 524400 47232
rect 519905 47227 519971 47230
rect 523200 47200 524400 47230
rect 110321 47154 110387 47157
rect 110321 47152 119140 47154
rect 110321 47096 110326 47152
rect 110382 47096 119140 47152
rect 110321 47094 119140 47096
rect 110321 47091 110387 47094
rect 519077 46066 519143 46069
rect 518788 46064 519143 46066
rect 518788 46008 519082 46064
rect 519138 46008 519143 46064
rect 518788 46006 519143 46008
rect 519077 46003 519143 46006
rect 519721 45794 519787 45797
rect 523200 45794 524400 45824
rect 519721 45792 524400 45794
rect 519721 45736 519726 45792
rect 519782 45736 524400 45792
rect 519721 45734 524400 45736
rect 519721 45731 519787 45734
rect 523200 45704 524400 45734
rect 110321 44298 110387 44301
rect 119110 44298 119170 45220
rect 519905 44706 519971 44709
rect 518788 44704 519971 44706
rect 518788 44648 519910 44704
rect 519966 44648 519971 44704
rect 518788 44646 519971 44648
rect 519905 44643 519971 44646
rect 110321 44296 119170 44298
rect 110321 44240 110326 44296
rect 110382 44240 119170 44296
rect 110321 44238 119170 44240
rect 520181 44298 520247 44301
rect 523200 44298 524400 44328
rect 520181 44296 524400 44298
rect 520181 44240 520186 44296
rect 520242 44240 524400 44296
rect 520181 44238 524400 44240
rect 110321 44235 110387 44238
rect 520181 44235 520247 44238
rect 523200 44208 524400 44238
rect 116117 43346 116183 43349
rect 519721 43346 519787 43349
rect 116117 43344 119140 43346
rect 116117 43288 116122 43344
rect 116178 43288 119140 43344
rect 116117 43286 119140 43288
rect 518788 43344 519787 43346
rect 518788 43288 519726 43344
rect 519782 43288 519787 43344
rect 518788 43286 519787 43288
rect 116117 43283 116183 43286
rect 519721 43283 519787 43286
rect 520733 42802 520799 42805
rect 523200 42802 524400 42832
rect 520733 42800 524400 42802
rect 520733 42744 520738 42800
rect 520794 42744 524400 42800
rect 520733 42742 524400 42744
rect 520733 42739 520799 42742
rect 523200 42712 524400 42742
rect 520181 41986 520247 41989
rect 518788 41984 520247 41986
rect 518788 41928 520186 41984
rect 520242 41928 520247 41984
rect 518788 41926 520247 41928
rect 520181 41923 520247 41926
rect 114093 41850 114159 41853
rect 110860 41848 114159 41850
rect 110860 41792 114098 41848
rect 114154 41792 114159 41848
rect 110860 41790 114159 41792
rect 114093 41787 114159 41790
rect 110321 41442 110387 41445
rect 110321 41440 119140 41442
rect 110321 41384 110326 41440
rect 110382 41384 119140 41440
rect 110321 41382 119140 41384
rect 110321 41379 110387 41382
rect 520733 41306 520799 41309
rect 518758 41304 520799 41306
rect 518758 41248 520738 41304
rect 520794 41248 520799 41304
rect 518758 41246 520799 41248
rect 518758 40596 518818 41246
rect 520733 41243 520799 41246
rect 520917 41306 520983 41309
rect 523200 41306 524400 41336
rect 520917 41304 524400 41306
rect 520917 41248 520922 41304
rect 520978 41248 524400 41304
rect 520917 41246 524400 41248
rect 520917 41243 520983 41246
rect 523200 41216 524400 41246
rect 520917 39946 520983 39949
rect 518758 39944 520983 39946
rect 518758 39888 520922 39944
rect 520978 39888 520983 39944
rect 518758 39886 520983 39888
rect 116945 39538 117011 39541
rect 116945 39536 119140 39538
rect 116945 39480 116950 39536
rect 117006 39480 119140 39536
rect 116945 39478 119140 39480
rect 116945 39475 117011 39478
rect 518758 39236 518818 39886
rect 520917 39883 520983 39886
rect 520917 39810 520983 39813
rect 523200 39810 524400 39840
rect 520917 39808 524400 39810
rect 520917 39752 520922 39808
rect 520978 39752 524400 39808
rect 520917 39750 524400 39752
rect 520917 39747 520983 39750
rect 523200 39720 524400 39750
rect 521101 38314 521167 38317
rect 523200 38314 524400 38344
rect 521101 38312 524400 38314
rect 521101 38256 521106 38312
rect 521162 38256 524400 38312
rect 521101 38254 524400 38256
rect 521101 38251 521167 38254
rect 523200 38224 524400 38254
rect 520917 37906 520983 37909
rect 518788 37904 520983 37906
rect 518788 37848 520922 37904
rect 520978 37848 520983 37904
rect 518788 37846 520983 37848
rect 520917 37843 520983 37846
rect 116853 37634 116919 37637
rect 116853 37632 119140 37634
rect 116853 37576 116858 37632
rect 116914 37576 119140 37632
rect 116853 37574 119140 37576
rect 116853 37571 116919 37574
rect 521101 37226 521167 37229
rect 518758 37224 521167 37226
rect 518758 37168 521106 37224
rect 521162 37168 521167 37224
rect 518758 37166 521167 37168
rect 518758 36516 518818 37166
rect 521101 37163 521167 37166
rect 521561 36818 521627 36821
rect 523200 36818 524400 36848
rect 521561 36816 524400 36818
rect 521561 36760 521566 36816
rect 521622 36760 524400 36816
rect 521561 36758 524400 36760
rect 521561 36755 521627 36758
rect 523200 36728 524400 36758
rect 521561 36002 521627 36005
rect 521561 36000 521670 36002
rect 521561 35944 521566 36000
rect 521622 35944 521670 36000
rect 521561 35939 521670 35944
rect 521610 35866 521670 35939
rect 518758 35806 521670 35866
rect 110321 34642 110387 34645
rect 119110 34642 119170 35700
rect 518758 35156 518818 35806
rect 520917 35322 520983 35325
rect 523200 35322 524400 35352
rect 520917 35320 524400 35322
rect 520917 35264 520922 35320
rect 520978 35264 524400 35320
rect 520917 35262 524400 35264
rect 520917 35259 520983 35262
rect 523200 35232 524400 35262
rect 110321 34640 119170 34642
rect 110321 34584 110326 34640
rect 110382 34584 119170 34640
rect 110321 34582 119170 34584
rect 110321 34579 110387 34582
rect 520917 34506 520983 34509
rect 518758 34504 520983 34506
rect 518758 34448 520922 34504
rect 520978 34448 520983 34504
rect 518758 34446 520983 34448
rect 117129 33826 117195 33829
rect 117129 33824 119140 33826
rect 117129 33768 117134 33824
rect 117190 33768 119140 33824
rect 518758 33796 518818 34446
rect 520917 34443 520983 34446
rect 521101 33826 521167 33829
rect 523200 33826 524400 33856
rect 521101 33824 524400 33826
rect 117129 33766 119140 33768
rect 521101 33768 521106 33824
rect 521162 33768 524400 33824
rect 521101 33766 524400 33768
rect 117129 33763 117195 33766
rect 521101 33763 521167 33766
rect 523200 33736 524400 33766
rect 521101 33146 521167 33149
rect 518758 33144 521167 33146
rect 518758 33088 521106 33144
rect 521162 33088 521167 33144
rect 518758 33086 521167 33088
rect 518758 32436 518818 33086
rect 521101 33083 521167 33086
rect 521101 32330 521167 32333
rect 523200 32330 524400 32360
rect 521101 32328 524400 32330
rect 521101 32272 521106 32328
rect 521162 32272 524400 32328
rect 521101 32270 524400 32272
rect 521101 32267 521167 32270
rect 523200 32240 524400 32270
rect 117037 31786 117103 31789
rect 117037 31784 119140 31786
rect 117037 31728 117042 31784
rect 117098 31728 119140 31784
rect 117037 31726 119140 31728
rect 117037 31723 117103 31726
rect 521101 31650 521167 31653
rect 518758 31648 521167 31650
rect 518758 31592 521106 31648
rect 521162 31592 521167 31648
rect 518758 31590 521167 31592
rect 518758 31076 518818 31590
rect 521101 31587 521167 31590
rect 523200 30834 524400 30864
rect 518850 30774 524400 30834
rect 114001 30426 114067 30429
rect 110860 30424 114067 30426
rect 110860 30368 114006 30424
rect 114062 30368 114067 30424
rect 110860 30366 114067 30368
rect 114001 30363 114067 30366
rect 518850 30290 518910 30774
rect 523200 30744 524400 30774
rect 518758 30230 518910 30290
rect 117221 29882 117287 29885
rect 117221 29880 119140 29882
rect 117221 29824 117226 29880
rect 117282 29824 119140 29880
rect 117221 29822 119140 29824
rect 117221 29819 117287 29822
rect 518758 29716 518818 30230
rect 520917 29338 520983 29341
rect 523200 29338 524400 29368
rect 520917 29336 524400 29338
rect 520917 29280 520922 29336
rect 520978 29280 524400 29336
rect 520917 29278 524400 29280
rect 520917 29275 520983 29278
rect 523200 29248 524400 29278
rect 520917 28386 520983 28389
rect 518788 28384 520983 28386
rect 518788 28328 520922 28384
rect 520978 28328 520983 28384
rect 518788 28326 520983 28328
rect 520917 28323 520983 28326
rect 116485 27978 116551 27981
rect 116485 27976 119140 27978
rect 116485 27920 116490 27976
rect 116546 27920 119140 27976
rect 116485 27918 119140 27920
rect 116485 27915 116551 27918
rect 523200 27842 524400 27872
rect 518850 27782 524400 27842
rect 518850 27570 518910 27782
rect 523200 27752 524400 27782
rect 518758 27510 518910 27570
rect 518758 26996 518818 27510
rect 523200 26346 524400 26376
rect 521610 26286 524400 26346
rect 521610 26210 521670 26286
rect 523200 26256 524400 26286
rect 518758 26150 521670 26210
rect 116301 26074 116367 26077
rect 116301 26072 119140 26074
rect 116301 26016 116306 26072
rect 116362 26016 119140 26072
rect 116301 26014 119140 26016
rect 116301 26011 116367 26014
rect 518758 25636 518818 26150
rect 521101 24850 521167 24853
rect 523200 24850 524400 24880
rect 521101 24848 524400 24850
rect 521101 24792 521106 24848
rect 521162 24792 524400 24848
rect 521101 24790 524400 24792
rect 521101 24787 521167 24790
rect 523200 24760 524400 24790
rect 116393 24170 116459 24173
rect 116393 24168 119140 24170
rect 116393 24112 116398 24168
rect 116454 24112 119140 24168
rect 116393 24110 119140 24112
rect 116393 24107 116459 24110
rect 518758 23626 518818 24276
rect 521101 23626 521167 23629
rect 518758 23624 521167 23626
rect 518758 23568 521106 23624
rect 521162 23568 521167 23624
rect 518758 23566 521167 23568
rect 521101 23563 521167 23566
rect 520365 23218 520431 23221
rect 523200 23218 524400 23248
rect 520365 23216 524400 23218
rect 520365 23160 520370 23216
rect 520426 23160 524400 23216
rect 520365 23158 524400 23160
rect 520365 23155 520431 23158
rect 523200 23128 524400 23158
rect 116209 22266 116275 22269
rect 518758 22266 518818 22916
rect 520365 22266 520431 22269
rect 116209 22264 119140 22266
rect 116209 22208 116214 22264
rect 116270 22208 119140 22264
rect 116209 22206 119140 22208
rect 518758 22264 520431 22266
rect 518758 22208 520370 22264
rect 520426 22208 520431 22264
rect 518758 22206 520431 22208
rect 116209 22203 116275 22206
rect 520365 22203 520431 22206
rect 520917 21722 520983 21725
rect 523200 21722 524400 21752
rect 520917 21720 524400 21722
rect 520917 21664 520922 21720
rect 520978 21664 524400 21720
rect 520917 21662 524400 21664
rect 520917 21659 520983 21662
rect 523200 21632 524400 21662
rect 518758 20906 518818 21556
rect 520917 20906 520983 20909
rect 518758 20904 520983 20906
rect 518758 20848 520922 20904
rect 520978 20848 520983 20904
rect 518758 20846 520983 20848
rect 520917 20843 520983 20846
rect 116025 20362 116091 20365
rect 116025 20360 119140 20362
rect 116025 20304 116030 20360
rect 116086 20304 119140 20360
rect 116025 20302 119140 20304
rect 116025 20299 116091 20302
rect 521101 20226 521167 20229
rect 523200 20226 524400 20256
rect 521101 20224 524400 20226
rect 518758 19546 518818 20196
rect 521101 20168 521106 20224
rect 521162 20168 524400 20224
rect 521101 20166 524400 20168
rect 521101 20163 521167 20166
rect 523200 20136 524400 20166
rect 521101 19546 521167 19549
rect 518758 19544 521167 19546
rect 518758 19488 521106 19544
rect 521162 19488 521167 19544
rect 518758 19486 521167 19488
rect 521101 19483 521167 19486
rect 113909 19002 113975 19005
rect 110860 19000 113975 19002
rect 110860 18944 113914 19000
rect 113970 18944 113975 19000
rect 110860 18942 113975 18944
rect 113909 18939 113975 18942
rect 116117 18458 116183 18461
rect 116117 18456 119140 18458
rect 116117 18400 116122 18456
rect 116178 18400 119140 18456
rect 116117 18398 119140 18400
rect 116117 18395 116183 18398
rect 518758 18186 518818 18836
rect 523200 18730 524400 18760
rect 521150 18670 524400 18730
rect 521150 18186 521210 18670
rect 523200 18640 524400 18670
rect 518758 18126 521210 18186
rect 518758 16826 518818 17476
rect 523200 17234 524400 17264
rect 521150 17174 524400 17234
rect 521150 16826 521210 17174
rect 523200 17144 524400 17174
rect 518758 16766 521210 16826
rect 115933 16418 115999 16421
rect 115933 16416 119140 16418
rect 115933 16360 115938 16416
rect 115994 16360 119140 16416
rect 115933 16358 119140 16360
rect 115933 16355 115999 16358
rect 518758 15466 518818 16116
rect 523200 15738 524400 15768
rect 521104 15678 524400 15738
rect 521104 15466 521164 15678
rect 523200 15648 524400 15678
rect 518758 15406 521164 15466
rect 116526 14452 116532 14516
rect 116596 14514 116602 14516
rect 116596 14454 119140 14514
rect 116596 14452 116602 14454
rect 518758 14106 518818 14756
rect 523200 14242 524400 14272
rect 521104 14182 524400 14242
rect 521104 14106 521164 14182
rect 523200 14152 524400 14182
rect 518758 14046 521164 14106
rect 518758 12746 518818 13396
rect 523200 12746 524400 12776
rect 518758 12686 524400 12746
rect 523200 12656 524400 12686
rect 116710 12548 116716 12612
rect 116780 12610 116786 12612
rect 116780 12550 119140 12610
rect 116780 12548 116786 12550
rect 518758 11386 518818 12036
rect 518758 11326 518910 11386
rect 518850 11250 518910 11326
rect 523200 11250 524400 11280
rect 518850 11190 524400 11250
rect 523200 11160 524400 11190
rect 116894 10644 116900 10708
rect 116964 10706 116970 10708
rect 116964 10646 119140 10706
rect 116964 10644 116970 10646
rect 518758 10026 518818 10676
rect 518758 9966 518910 10026
rect 518850 9754 518910 9966
rect 523200 9754 524400 9784
rect 518850 9694 524400 9754
rect 523200 9664 524400 9694
rect 521101 9346 521167 9349
rect 518788 9344 521167 9346
rect 518788 9288 521106 9344
rect 521162 9288 521167 9344
rect 518788 9286 521167 9288
rect 521101 9283 521167 9286
rect 117262 8740 117268 8804
rect 117332 8802 117338 8804
rect 117332 8742 119140 8802
rect 117332 8740 117338 8742
rect 110321 8258 110387 8261
rect 110505 8258 110571 8261
rect 110321 8256 110571 8258
rect 110321 8200 110326 8256
rect 110382 8200 110510 8256
rect 110566 8200 110571 8256
rect 110321 8198 110571 8200
rect 110321 8195 110387 8198
rect 110505 8195 110571 8198
rect 521101 8258 521167 8261
rect 523200 8258 524400 8288
rect 521101 8256 524400 8258
rect 521101 8200 521106 8256
rect 521162 8200 524400 8256
rect 521101 8198 524400 8200
rect 521101 8195 521167 8198
rect 523200 8168 524400 8198
rect 111057 7986 111123 7989
rect 116761 7986 116827 7989
rect 520365 7986 520431 7989
rect 111057 7984 116827 7986
rect 111057 7928 111062 7984
rect 111118 7928 116766 7984
rect 116822 7928 116827 7984
rect 111057 7926 116827 7928
rect 518788 7984 520431 7986
rect 518788 7928 520370 7984
rect 520426 7928 520431 7984
rect 518788 7926 520431 7928
rect 111057 7923 111123 7926
rect 116761 7923 116827 7926
rect 520365 7923 520431 7926
rect 113817 7714 113883 7717
rect 110860 7712 113883 7714
rect 110860 7656 113822 7712
rect 113878 7656 113883 7712
rect 110860 7654 113883 7656
rect 113817 7651 113883 7654
rect 117129 6898 117195 6901
rect 117129 6896 119140 6898
rect 117129 6840 117134 6896
rect 117190 6840 119140 6896
rect 117129 6838 119140 6840
rect 117129 6835 117195 6838
rect 520365 6762 520431 6765
rect 523200 6762 524400 6792
rect 520365 6760 524400 6762
rect 520365 6704 520370 6760
rect 520426 6704 524400 6760
rect 520365 6702 524400 6704
rect 520365 6699 520431 6702
rect 523200 6672 524400 6702
rect 521101 6626 521167 6629
rect 518788 6624 521167 6626
rect 518788 6568 521106 6624
rect 521162 6568 521167 6624
rect 518788 6566 521167 6568
rect 521101 6563 521167 6566
rect 110597 5674 110663 5677
rect 117037 5674 117103 5677
rect 110597 5672 117103 5674
rect 110597 5616 110602 5672
rect 110658 5616 117042 5672
rect 117098 5616 117103 5672
rect 110597 5614 117103 5616
rect 110597 5611 110663 5614
rect 117037 5611 117103 5614
rect 520917 5266 520983 5269
rect 518788 5264 520983 5266
rect 518788 5208 520922 5264
rect 520978 5208 520983 5264
rect 518788 5206 520983 5208
rect 520917 5203 520983 5206
rect 521101 5266 521167 5269
rect 523200 5266 524400 5296
rect 521101 5264 524400 5266
rect 521101 5208 521106 5264
rect 521162 5208 524400 5264
rect 521101 5206 524400 5208
rect 521101 5203 521167 5206
rect 523200 5176 524400 5206
rect 119110 4178 119170 4964
rect 110462 4118 119170 4178
rect 68326 3982 82830 4042
rect 55170 3438 59370 3498
rect 55170 3090 55230 3438
rect 45510 3030 55230 3090
rect 45510 2818 45570 3030
rect 32446 2758 45570 2818
rect 59310 2818 59370 3438
rect 59310 2758 63234 2818
rect 32446 2685 32506 2758
rect 32397 2680 32506 2685
rect 32397 2624 32402 2680
rect 32458 2624 32506 2680
rect 32397 2622 32506 2624
rect 36353 2682 36419 2685
rect 62389 2682 62455 2685
rect 36353 2680 62455 2682
rect 36353 2624 36358 2680
rect 36414 2624 62394 2680
rect 62450 2624 62455 2680
rect 36353 2622 62455 2624
rect 63174 2682 63234 2758
rect 68326 2685 68386 3982
rect 82770 3906 82830 3982
rect 88290 3982 109786 4042
rect 88290 3906 88350 3982
rect 109493 3906 109559 3909
rect 77342 3846 78690 3906
rect 82770 3846 88350 3906
rect 104390 3904 109559 3906
rect 104390 3848 109498 3904
rect 109554 3848 109559 3904
rect 104390 3846 109559 3848
rect 77342 3770 77402 3846
rect 77250 3710 77402 3770
rect 78630 3770 78690 3846
rect 78630 3710 82830 3770
rect 77250 2954 77310 3710
rect 82770 3498 82830 3710
rect 104390 3634 104450 3846
rect 109493 3843 109559 3846
rect 109726 3770 109786 3982
rect 110229 3906 110295 3909
rect 110462 3906 110522 4118
rect 521009 3906 521075 3909
rect 110229 3904 110522 3906
rect 110229 3848 110234 3904
rect 110290 3848 110522 3904
rect 110229 3846 110522 3848
rect 518788 3904 521075 3906
rect 518788 3848 521014 3904
rect 521070 3848 521075 3904
rect 518788 3846 521075 3848
rect 110229 3843 110295 3846
rect 521009 3843 521075 3846
rect 520917 3770 520983 3773
rect 523200 3770 524400 3800
rect 109726 3710 114570 3770
rect 109861 3634 109927 3637
rect 99054 3574 104450 3634
rect 106230 3632 109927 3634
rect 106230 3576 109866 3632
rect 109922 3576 109927 3632
rect 106230 3574 109927 3576
rect 114510 3634 114570 3710
rect 520917 3768 524400 3770
rect 520917 3712 520922 3768
rect 520978 3712 524400 3768
rect 520917 3710 524400 3712
rect 520917 3707 520983 3710
rect 523200 3680 524400 3710
rect 116301 3634 116367 3637
rect 114510 3632 116367 3634
rect 114510 3576 116306 3632
rect 116362 3576 116367 3632
rect 114510 3574 116367 3576
rect 82770 3438 88350 3498
rect 88290 3226 88350 3438
rect 88290 3166 89730 3226
rect 89670 3090 89730 3166
rect 68464 2894 77310 2954
rect 85530 3030 86970 3090
rect 89670 3030 91110 3090
rect 68464 2685 68524 2894
rect 85530 2818 85590 3030
rect 82770 2758 85590 2818
rect 64137 2682 64203 2685
rect 63174 2680 64203 2682
rect 63174 2624 64142 2680
rect 64198 2624 64203 2680
rect 63174 2622 64203 2624
rect 32397 2619 32463 2622
rect 36353 2619 36419 2622
rect 62389 2619 62455 2622
rect 64137 2619 64203 2622
rect 65333 2682 65399 2685
rect 68001 2682 68067 2685
rect 65333 2680 68067 2682
rect 65333 2624 65338 2680
rect 65394 2624 68006 2680
rect 68062 2624 68067 2680
rect 65333 2622 68067 2624
rect 65333 2619 65399 2622
rect 68001 2619 68067 2622
rect 68277 2680 68386 2685
rect 68277 2624 68282 2680
rect 68338 2624 68386 2680
rect 68277 2622 68386 2624
rect 68461 2680 68527 2685
rect 68461 2624 68466 2680
rect 68522 2624 68527 2680
rect 68277 2619 68343 2622
rect 68461 2619 68527 2624
rect 69381 2682 69447 2685
rect 75637 2682 75703 2685
rect 69381 2680 75703 2682
rect 69381 2624 69386 2680
rect 69442 2624 75642 2680
rect 75698 2624 75703 2680
rect 69381 2622 75703 2624
rect 69381 2619 69447 2622
rect 75637 2619 75703 2622
rect 77477 2682 77543 2685
rect 82770 2682 82830 2758
rect 77477 2680 82830 2682
rect 77477 2624 77482 2680
rect 77538 2624 82830 2680
rect 77477 2622 82830 2624
rect 85389 2682 85455 2685
rect 86677 2682 86743 2685
rect 85389 2680 86743 2682
rect 85389 2624 85394 2680
rect 85450 2624 86682 2680
rect 86738 2624 86743 2680
rect 85389 2622 86743 2624
rect 86910 2682 86970 3030
rect 91050 2954 91110 3030
rect 91050 2894 92490 2954
rect 91737 2682 91803 2685
rect 86910 2680 91803 2682
rect 86910 2624 91742 2680
rect 91798 2624 91803 2680
rect 86910 2622 91803 2624
rect 77477 2619 77543 2622
rect 85389 2619 85455 2622
rect 86677 2619 86743 2622
rect 91737 2619 91803 2622
rect 33041 2546 33107 2549
rect 91645 2546 91711 2549
rect 33041 2544 91711 2546
rect 33041 2488 33046 2544
rect 33102 2488 91650 2544
rect 91706 2488 91711 2544
rect 33041 2486 91711 2488
rect 92430 2546 92490 2894
rect 93025 2682 93091 2685
rect 98913 2682 98979 2685
rect 93025 2680 98979 2682
rect 93025 2624 93030 2680
rect 93086 2624 98918 2680
rect 98974 2624 98979 2680
rect 93025 2622 98979 2624
rect 93025 2619 93091 2622
rect 98913 2619 98979 2622
rect 95693 2546 95759 2549
rect 92430 2544 95759 2546
rect 92430 2488 95698 2544
rect 95754 2488 95759 2544
rect 92430 2486 95759 2488
rect 33041 2483 33107 2486
rect 91645 2483 91711 2486
rect 95693 2483 95759 2486
rect 96337 2546 96403 2549
rect 99054 2546 99114 3574
rect 106230 3498 106290 3574
rect 109861 3571 109927 3574
rect 116301 3571 116367 3574
rect 99422 3438 106290 3498
rect 109493 3498 109559 3501
rect 110229 3498 110295 3501
rect 109493 3496 110295 3498
rect 109493 3440 109498 3496
rect 109554 3440 110234 3496
rect 110290 3440 110295 3496
rect 109493 3438 110295 3440
rect 99189 2682 99255 2685
rect 99422 2682 99482 3438
rect 109493 3435 109559 3438
rect 110229 3435 110295 3438
rect 116945 3362 117011 3365
rect 103102 3360 117011 3362
rect 103102 3304 116950 3360
rect 117006 3304 117011 3360
rect 103102 3302 117011 3304
rect 103102 2954 103162 3302
rect 116945 3299 117011 3302
rect 110689 3226 110755 3229
rect 116669 3226 116735 3229
rect 102090 2894 103162 2954
rect 103286 3224 110755 3226
rect 103286 3168 110694 3224
rect 110750 3168 110755 3224
rect 103286 3166 110755 3168
rect 102090 2818 102150 2894
rect 99606 2758 102150 2818
rect 99606 2685 99666 2758
rect 99189 2680 99482 2682
rect 99189 2624 99194 2680
rect 99250 2624 99482 2680
rect 99189 2622 99482 2624
rect 99557 2680 99666 2685
rect 99557 2624 99562 2680
rect 99618 2624 99666 2680
rect 99557 2622 99666 2624
rect 99741 2682 99807 2685
rect 103286 2682 103346 3166
rect 110689 3163 110755 3166
rect 113038 3224 116735 3226
rect 113038 3168 116674 3224
rect 116730 3168 116735 3224
rect 113038 3166 116735 3168
rect 113038 3090 113098 3166
rect 116669 3163 116735 3166
rect 103470 3030 113098 3090
rect 116301 3090 116367 3093
rect 116301 3088 119140 3090
rect 116301 3032 116306 3088
rect 116362 3032 119140 3088
rect 116301 3030 119140 3032
rect 103470 2685 103530 3030
rect 116301 3027 116367 3030
rect 110137 2954 110203 2957
rect 111701 2954 111767 2957
rect 110137 2952 111767 2954
rect 110137 2896 110142 2952
rect 110198 2896 111706 2952
rect 111762 2896 111767 2952
rect 110137 2894 111767 2896
rect 110137 2891 110203 2894
rect 111701 2891 111767 2894
rect 109861 2818 109927 2821
rect 110597 2818 110663 2821
rect 109861 2816 110663 2818
rect 109861 2760 109866 2816
rect 109922 2760 110602 2816
rect 110658 2760 110663 2816
rect 109861 2758 110663 2760
rect 109861 2755 109927 2758
rect 110597 2755 110663 2758
rect 99741 2680 103346 2682
rect 99741 2624 99746 2680
rect 99802 2624 103346 2680
rect 99741 2622 103346 2624
rect 103421 2680 103530 2685
rect 116209 2682 116275 2685
rect 521101 2682 521167 2685
rect 103421 2624 103426 2680
rect 103482 2624 103530 2680
rect 103421 2622 103530 2624
rect 104022 2680 116275 2682
rect 104022 2624 116214 2680
rect 116270 2624 116275 2680
rect 104022 2622 116275 2624
rect 518788 2680 521167 2682
rect 518788 2624 521106 2680
rect 521162 2624 521167 2680
rect 518788 2622 521167 2624
rect 99189 2619 99255 2622
rect 99557 2619 99623 2622
rect 99741 2619 99807 2622
rect 103421 2619 103487 2622
rect 96337 2544 99114 2546
rect 96337 2488 96342 2544
rect 96398 2488 99114 2544
rect 96337 2486 99114 2488
rect 99833 2546 99899 2549
rect 104022 2546 104082 2622
rect 116209 2619 116275 2622
rect 521101 2619 521167 2622
rect 99833 2544 104082 2546
rect 99833 2488 99838 2544
rect 99894 2488 104082 2544
rect 99833 2486 104082 2488
rect 104157 2546 104223 2549
rect 116025 2546 116091 2549
rect 104157 2544 116091 2546
rect 104157 2488 104162 2544
rect 104218 2488 116030 2544
rect 116086 2488 116091 2544
rect 104157 2486 116091 2488
rect 96337 2483 96403 2486
rect 99833 2483 99899 2486
rect 104157 2483 104223 2486
rect 116025 2483 116091 2486
rect 29545 2410 29611 2413
rect 116117 2410 116183 2413
rect 29545 2408 116183 2410
rect 29545 2352 29550 2408
rect 29606 2352 116122 2408
rect 116178 2352 116183 2408
rect 29545 2350 116183 2352
rect 29545 2347 29611 2350
rect 116117 2347 116183 2350
rect 26049 2274 26115 2277
rect 115933 2274 115999 2277
rect 26049 2272 115999 2274
rect 26049 2216 26054 2272
rect 26110 2216 115938 2272
rect 115994 2216 115999 2272
rect 26049 2214 115999 2216
rect 26049 2211 26115 2214
rect 115933 2211 115999 2214
rect 521009 2274 521075 2277
rect 523200 2274 524400 2304
rect 521009 2272 524400 2274
rect 521009 2216 521014 2272
rect 521070 2216 524400 2272
rect 521009 2214 524400 2216
rect 521009 2211 521075 2214
rect 523200 2184 524400 2214
rect 22921 2138 22987 2141
rect 87965 2138 88031 2141
rect 22921 2136 88031 2138
rect 22921 2080 22926 2136
rect 22982 2080 87970 2136
rect 88026 2080 88031 2136
rect 22921 2078 88031 2080
rect 22921 2075 22987 2078
rect 87965 2075 88031 2078
rect 91645 2138 91711 2141
rect 104157 2138 104223 2141
rect 91645 2136 104223 2138
rect 91645 2080 91650 2136
rect 91706 2080 104162 2136
rect 104218 2080 104223 2136
rect 91645 2078 104223 2080
rect 91645 2075 91711 2078
rect 104157 2075 104223 2078
rect 104341 2138 104407 2141
rect 116526 2138 116532 2140
rect 104341 2136 116532 2138
rect 104341 2080 104346 2136
rect 104402 2080 116532 2136
rect 104341 2078 116532 2080
rect 104341 2075 104407 2078
rect 116526 2076 116532 2078
rect 116596 2076 116602 2140
rect 19609 2002 19675 2005
rect 116710 2002 116716 2004
rect 19609 2000 116716 2002
rect 19609 1944 19614 2000
rect 19670 1944 116716 2000
rect 19609 1942 116716 1944
rect 19609 1939 19675 1942
rect 116710 1940 116716 1942
rect 116780 1940 116786 2004
rect 15929 1866 15995 1869
rect 116894 1866 116900 1868
rect 15929 1864 116900 1866
rect 15929 1808 15934 1864
rect 15990 1808 116900 1864
rect 15929 1806 116900 1808
rect 15929 1803 15995 1806
rect 116894 1804 116900 1806
rect 116964 1804 116970 1868
rect 5993 1730 6059 1733
rect 109493 1730 109559 1733
rect 5993 1728 109559 1730
rect 5993 1672 5998 1728
rect 6054 1672 109498 1728
rect 109554 1672 109559 1728
rect 5993 1670 109559 1672
rect 5993 1667 6059 1670
rect 109493 1667 109559 1670
rect 12617 1594 12683 1597
rect 117262 1594 117268 1596
rect 12617 1592 117268 1594
rect 12617 1536 12622 1592
rect 12678 1536 117268 1592
rect 12617 1534 117268 1536
rect 12617 1531 12683 1534
rect 117262 1532 117268 1534
rect 117332 1532 117338 1596
rect 229277 1594 229343 1597
rect 293585 1594 293651 1597
rect 229277 1592 293651 1594
rect 229277 1536 229282 1592
rect 229338 1536 293590 1592
rect 293646 1536 293651 1592
rect 229277 1534 293651 1536
rect 229277 1531 229343 1534
rect 293585 1531 293651 1534
rect 9305 1458 9371 1461
rect 117129 1458 117195 1461
rect 9305 1456 117195 1458
rect 9305 1400 9310 1456
rect 9366 1400 117134 1456
rect 117190 1400 117195 1456
rect 9305 1398 117195 1400
rect 9305 1395 9371 1398
rect 117129 1395 117195 1398
rect 163773 1458 163839 1461
rect 243629 1458 243695 1461
rect 163773 1456 243695 1458
rect 163773 1400 163778 1456
rect 163834 1400 243634 1456
rect 243690 1400 243695 1456
rect 163773 1398 243695 1400
rect 163773 1395 163839 1398
rect 243629 1395 243695 1398
rect 360285 1458 360351 1461
rect 393589 1458 393655 1461
rect 360285 1456 393655 1458
rect 360285 1400 360290 1456
rect 360346 1400 393594 1456
rect 393650 1400 393655 1456
rect 360285 1398 393655 1400
rect 360285 1395 360351 1398
rect 393589 1395 393655 1398
rect 86677 1322 86743 1325
rect 103329 1322 103395 1325
rect 86677 1320 103395 1322
rect 86677 1264 86682 1320
rect 86738 1264 103334 1320
rect 103390 1264 103395 1320
rect 86677 1262 103395 1264
rect 86677 1259 86743 1262
rect 103329 1259 103395 1262
rect 108205 1322 108271 1325
rect 110229 1322 110295 1325
rect 108205 1320 110295 1322
rect 108205 1264 108210 1320
rect 108266 1264 110234 1320
rect 110290 1264 110295 1320
rect 108205 1262 110295 1264
rect 108205 1259 108271 1262
rect 110229 1259 110295 1262
rect 89253 1186 89319 1189
rect 98269 1186 98335 1189
rect 110137 1186 110203 1189
rect 89253 1184 92490 1186
rect 89253 1128 89258 1184
rect 89314 1128 92490 1184
rect 89253 1126 92490 1128
rect 89253 1123 89319 1126
rect 92430 1050 92490 1126
rect 98269 1184 110203 1186
rect 98269 1128 98274 1184
rect 98330 1128 110142 1184
rect 110198 1128 110203 1184
rect 98269 1126 110203 1128
rect 98269 1123 98335 1126
rect 110137 1123 110203 1126
rect 99833 1050 99899 1053
rect 92430 1048 99899 1050
rect 92430 992 99838 1048
rect 99894 992 99899 1048
rect 92430 990 99899 992
rect 99833 987 99899 990
rect 521101 778 521167 781
rect 523200 778 524400 808
rect 521101 776 524400 778
rect 521101 720 521106 776
rect 521162 720 524400 776
rect 521101 718 524400 720
rect 521101 715 521167 718
rect 523200 688 524400 718
<< via3 >>
rect 116532 14452 116596 14516
rect 116716 12548 116780 12612
rect 116900 10644 116964 10708
rect 117268 8740 117332 8804
rect 116532 2076 116596 2140
rect 116716 1940 116780 2004
rect 116900 1804 116964 1868
rect 117268 1532 117332 1596
<< metal4 >>
rect 1664 144454 1984 144496
rect 1664 144218 1706 144454
rect 1942 144218 1984 144454
rect 1664 144134 1984 144218
rect 1664 143898 1706 144134
rect 1942 143898 1984 144134
rect 1664 143856 1984 143898
rect 109956 144454 110276 144496
rect 109956 144218 109998 144454
rect 110234 144218 110276 144454
rect 109956 144134 110276 144218
rect 109956 143898 109998 144134
rect 110234 143898 110276 144134
rect 109956 143856 110276 143898
rect 119664 144454 119984 144496
rect 119664 144218 119706 144454
rect 119942 144218 119984 144454
rect 119664 144134 119984 144218
rect 119664 143898 119706 144134
rect 119942 143898 119984 144134
rect 119664 143856 119984 143898
rect 517940 144454 518260 144496
rect 517940 144218 517982 144454
rect 518218 144218 518260 144454
rect 517940 144134 518260 144218
rect 517940 143898 517982 144134
rect 518218 143898 518260 144134
rect 517940 143856 518260 143898
rect 1096 131454 1332 131496
rect 1096 131134 1332 131218
rect 1096 130856 1332 130898
rect 110616 131454 110936 131496
rect 110616 131218 110658 131454
rect 110894 131218 110936 131454
rect 110616 131134 110936 131218
rect 110616 130898 110658 131134
rect 110894 130898 110936 131134
rect 110616 130856 110936 130898
rect 119004 131454 119324 131496
rect 119004 131218 119046 131454
rect 119282 131218 119324 131454
rect 119004 131134 119324 131218
rect 119004 130898 119046 131134
rect 119282 130898 119324 131134
rect 119004 130856 119324 130898
rect 518600 131454 518920 131496
rect 518600 131218 518642 131454
rect 518878 131218 518920 131454
rect 518600 131134 518920 131218
rect 518600 130898 518642 131134
rect 518878 130898 518920 131134
rect 518600 130856 518920 130898
rect 1664 118454 1984 118496
rect 1664 118218 1706 118454
rect 1942 118218 1984 118454
rect 1664 118134 1984 118218
rect 1664 117898 1706 118134
rect 1942 117898 1984 118134
rect 1664 117856 1984 117898
rect 109956 118454 110276 118496
rect 109956 118218 109998 118454
rect 110234 118218 110276 118454
rect 109956 118134 110276 118218
rect 109956 117898 109998 118134
rect 110234 117898 110276 118134
rect 109956 117856 110276 117898
rect 119664 118454 119984 118496
rect 119664 118218 119706 118454
rect 119942 118218 119984 118454
rect 119664 118134 119984 118218
rect 119664 117898 119706 118134
rect 119942 117898 119984 118134
rect 119664 117856 119984 117898
rect 517940 118454 518260 118496
rect 517940 118218 517982 118454
rect 518218 118218 518260 118454
rect 517940 118134 518260 118218
rect 517940 117898 517982 118134
rect 518218 117898 518260 118134
rect 517940 117856 518260 117898
rect 1096 105454 1332 105496
rect 1096 105134 1332 105218
rect 1096 104856 1332 104898
rect 110616 105454 110936 105496
rect 110616 105218 110658 105454
rect 110894 105218 110936 105454
rect 110616 105134 110936 105218
rect 110616 104898 110658 105134
rect 110894 104898 110936 105134
rect 110616 104856 110936 104898
rect 119004 105454 119324 105496
rect 119004 105218 119046 105454
rect 119282 105218 119324 105454
rect 119004 105134 119324 105218
rect 119004 104898 119046 105134
rect 119282 104898 119324 105134
rect 119004 104856 119324 104898
rect 518600 105454 518920 105496
rect 518600 105218 518642 105454
rect 518878 105218 518920 105454
rect 518600 105134 518920 105218
rect 518600 104898 518642 105134
rect 518878 104898 518920 105134
rect 518600 104856 518920 104898
rect 1664 92454 1984 92496
rect 1664 92218 1706 92454
rect 1942 92218 1984 92454
rect 1664 92134 1984 92218
rect 1664 91898 1706 92134
rect 1942 91898 1984 92134
rect 1664 91856 1984 91898
rect 109956 92454 110276 92496
rect 109956 92218 109998 92454
rect 110234 92218 110276 92454
rect 109956 92134 110276 92218
rect 109956 91898 109998 92134
rect 110234 91898 110276 92134
rect 109956 91856 110276 91898
rect 119664 92454 119984 92496
rect 119664 92218 119706 92454
rect 119942 92218 119984 92454
rect 119664 92134 119984 92218
rect 119664 91898 119706 92134
rect 119942 91898 119984 92134
rect 119664 91856 119984 91898
rect 517940 92454 518260 92496
rect 517940 92218 517982 92454
rect 518218 92218 518260 92454
rect 517940 92134 518260 92218
rect 517940 91898 517982 92134
rect 518218 91898 518260 92134
rect 517940 91856 518260 91898
rect 1096 79454 1332 79496
rect 1096 79134 1332 79218
rect 1096 78856 1332 78898
rect 110616 79454 110936 79496
rect 110616 79218 110658 79454
rect 110894 79218 110936 79454
rect 110616 79134 110936 79218
rect 110616 78898 110658 79134
rect 110894 78898 110936 79134
rect 110616 78856 110936 78898
rect 119004 79454 119324 79496
rect 119004 79218 119046 79454
rect 119282 79218 119324 79454
rect 119004 79134 119324 79218
rect 119004 78898 119046 79134
rect 119282 78898 119324 79134
rect 119004 78856 119324 78898
rect 518600 79454 518920 79496
rect 518600 79218 518642 79454
rect 518878 79218 518920 79454
rect 518600 79134 518920 79218
rect 518600 78898 518642 79134
rect 518878 78898 518920 79134
rect 518600 78856 518920 78898
rect 1664 66454 1984 66496
rect 1664 66218 1706 66454
rect 1942 66218 1984 66454
rect 1664 66134 1984 66218
rect 1664 65898 1706 66134
rect 1942 65898 1984 66134
rect 1664 65856 1984 65898
rect 109956 66454 110276 66496
rect 109956 66218 109998 66454
rect 110234 66218 110276 66454
rect 109956 66134 110276 66218
rect 109956 65898 109998 66134
rect 110234 65898 110276 66134
rect 109956 65856 110276 65898
rect 119664 66454 119984 66496
rect 119664 66218 119706 66454
rect 119942 66218 119984 66454
rect 119664 66134 119984 66218
rect 119664 65898 119706 66134
rect 119942 65898 119984 66134
rect 119664 65856 119984 65898
rect 517940 66454 518260 66496
rect 517940 66218 517982 66454
rect 518218 66218 518260 66454
rect 517940 66134 518260 66218
rect 517940 65898 517982 66134
rect 518218 65898 518260 66134
rect 517940 65856 518260 65898
rect 1096 53454 1332 53496
rect 1096 53134 1332 53218
rect 1096 52856 1332 52898
rect 110616 53454 110936 53496
rect 110616 53218 110658 53454
rect 110894 53218 110936 53454
rect 110616 53134 110936 53218
rect 110616 52898 110658 53134
rect 110894 52898 110936 53134
rect 110616 52856 110936 52898
rect 119004 53454 119324 53496
rect 119004 53218 119046 53454
rect 119282 53218 119324 53454
rect 119004 53134 119324 53218
rect 119004 52898 119046 53134
rect 119282 52898 119324 53134
rect 119004 52856 119324 52898
rect 518600 53454 518920 53496
rect 518600 53218 518642 53454
rect 518878 53218 518920 53454
rect 518600 53134 518920 53218
rect 518600 52898 518642 53134
rect 518878 52898 518920 53134
rect 518600 52856 518920 52898
rect 1664 40454 1984 40496
rect 1664 40218 1706 40454
rect 1942 40218 1984 40454
rect 1664 40134 1984 40218
rect 1664 39898 1706 40134
rect 1942 39898 1984 40134
rect 1664 39856 1984 39898
rect 109956 40454 110276 40496
rect 109956 40218 109998 40454
rect 110234 40218 110276 40454
rect 109956 40134 110276 40218
rect 109956 39898 109998 40134
rect 110234 39898 110276 40134
rect 109956 39856 110276 39898
rect 119664 40454 119984 40496
rect 119664 40218 119706 40454
rect 119942 40218 119984 40454
rect 119664 40134 119984 40218
rect 119664 39898 119706 40134
rect 119942 39898 119984 40134
rect 119664 39856 119984 39898
rect 517940 40454 518260 40496
rect 517940 40218 517982 40454
rect 518218 40218 518260 40454
rect 517940 40134 518260 40218
rect 517940 39898 517982 40134
rect 518218 39898 518260 40134
rect 517940 39856 518260 39898
rect 1096 27454 1332 27496
rect 1096 27134 1332 27218
rect 1096 26856 1332 26898
rect 110616 27454 110936 27496
rect 110616 27218 110658 27454
rect 110894 27218 110936 27454
rect 110616 27134 110936 27218
rect 110616 26898 110658 27134
rect 110894 26898 110936 27134
rect 110616 26856 110936 26898
rect 119004 27454 119324 27496
rect 119004 27218 119046 27454
rect 119282 27218 119324 27454
rect 119004 27134 119324 27218
rect 119004 26898 119046 27134
rect 119282 26898 119324 27134
rect 119004 26856 119324 26898
rect 518600 27454 518920 27496
rect 518600 27218 518642 27454
rect 518878 27218 518920 27454
rect 518600 27134 518920 27218
rect 518600 26898 518642 27134
rect 518878 26898 518920 27134
rect 518600 26856 518920 26898
rect 116531 14516 116597 14517
rect 1664 14454 1984 14496
rect 1664 14218 1706 14454
rect 1942 14218 1984 14454
rect 1664 14134 1984 14218
rect 1664 13898 1706 14134
rect 1942 13898 1984 14134
rect 1664 13856 1984 13898
rect 109956 14454 110276 14496
rect 109956 14218 109998 14454
rect 110234 14218 110276 14454
rect 116531 14452 116532 14516
rect 116596 14452 116597 14516
rect 116531 14451 116597 14452
rect 119664 14454 119984 14496
rect 109956 14134 110276 14218
rect 109956 13898 109998 14134
rect 110234 13898 110276 14134
rect 109956 13856 110276 13898
rect 116534 2141 116594 14451
rect 119664 14218 119706 14454
rect 119942 14218 119984 14454
rect 119664 14134 119984 14218
rect 119664 13898 119706 14134
rect 119942 13898 119984 14134
rect 119664 13856 119984 13898
rect 517940 14454 518260 14496
rect 517940 14218 517982 14454
rect 518218 14218 518260 14454
rect 517940 14134 518260 14218
rect 517940 13898 517982 14134
rect 518218 13898 518260 14134
rect 517940 13856 518260 13898
rect 116715 12612 116781 12613
rect 116715 12548 116716 12612
rect 116780 12548 116781 12612
rect 116715 12547 116781 12548
rect 116531 2140 116597 2141
rect 116531 2076 116532 2140
rect 116596 2076 116597 2140
rect 116531 2075 116597 2076
rect 116718 2005 116778 12547
rect 116899 10708 116965 10709
rect 116899 10644 116900 10708
rect 116964 10644 116965 10708
rect 116899 10643 116965 10644
rect 116715 2004 116781 2005
rect 116715 1940 116716 2004
rect 116780 1940 116781 2004
rect 116715 1939 116781 1940
rect 116902 1869 116962 10643
rect 117267 8804 117333 8805
rect 117267 8740 117268 8804
rect 117332 8740 117333 8804
rect 117267 8739 117333 8740
rect 116899 1868 116965 1869
rect 116899 1804 116900 1868
rect 116964 1804 116965 1868
rect 116899 1803 116965 1804
rect 117270 1597 117330 8739
rect 117267 1596 117333 1597
rect 117267 1532 117268 1596
rect 117332 1532 117333 1596
rect 117267 1531 117333 1532
<< via4 >>
rect 1706 144218 1942 144454
rect 1706 143898 1942 144134
rect 109998 144218 110234 144454
rect 109998 143898 110234 144134
rect 119706 144218 119942 144454
rect 119706 143898 119942 144134
rect 517982 144218 518218 144454
rect 517982 143898 518218 144134
rect 1096 131218 1332 131454
rect 1096 130898 1332 131134
rect 110658 131218 110894 131454
rect 110658 130898 110894 131134
rect 119046 131218 119282 131454
rect 119046 130898 119282 131134
rect 518642 131218 518878 131454
rect 518642 130898 518878 131134
rect 1706 118218 1942 118454
rect 1706 117898 1942 118134
rect 109998 118218 110234 118454
rect 109998 117898 110234 118134
rect 119706 118218 119942 118454
rect 119706 117898 119942 118134
rect 517982 118218 518218 118454
rect 517982 117898 518218 118134
rect 1096 105218 1332 105454
rect 1096 104898 1332 105134
rect 110658 105218 110894 105454
rect 110658 104898 110894 105134
rect 119046 105218 119282 105454
rect 119046 104898 119282 105134
rect 518642 105218 518878 105454
rect 518642 104898 518878 105134
rect 1706 92218 1942 92454
rect 1706 91898 1942 92134
rect 109998 92218 110234 92454
rect 109998 91898 110234 92134
rect 119706 92218 119942 92454
rect 119706 91898 119942 92134
rect 517982 92218 518218 92454
rect 517982 91898 518218 92134
rect 1096 79218 1332 79454
rect 1096 78898 1332 79134
rect 110658 79218 110894 79454
rect 110658 78898 110894 79134
rect 119046 79218 119282 79454
rect 119046 78898 119282 79134
rect 518642 79218 518878 79454
rect 518642 78898 518878 79134
rect 1706 66218 1942 66454
rect 1706 65898 1942 66134
rect 109998 66218 110234 66454
rect 109998 65898 110234 66134
rect 119706 66218 119942 66454
rect 119706 65898 119942 66134
rect 517982 66218 518218 66454
rect 517982 65898 518218 66134
rect 1096 53218 1332 53454
rect 1096 52898 1332 53134
rect 110658 53218 110894 53454
rect 110658 52898 110894 53134
rect 119046 53218 119282 53454
rect 119046 52898 119282 53134
rect 518642 53218 518878 53454
rect 518642 52898 518878 53134
rect 1706 40218 1942 40454
rect 1706 39898 1942 40134
rect 109998 40218 110234 40454
rect 109998 39898 110234 40134
rect 119706 40218 119942 40454
rect 119706 39898 119942 40134
rect 517982 40218 518218 40454
rect 517982 39898 518218 40134
rect 1096 27218 1332 27454
rect 1096 26898 1332 27134
rect 110658 27218 110894 27454
rect 110658 26898 110894 27134
rect 119046 27218 119282 27454
rect 119046 26898 119282 27134
rect 518642 27218 518878 27454
rect 518642 26898 518878 27134
rect 1706 14218 1942 14454
rect 1706 13898 1942 14134
rect 109998 14218 110234 14454
rect 109998 13898 110234 14134
rect 119706 14218 119942 14454
rect 119706 13898 119942 14134
rect 517982 14218 518218 14454
rect 517982 13898 518218 14134
<< metal5 >>
rect 1104 156856 522836 157496
rect 1104 144454 2200 144496
rect 1104 144218 1706 144454
rect 1942 144218 2200 144454
rect 1104 144134 2200 144218
rect 1104 143898 1706 144134
rect 1942 143898 2200 144134
rect 1104 143856 2200 143898
rect 109800 144454 120200 144496
rect 109800 144218 109998 144454
rect 110234 144218 119706 144454
rect 119942 144218 120200 144454
rect 109800 144134 120200 144218
rect 109800 143898 109998 144134
rect 110234 143898 119706 144134
rect 119942 143898 120200 144134
rect 109800 143856 120200 143898
rect 517800 144454 522836 144496
rect 517800 144218 517982 144454
rect 518218 144218 522836 144454
rect 517800 144134 522836 144218
rect 517800 143898 517982 144134
rect 518218 143898 522836 144134
rect 517800 143856 522836 143898
rect 1072 131454 2200 131496
rect 1072 131218 1096 131454
rect 1332 131218 2200 131454
rect 1072 131134 2200 131218
rect 1072 130898 1096 131134
rect 1332 130898 2200 131134
rect 1072 130856 2200 130898
rect 109800 131454 120200 131496
rect 109800 131218 110658 131454
rect 110894 131218 119046 131454
rect 119282 131218 120200 131454
rect 109800 131134 120200 131218
rect 109800 130898 110658 131134
rect 110894 130898 119046 131134
rect 119282 130898 120200 131134
rect 109800 130856 120200 130898
rect 517800 131454 522836 131496
rect 517800 131218 518642 131454
rect 518878 131218 522836 131454
rect 517800 131134 522836 131218
rect 517800 130898 518642 131134
rect 518878 130898 522836 131134
rect 517800 130856 522836 130898
rect 1104 118454 2200 118496
rect 1104 118218 1706 118454
rect 1942 118218 2200 118454
rect 1104 118134 2200 118218
rect 1104 117898 1706 118134
rect 1942 117898 2200 118134
rect 1104 117856 2200 117898
rect 109800 118454 120200 118496
rect 109800 118218 109998 118454
rect 110234 118218 119706 118454
rect 119942 118218 120200 118454
rect 109800 118134 120200 118218
rect 109800 117898 109998 118134
rect 110234 117898 119706 118134
rect 119942 117898 120200 118134
rect 109800 117856 120200 117898
rect 517800 118454 522836 118496
rect 517800 118218 517982 118454
rect 518218 118218 522836 118454
rect 517800 118134 522836 118218
rect 517800 117898 517982 118134
rect 518218 117898 522836 118134
rect 517800 117856 522836 117898
rect 1072 105454 2200 105496
rect 1072 105218 1096 105454
rect 1332 105218 2200 105454
rect 1072 105134 2200 105218
rect 1072 104898 1096 105134
rect 1332 104898 2200 105134
rect 1072 104856 2200 104898
rect 109800 105454 120200 105496
rect 109800 105218 110658 105454
rect 110894 105218 119046 105454
rect 119282 105218 120200 105454
rect 109800 105134 120200 105218
rect 109800 104898 110658 105134
rect 110894 104898 119046 105134
rect 119282 104898 120200 105134
rect 109800 104856 120200 104898
rect 517800 105454 522836 105496
rect 517800 105218 518642 105454
rect 518878 105218 522836 105454
rect 517800 105134 522836 105218
rect 517800 104898 518642 105134
rect 518878 104898 522836 105134
rect 517800 104856 522836 104898
rect 1104 92454 2200 92496
rect 1104 92218 1706 92454
rect 1942 92218 2200 92454
rect 1104 92134 2200 92218
rect 1104 91898 1706 92134
rect 1942 91898 2200 92134
rect 1104 91856 2200 91898
rect 109800 92454 120200 92496
rect 109800 92218 109998 92454
rect 110234 92218 119706 92454
rect 119942 92218 120200 92454
rect 109800 92134 120200 92218
rect 109800 91898 109998 92134
rect 110234 91898 119706 92134
rect 119942 91898 120200 92134
rect 109800 91856 120200 91898
rect 517800 92454 522836 92496
rect 517800 92218 517982 92454
rect 518218 92218 522836 92454
rect 517800 92134 522836 92218
rect 517800 91898 517982 92134
rect 518218 91898 522836 92134
rect 517800 91856 522836 91898
rect 1072 79454 2200 79496
rect 1072 79218 1096 79454
rect 1332 79218 2200 79454
rect 1072 79134 2200 79218
rect 1072 78898 1096 79134
rect 1332 78898 2200 79134
rect 1072 78856 2200 78898
rect 109800 79454 120200 79496
rect 109800 79218 110658 79454
rect 110894 79218 119046 79454
rect 119282 79218 120200 79454
rect 109800 79134 120200 79218
rect 109800 78898 110658 79134
rect 110894 78898 119046 79134
rect 119282 78898 120200 79134
rect 109800 78856 120200 78898
rect 517800 79454 522836 79496
rect 517800 79218 518642 79454
rect 518878 79218 522836 79454
rect 517800 79134 522836 79218
rect 517800 78898 518642 79134
rect 518878 78898 522836 79134
rect 517800 78856 522836 78898
rect 1104 66454 2200 66496
rect 1104 66218 1706 66454
rect 1942 66218 2200 66454
rect 1104 66134 2200 66218
rect 1104 65898 1706 66134
rect 1942 65898 2200 66134
rect 1104 65856 2200 65898
rect 109800 66454 120200 66496
rect 109800 66218 109998 66454
rect 110234 66218 119706 66454
rect 119942 66218 120200 66454
rect 109800 66134 120200 66218
rect 109800 65898 109998 66134
rect 110234 65898 119706 66134
rect 119942 65898 120200 66134
rect 109800 65856 120200 65898
rect 517800 66454 522836 66496
rect 517800 66218 517982 66454
rect 518218 66218 522836 66454
rect 517800 66134 522836 66218
rect 517800 65898 517982 66134
rect 518218 65898 522836 66134
rect 517800 65856 522836 65898
rect 1072 53454 2200 53496
rect 1072 53218 1096 53454
rect 1332 53218 2200 53454
rect 1072 53134 2200 53218
rect 1072 52898 1096 53134
rect 1332 52898 2200 53134
rect 1072 52856 2200 52898
rect 109800 53454 120200 53496
rect 109800 53218 110658 53454
rect 110894 53218 119046 53454
rect 119282 53218 120200 53454
rect 109800 53134 120200 53218
rect 109800 52898 110658 53134
rect 110894 52898 119046 53134
rect 119282 52898 120200 53134
rect 109800 52856 120200 52898
rect 517800 53454 522836 53496
rect 517800 53218 518642 53454
rect 518878 53218 522836 53454
rect 517800 53134 522836 53218
rect 517800 52898 518642 53134
rect 518878 52898 522836 53134
rect 517800 52856 522836 52898
rect 1104 40454 2200 40496
rect 1104 40218 1706 40454
rect 1942 40218 2200 40454
rect 1104 40134 2200 40218
rect 1104 39898 1706 40134
rect 1942 39898 2200 40134
rect 1104 39856 2200 39898
rect 109800 40454 120200 40496
rect 109800 40218 109998 40454
rect 110234 40218 119706 40454
rect 119942 40218 120200 40454
rect 109800 40134 120200 40218
rect 109800 39898 109998 40134
rect 110234 39898 119706 40134
rect 119942 39898 120200 40134
rect 109800 39856 120200 39898
rect 517800 40454 522836 40496
rect 517800 40218 517982 40454
rect 518218 40218 522836 40454
rect 517800 40134 522836 40218
rect 517800 39898 517982 40134
rect 518218 39898 522836 40134
rect 517800 39856 522836 39898
rect 1072 27454 2200 27496
rect 1072 27218 1096 27454
rect 1332 27218 2200 27454
rect 1072 27134 2200 27218
rect 1072 26898 1096 27134
rect 1332 26898 2200 27134
rect 1072 26856 2200 26898
rect 109800 27454 120200 27496
rect 109800 27218 110658 27454
rect 110894 27218 119046 27454
rect 119282 27218 120200 27454
rect 109800 27134 120200 27218
rect 109800 26898 110658 27134
rect 110894 26898 119046 27134
rect 119282 26898 120200 27134
rect 109800 26856 120200 26898
rect 517800 27454 522836 27496
rect 517800 27218 518642 27454
rect 518878 27218 522836 27454
rect 517800 27134 522836 27218
rect 517800 26898 518642 27134
rect 518878 26898 522836 27134
rect 517800 26856 522836 26898
rect 1104 14454 2200 14496
rect 1104 14218 1706 14454
rect 1942 14218 2200 14454
rect 1104 14134 2200 14218
rect 1104 13898 1706 14134
rect 1942 13898 2200 14134
rect 1104 13856 2200 13898
rect 109800 14454 120200 14496
rect 109800 14218 109998 14454
rect 110234 14218 119706 14454
rect 119942 14218 120200 14454
rect 109800 14134 120200 14218
rect 109800 13898 109998 14134
rect 110234 13898 119706 14134
rect 119942 13898 120200 14134
rect 109800 13856 120200 13898
rect 517800 14454 522836 14496
rect 517800 14218 517982 14454
rect 518218 14218 522836 14454
rect 517800 14134 522836 14218
rect 517800 13898 517982 14134
rect 518218 13898 522836 14134
rect 517800 13856 522836 13898
use mgmt_core  core
timestamp 1638728696
transform 1 0 119000 0 1 2000
box 0 0 400000 148000
use DFFRAM  DFFRAM_0
timestamp 1638728696
transform 1 0 1000 0 1 2000
box 4 0 110000 148000
<< labels >>
rlabel metal5 s 1104 26856 2200 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 26856 120200 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 26856 522836 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 52856 2200 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 52856 120200 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 52856 522836 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 78856 2200 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 78856 120200 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 78856 522836 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 104856 2200 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 104856 120200 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 104856 522836 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 130856 2200 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 130856 120200 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 130856 522836 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 156856 522836 157496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 13856 2200 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 13856 120200 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 13856 522836 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 39856 2200 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 39856 120200 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 39856 522836 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 65856 2200 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 65856 120200 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 65856 522836 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 91856 2200 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 91856 120200 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 91856 522836 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 117856 2200 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 117856 120200 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 117856 522836 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 143856 2200 144496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 143856 120200 144496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 143856 522836 144496 6 VPWR
port 1 nsew power input
rlabel metal2 s 294786 -400 294842 800 6 core_clk
port 2 nsew signal input
rlabel metal2 s 98274 -400 98330 800 6 core_rstn
port 3 nsew signal input
rlabel metal3 s 523200 63792 524400 63912 6 debug_in
port 4 nsew signal input
rlabel metal3 s 523200 65288 524400 65408 6 debug_mode
port 5 nsew signal tristate
rlabel metal3 s 523200 66784 524400 66904 6 debug_oeb
port 6 nsew signal tristate
rlabel metal3 s 523200 68280 524400 68400 6 debug_out
port 7 nsew signal tristate
rlabel metal3 s 523200 145120 524400 145240 6 flash_clk
port 8 nsew signal tristate
rlabel metal3 s 523200 143624 524400 143744 6 flash_csb
port 9 nsew signal tristate
rlabel metal3 s 523200 146616 524400 146736 6 flash_io0_di
port 10 nsew signal input
rlabel metal3 s 523200 148112 524400 148232 6 flash_io0_do
port 11 nsew signal tristate
rlabel metal3 s 523200 149608 524400 149728 6 flash_io0_oeb
port 12 nsew signal tristate
rlabel metal3 s 523200 151104 524400 151224 6 flash_io1_di
port 13 nsew signal input
rlabel metal3 s 523200 152600 524400 152720 6 flash_io1_do
port 14 nsew signal tristate
rlabel metal3 s 523200 154096 524400 154216 6 flash_io1_oeb
port 15 nsew signal tristate
rlabel metal3 s 523200 155592 524400 155712 6 flash_io2_di
port 16 nsew signal input
rlabel metal3 s 523200 157088 524400 157208 6 flash_io2_do
port 17 nsew signal tristate
rlabel metal3 s 523200 158584 524400 158704 6 flash_io2_oeb
port 18 nsew signal tristate
rlabel metal3 s 523200 160080 524400 160200 6 flash_io3_di
port 19 nsew signal input
rlabel metal3 s 523200 161576 524400 161696 6 flash_io3_do
port 20 nsew signal tristate
rlabel metal3 s 523200 163072 524400 163192 6 flash_io3_oeb
port 21 nsew signal tristate
rlabel metal2 s 32770 -400 32826 800 6 gpio_in_pad
port 22 nsew signal input
rlabel metal2 s 163778 -400 163834 800 6 gpio_inenb_pad
port 23 nsew signal tristate
rlabel metal2 s 229282 -400 229338 800 6 gpio_mode0_pad
port 24 nsew signal tristate
rlabel metal2 s 360290 -400 360346 800 6 gpio_mode1_pad
port 25 nsew signal tristate
rlabel metal2 s 425794 -400 425850 800 6 gpio_out_pad
port 26 nsew signal tristate
rlabel metal2 s 491298 -400 491354 800 6 gpio_outenb_pad
port 27 nsew signal tristate
rlabel metal3 s 523200 90856 524400 90976 6 hk_ack_i
port 28 nsew signal input
rlabel metal3 s 523200 93848 524400 93968 6 hk_cyc_o
port 29 nsew signal tristate
rlabel metal3 s 523200 95480 524400 95600 6 hk_dat_i[0]
port 30 nsew signal input
rlabel metal3 s 523200 110440 524400 110560 6 hk_dat_i[10]
port 31 nsew signal input
rlabel metal3 s 523200 111936 524400 112056 6 hk_dat_i[11]
port 32 nsew signal input
rlabel metal3 s 523200 113432 524400 113552 6 hk_dat_i[12]
port 33 nsew signal input
rlabel metal3 s 523200 114928 524400 115048 6 hk_dat_i[13]
port 34 nsew signal input
rlabel metal3 s 523200 116424 524400 116544 6 hk_dat_i[14]
port 35 nsew signal input
rlabel metal3 s 523200 118056 524400 118176 6 hk_dat_i[15]
port 36 nsew signal input
rlabel metal3 s 523200 119552 524400 119672 6 hk_dat_i[16]
port 37 nsew signal input
rlabel metal3 s 523200 121048 524400 121168 6 hk_dat_i[17]
port 38 nsew signal input
rlabel metal3 s 523200 122544 524400 122664 6 hk_dat_i[18]
port 39 nsew signal input
rlabel metal3 s 523200 124040 524400 124160 6 hk_dat_i[19]
port 40 nsew signal input
rlabel metal3 s 523200 96976 524400 97096 6 hk_dat_i[1]
port 41 nsew signal input
rlabel metal3 s 523200 125536 524400 125656 6 hk_dat_i[20]
port 42 nsew signal input
rlabel metal3 s 523200 127032 524400 127152 6 hk_dat_i[21]
port 43 nsew signal input
rlabel metal3 s 523200 128528 524400 128648 6 hk_dat_i[22]
port 44 nsew signal input
rlabel metal3 s 523200 130024 524400 130144 6 hk_dat_i[23]
port 45 nsew signal input
rlabel metal3 s 523200 131520 524400 131640 6 hk_dat_i[24]
port 46 nsew signal input
rlabel metal3 s 523200 133016 524400 133136 6 hk_dat_i[25]
port 47 nsew signal input
rlabel metal3 s 523200 134512 524400 134632 6 hk_dat_i[26]
port 48 nsew signal input
rlabel metal3 s 523200 136008 524400 136128 6 hk_dat_i[27]
port 49 nsew signal input
rlabel metal3 s 523200 137504 524400 137624 6 hk_dat_i[28]
port 50 nsew signal input
rlabel metal3 s 523200 139000 524400 139120 6 hk_dat_i[29]
port 51 nsew signal input
rlabel metal3 s 523200 98472 524400 98592 6 hk_dat_i[2]
port 52 nsew signal input
rlabel metal3 s 523200 140496 524400 140616 6 hk_dat_i[30]
port 53 nsew signal input
rlabel metal3 s 523200 142128 524400 142248 6 hk_dat_i[31]
port 54 nsew signal input
rlabel metal3 s 523200 99968 524400 100088 6 hk_dat_i[3]
port 55 nsew signal input
rlabel metal3 s 523200 101464 524400 101584 6 hk_dat_i[4]
port 56 nsew signal input
rlabel metal3 s 523200 102960 524400 103080 6 hk_dat_i[5]
port 57 nsew signal input
rlabel metal3 s 523200 104456 524400 104576 6 hk_dat_i[6]
port 58 nsew signal input
rlabel metal3 s 523200 105952 524400 106072 6 hk_dat_i[7]
port 59 nsew signal input
rlabel metal3 s 523200 107448 524400 107568 6 hk_dat_i[8]
port 60 nsew signal input
rlabel metal3 s 523200 108944 524400 109064 6 hk_dat_i[9]
port 61 nsew signal input
rlabel metal3 s 523200 92352 524400 92472 6 hk_stb_o
port 62 nsew signal tristate
rlabel metal2 s 521842 163200 521898 164400 6 irq[0]
port 63 nsew signal input
rlabel metal2 s 522670 163200 522726 164400 6 irq[1]
port 64 nsew signal input
rlabel metal2 s 523498 163200 523554 164400 6 irq[2]
port 65 nsew signal input
rlabel metal3 s 523200 74400 524400 74520 6 irq[3]
port 66 nsew signal input
rlabel metal3 s 523200 72904 524400 73024 6 irq[4]
port 67 nsew signal input
rlabel metal3 s 523200 71408 524400 71528 6 irq[5]
port 68 nsew signal input
rlabel metal2 s 386 163200 442 164400 6 la_iena[0]
port 69 nsew signal tristate
rlabel metal2 s 336830 163200 336886 164400 6 la_iena[100]
port 70 nsew signal tristate
rlabel metal2 s 340142 163200 340198 164400 6 la_iena[101]
port 71 nsew signal tristate
rlabel metal2 s 343546 163200 343602 164400 6 la_iena[102]
port 72 nsew signal tristate
rlabel metal2 s 346858 163200 346914 164400 6 la_iena[103]
port 73 nsew signal tristate
rlabel metal2 s 350262 163200 350318 164400 6 la_iena[104]
port 74 nsew signal tristate
rlabel metal2 s 353666 163200 353722 164400 6 la_iena[105]
port 75 nsew signal tristate
rlabel metal2 s 356978 163200 357034 164400 6 la_iena[106]
port 76 nsew signal tristate
rlabel metal2 s 360382 163200 360438 164400 6 la_iena[107]
port 77 nsew signal tristate
rlabel metal2 s 363694 163200 363750 164400 6 la_iena[108]
port 78 nsew signal tristate
rlabel metal2 s 367098 163200 367154 164400 6 la_iena[109]
port 79 nsew signal tristate
rlabel metal2 s 33966 163200 34022 164400 6 la_iena[10]
port 80 nsew signal tristate
rlabel metal2 s 370410 163200 370466 164400 6 la_iena[110]
port 81 nsew signal tristate
rlabel metal2 s 373814 163200 373870 164400 6 la_iena[111]
port 82 nsew signal tristate
rlabel metal2 s 377218 163200 377274 164400 6 la_iena[112]
port 83 nsew signal tristate
rlabel metal2 s 380530 163200 380586 164400 6 la_iena[113]
port 84 nsew signal tristate
rlabel metal2 s 383934 163200 383990 164400 6 la_iena[114]
port 85 nsew signal tristate
rlabel metal2 s 387246 163200 387302 164400 6 la_iena[115]
port 86 nsew signal tristate
rlabel metal2 s 390650 163200 390706 164400 6 la_iena[116]
port 87 nsew signal tristate
rlabel metal2 s 393962 163200 394018 164400 6 la_iena[117]
port 88 nsew signal tristate
rlabel metal2 s 397366 163200 397422 164400 6 la_iena[118]
port 89 nsew signal tristate
rlabel metal2 s 400770 163200 400826 164400 6 la_iena[119]
port 90 nsew signal tristate
rlabel metal2 s 37370 163200 37426 164400 6 la_iena[11]
port 91 nsew signal tristate
rlabel metal2 s 404082 163200 404138 164400 6 la_iena[120]
port 92 nsew signal tristate
rlabel metal2 s 407486 163200 407542 164400 6 la_iena[121]
port 93 nsew signal tristate
rlabel metal2 s 410798 163200 410854 164400 6 la_iena[122]
port 94 nsew signal tristate
rlabel metal2 s 414202 163200 414258 164400 6 la_iena[123]
port 95 nsew signal tristate
rlabel metal2 s 417514 163200 417570 164400 6 la_iena[124]
port 96 nsew signal tristate
rlabel metal2 s 420918 163200 420974 164400 6 la_iena[125]
port 97 nsew signal tristate
rlabel metal2 s 424322 163200 424378 164400 6 la_iena[126]
port 98 nsew signal tristate
rlabel metal2 s 427634 163200 427690 164400 6 la_iena[127]
port 99 nsew signal tristate
rlabel metal2 s 40682 163200 40738 164400 6 la_iena[12]
port 100 nsew signal tristate
rlabel metal2 s 44086 163200 44142 164400 6 la_iena[13]
port 101 nsew signal tristate
rlabel metal2 s 47490 163200 47546 164400 6 la_iena[14]
port 102 nsew signal tristate
rlabel metal2 s 50802 163200 50858 164400 6 la_iena[15]
port 103 nsew signal tristate
rlabel metal2 s 54206 163200 54262 164400 6 la_iena[16]
port 104 nsew signal tristate
rlabel metal2 s 57518 163200 57574 164400 6 la_iena[17]
port 105 nsew signal tristate
rlabel metal2 s 60922 163200 60978 164400 6 la_iena[18]
port 106 nsew signal tristate
rlabel metal2 s 64234 163200 64290 164400 6 la_iena[19]
port 107 nsew signal tristate
rlabel metal2 s 3698 163200 3754 164400 6 la_iena[1]
port 108 nsew signal tristate
rlabel metal2 s 67638 163200 67694 164400 6 la_iena[20]
port 109 nsew signal tristate
rlabel metal2 s 71042 163200 71098 164400 6 la_iena[21]
port 110 nsew signal tristate
rlabel metal2 s 74354 163200 74410 164400 6 la_iena[22]
port 111 nsew signal tristate
rlabel metal2 s 77758 163200 77814 164400 6 la_iena[23]
port 112 nsew signal tristate
rlabel metal2 s 81070 163200 81126 164400 6 la_iena[24]
port 113 nsew signal tristate
rlabel metal2 s 84474 163200 84530 164400 6 la_iena[25]
port 114 nsew signal tristate
rlabel metal2 s 87786 163200 87842 164400 6 la_iena[26]
port 115 nsew signal tristate
rlabel metal2 s 91190 163200 91246 164400 6 la_iena[27]
port 116 nsew signal tristate
rlabel metal2 s 94594 163200 94650 164400 6 la_iena[28]
port 117 nsew signal tristate
rlabel metal2 s 97906 163200 97962 164400 6 la_iena[29]
port 118 nsew signal tristate
rlabel metal2 s 7102 163200 7158 164400 6 la_iena[2]
port 119 nsew signal tristate
rlabel metal2 s 101310 163200 101366 164400 6 la_iena[30]
port 120 nsew signal tristate
rlabel metal2 s 104622 163200 104678 164400 6 la_iena[31]
port 121 nsew signal tristate
rlabel metal2 s 108026 163200 108082 164400 6 la_iena[32]
port 122 nsew signal tristate
rlabel metal2 s 111338 163200 111394 164400 6 la_iena[33]
port 123 nsew signal tristate
rlabel metal2 s 114742 163200 114798 164400 6 la_iena[34]
port 124 nsew signal tristate
rlabel metal2 s 118146 163200 118202 164400 6 la_iena[35]
port 125 nsew signal tristate
rlabel metal2 s 121458 163200 121514 164400 6 la_iena[36]
port 126 nsew signal tristate
rlabel metal2 s 124862 163200 124918 164400 6 la_iena[37]
port 127 nsew signal tristate
rlabel metal2 s 128174 163200 128230 164400 6 la_iena[38]
port 128 nsew signal tristate
rlabel metal2 s 131578 163200 131634 164400 6 la_iena[39]
port 129 nsew signal tristate
rlabel metal2 s 10414 163200 10470 164400 6 la_iena[3]
port 130 nsew signal tristate
rlabel metal2 s 134890 163200 134946 164400 6 la_iena[40]
port 131 nsew signal tristate
rlabel metal2 s 138294 163200 138350 164400 6 la_iena[41]
port 132 nsew signal tristate
rlabel metal2 s 141698 163200 141754 164400 6 la_iena[42]
port 133 nsew signal tristate
rlabel metal2 s 145010 163200 145066 164400 6 la_iena[43]
port 134 nsew signal tristate
rlabel metal2 s 148414 163200 148470 164400 6 la_iena[44]
port 135 nsew signal tristate
rlabel metal2 s 151726 163200 151782 164400 6 la_iena[45]
port 136 nsew signal tristate
rlabel metal2 s 155130 163200 155186 164400 6 la_iena[46]
port 137 nsew signal tristate
rlabel metal2 s 158442 163200 158498 164400 6 la_iena[47]
port 138 nsew signal tristate
rlabel metal2 s 161846 163200 161902 164400 6 la_iena[48]
port 139 nsew signal tristate
rlabel metal2 s 165250 163200 165306 164400 6 la_iena[49]
port 140 nsew signal tristate
rlabel metal2 s 13818 163200 13874 164400 6 la_iena[4]
port 141 nsew signal tristate
rlabel metal2 s 168562 163200 168618 164400 6 la_iena[50]
port 142 nsew signal tristate
rlabel metal2 s 171966 163200 172022 164400 6 la_iena[51]
port 143 nsew signal tristate
rlabel metal2 s 175278 163200 175334 164400 6 la_iena[52]
port 144 nsew signal tristate
rlabel metal2 s 178682 163200 178738 164400 6 la_iena[53]
port 145 nsew signal tristate
rlabel metal2 s 181994 163200 182050 164400 6 la_iena[54]
port 146 nsew signal tristate
rlabel metal2 s 185398 163200 185454 164400 6 la_iena[55]
port 147 nsew signal tristate
rlabel metal2 s 188802 163200 188858 164400 6 la_iena[56]
port 148 nsew signal tristate
rlabel metal2 s 192114 163200 192170 164400 6 la_iena[57]
port 149 nsew signal tristate
rlabel metal2 s 195518 163200 195574 164400 6 la_iena[58]
port 150 nsew signal tristate
rlabel metal2 s 198830 163200 198886 164400 6 la_iena[59]
port 151 nsew signal tristate
rlabel metal2 s 17130 163200 17186 164400 6 la_iena[5]
port 152 nsew signal tristate
rlabel metal2 s 202234 163200 202290 164400 6 la_iena[60]
port 153 nsew signal tristate
rlabel metal2 s 205546 163200 205602 164400 6 la_iena[61]
port 154 nsew signal tristate
rlabel metal2 s 208950 163200 209006 164400 6 la_iena[62]
port 155 nsew signal tristate
rlabel metal2 s 212354 163200 212410 164400 6 la_iena[63]
port 156 nsew signal tristate
rlabel metal2 s 215666 163200 215722 164400 6 la_iena[64]
port 157 nsew signal tristate
rlabel metal2 s 219070 163200 219126 164400 6 la_iena[65]
port 158 nsew signal tristate
rlabel metal2 s 222382 163200 222438 164400 6 la_iena[66]
port 159 nsew signal tristate
rlabel metal2 s 225786 163200 225842 164400 6 la_iena[67]
port 160 nsew signal tristate
rlabel metal2 s 229098 163200 229154 164400 6 la_iena[68]
port 161 nsew signal tristate
rlabel metal2 s 232502 163200 232558 164400 6 la_iena[69]
port 162 nsew signal tristate
rlabel metal2 s 20534 163200 20590 164400 6 la_iena[6]
port 163 nsew signal tristate
rlabel metal2 s 235906 163200 235962 164400 6 la_iena[70]
port 164 nsew signal tristate
rlabel metal2 s 239218 163200 239274 164400 6 la_iena[71]
port 165 nsew signal tristate
rlabel metal2 s 242622 163200 242678 164400 6 la_iena[72]
port 166 nsew signal tristate
rlabel metal2 s 245934 163200 245990 164400 6 la_iena[73]
port 167 nsew signal tristate
rlabel metal2 s 249338 163200 249394 164400 6 la_iena[74]
port 168 nsew signal tristate
rlabel metal2 s 252650 163200 252706 164400 6 la_iena[75]
port 169 nsew signal tristate
rlabel metal2 s 256054 163200 256110 164400 6 la_iena[76]
port 170 nsew signal tristate
rlabel metal2 s 259458 163200 259514 164400 6 la_iena[77]
port 171 nsew signal tristate
rlabel metal2 s 262770 163200 262826 164400 6 la_iena[78]
port 172 nsew signal tristate
rlabel metal2 s 266174 163200 266230 164400 6 la_iena[79]
port 173 nsew signal tristate
rlabel metal2 s 23938 163200 23994 164400 6 la_iena[7]
port 174 nsew signal tristate
rlabel metal2 s 269486 163200 269542 164400 6 la_iena[80]
port 175 nsew signal tristate
rlabel metal2 s 272890 163200 272946 164400 6 la_iena[81]
port 176 nsew signal tristate
rlabel metal2 s 276202 163200 276258 164400 6 la_iena[82]
port 177 nsew signal tristate
rlabel metal2 s 279606 163200 279662 164400 6 la_iena[83]
port 178 nsew signal tristate
rlabel metal2 s 283010 163200 283066 164400 6 la_iena[84]
port 179 nsew signal tristate
rlabel metal2 s 286322 163200 286378 164400 6 la_iena[85]
port 180 nsew signal tristate
rlabel metal2 s 289726 163200 289782 164400 6 la_iena[86]
port 181 nsew signal tristate
rlabel metal2 s 293038 163200 293094 164400 6 la_iena[87]
port 182 nsew signal tristate
rlabel metal2 s 296442 163200 296498 164400 6 la_iena[88]
port 183 nsew signal tristate
rlabel metal2 s 299754 163200 299810 164400 6 la_iena[89]
port 184 nsew signal tristate
rlabel metal2 s 27250 163200 27306 164400 6 la_iena[8]
port 185 nsew signal tristate
rlabel metal2 s 303158 163200 303214 164400 6 la_iena[90]
port 186 nsew signal tristate
rlabel metal2 s 306562 163200 306618 164400 6 la_iena[91]
port 187 nsew signal tristate
rlabel metal2 s 309874 163200 309930 164400 6 la_iena[92]
port 188 nsew signal tristate
rlabel metal2 s 313278 163200 313334 164400 6 la_iena[93]
port 189 nsew signal tristate
rlabel metal2 s 316590 163200 316646 164400 6 la_iena[94]
port 190 nsew signal tristate
rlabel metal2 s 319994 163200 320050 164400 6 la_iena[95]
port 191 nsew signal tristate
rlabel metal2 s 323306 163200 323362 164400 6 la_iena[96]
port 192 nsew signal tristate
rlabel metal2 s 326710 163200 326766 164400 6 la_iena[97]
port 193 nsew signal tristate
rlabel metal2 s 330114 163200 330170 164400 6 la_iena[98]
port 194 nsew signal tristate
rlabel metal2 s 333426 163200 333482 164400 6 la_iena[99]
port 195 nsew signal tristate
rlabel metal2 s 30654 163200 30710 164400 6 la_iena[9]
port 196 nsew signal tristate
rlabel metal2 s 1214 163200 1270 164400 6 la_input[0]
port 197 nsew signal input
rlabel metal2 s 337658 163200 337714 164400 6 la_input[100]
port 198 nsew signal input
rlabel metal2 s 340970 163200 341026 164400 6 la_input[101]
port 199 nsew signal input
rlabel metal2 s 344374 163200 344430 164400 6 la_input[102]
port 200 nsew signal input
rlabel metal2 s 347778 163200 347834 164400 6 la_input[103]
port 201 nsew signal input
rlabel metal2 s 351090 163200 351146 164400 6 la_input[104]
port 202 nsew signal input
rlabel metal2 s 354494 163200 354550 164400 6 la_input[105]
port 203 nsew signal input
rlabel metal2 s 357806 163200 357862 164400 6 la_input[106]
port 204 nsew signal input
rlabel metal2 s 361210 163200 361266 164400 6 la_input[107]
port 205 nsew signal input
rlabel metal2 s 364522 163200 364578 164400 6 la_input[108]
port 206 nsew signal input
rlabel metal2 s 367926 163200 367982 164400 6 la_input[109]
port 207 nsew signal input
rlabel metal2 s 34794 163200 34850 164400 6 la_input[10]
port 208 nsew signal input
rlabel metal2 s 371330 163200 371386 164400 6 la_input[110]
port 209 nsew signal input
rlabel metal2 s 374642 163200 374698 164400 6 la_input[111]
port 210 nsew signal input
rlabel metal2 s 378046 163200 378102 164400 6 la_input[112]
port 211 nsew signal input
rlabel metal2 s 381358 163200 381414 164400 6 la_input[113]
port 212 nsew signal input
rlabel metal2 s 384762 163200 384818 164400 6 la_input[114]
port 213 nsew signal input
rlabel metal2 s 388074 163200 388130 164400 6 la_input[115]
port 214 nsew signal input
rlabel metal2 s 391478 163200 391534 164400 6 la_input[116]
port 215 nsew signal input
rlabel metal2 s 394882 163200 394938 164400 6 la_input[117]
port 216 nsew signal input
rlabel metal2 s 398194 163200 398250 164400 6 la_input[118]
port 217 nsew signal input
rlabel metal2 s 401598 163200 401654 164400 6 la_input[119]
port 218 nsew signal input
rlabel metal2 s 38198 163200 38254 164400 6 la_input[11]
port 219 nsew signal input
rlabel metal2 s 404910 163200 404966 164400 6 la_input[120]
port 220 nsew signal input
rlabel metal2 s 408314 163200 408370 164400 6 la_input[121]
port 221 nsew signal input
rlabel metal2 s 411626 163200 411682 164400 6 la_input[122]
port 222 nsew signal input
rlabel metal2 s 415030 163200 415086 164400 6 la_input[123]
port 223 nsew signal input
rlabel metal2 s 418434 163200 418490 164400 6 la_input[124]
port 224 nsew signal input
rlabel metal2 s 421746 163200 421802 164400 6 la_input[125]
port 225 nsew signal input
rlabel metal2 s 425150 163200 425206 164400 6 la_input[126]
port 226 nsew signal input
rlabel metal2 s 428462 163200 428518 164400 6 la_input[127]
port 227 nsew signal input
rlabel metal2 s 41602 163200 41658 164400 6 la_input[12]
port 228 nsew signal input
rlabel metal2 s 44914 163200 44970 164400 6 la_input[13]
port 229 nsew signal input
rlabel metal2 s 48318 163200 48374 164400 6 la_input[14]
port 230 nsew signal input
rlabel metal2 s 51630 163200 51686 164400 6 la_input[15]
port 231 nsew signal input
rlabel metal2 s 55034 163200 55090 164400 6 la_input[16]
port 232 nsew signal input
rlabel metal2 s 58346 163200 58402 164400 6 la_input[17]
port 233 nsew signal input
rlabel metal2 s 61750 163200 61806 164400 6 la_input[18]
port 234 nsew signal input
rlabel metal2 s 65154 163200 65210 164400 6 la_input[19]
port 235 nsew signal input
rlabel metal2 s 4526 163200 4582 164400 6 la_input[1]
port 236 nsew signal input
rlabel metal2 s 68466 163200 68522 164400 6 la_input[20]
port 237 nsew signal input
rlabel metal2 s 71870 163200 71926 164400 6 la_input[21]
port 238 nsew signal input
rlabel metal2 s 75182 163200 75238 164400 6 la_input[22]
port 239 nsew signal input
rlabel metal2 s 78586 163200 78642 164400 6 la_input[23]
port 240 nsew signal input
rlabel metal2 s 81898 163200 81954 164400 6 la_input[24]
port 241 nsew signal input
rlabel metal2 s 85302 163200 85358 164400 6 la_input[25]
port 242 nsew signal input
rlabel metal2 s 88706 163200 88762 164400 6 la_input[26]
port 243 nsew signal input
rlabel metal2 s 92018 163200 92074 164400 6 la_input[27]
port 244 nsew signal input
rlabel metal2 s 95422 163200 95478 164400 6 la_input[28]
port 245 nsew signal input
rlabel metal2 s 98734 163200 98790 164400 6 la_input[29]
port 246 nsew signal input
rlabel metal2 s 7930 163200 7986 164400 6 la_input[2]
port 247 nsew signal input
rlabel metal2 s 102138 163200 102194 164400 6 la_input[30]
port 248 nsew signal input
rlabel metal2 s 105450 163200 105506 164400 6 la_input[31]
port 249 nsew signal input
rlabel metal2 s 108854 163200 108910 164400 6 la_input[32]
port 250 nsew signal input
rlabel metal2 s 112258 163200 112314 164400 6 la_input[33]
port 251 nsew signal input
rlabel metal2 s 115570 163200 115626 164400 6 la_input[34]
port 252 nsew signal input
rlabel metal2 s 118974 163200 119030 164400 6 la_input[35]
port 253 nsew signal input
rlabel metal2 s 122286 163200 122342 164400 6 la_input[36]
port 254 nsew signal input
rlabel metal2 s 125690 163200 125746 164400 6 la_input[37]
port 255 nsew signal input
rlabel metal2 s 129002 163200 129058 164400 6 la_input[38]
port 256 nsew signal input
rlabel metal2 s 132406 163200 132462 164400 6 la_input[39]
port 257 nsew signal input
rlabel metal2 s 11242 163200 11298 164400 6 la_input[3]
port 258 nsew signal input
rlabel metal2 s 135810 163200 135866 164400 6 la_input[40]
port 259 nsew signal input
rlabel metal2 s 139122 163200 139178 164400 6 la_input[41]
port 260 nsew signal input
rlabel metal2 s 142526 163200 142582 164400 6 la_input[42]
port 261 nsew signal input
rlabel metal2 s 145838 163200 145894 164400 6 la_input[43]
port 262 nsew signal input
rlabel metal2 s 149242 163200 149298 164400 6 la_input[44]
port 263 nsew signal input
rlabel metal2 s 152554 163200 152610 164400 6 la_input[45]
port 264 nsew signal input
rlabel metal2 s 155958 163200 156014 164400 6 la_input[46]
port 265 nsew signal input
rlabel metal2 s 159362 163200 159418 164400 6 la_input[47]
port 266 nsew signal input
rlabel metal2 s 162674 163200 162730 164400 6 la_input[48]
port 267 nsew signal input
rlabel metal2 s 166078 163200 166134 164400 6 la_input[49]
port 268 nsew signal input
rlabel metal2 s 14646 163200 14702 164400 6 la_input[4]
port 269 nsew signal input
rlabel metal2 s 169390 163200 169446 164400 6 la_input[50]
port 270 nsew signal input
rlabel metal2 s 172794 163200 172850 164400 6 la_input[51]
port 271 nsew signal input
rlabel metal2 s 176106 163200 176162 164400 6 la_input[52]
port 272 nsew signal input
rlabel metal2 s 179510 163200 179566 164400 6 la_input[53]
port 273 nsew signal input
rlabel metal2 s 182914 163200 182970 164400 6 la_input[54]
port 274 nsew signal input
rlabel metal2 s 186226 163200 186282 164400 6 la_input[55]
port 275 nsew signal input
rlabel metal2 s 189630 163200 189686 164400 6 la_input[56]
port 276 nsew signal input
rlabel metal2 s 192942 163200 192998 164400 6 la_input[57]
port 277 nsew signal input
rlabel metal2 s 196346 163200 196402 164400 6 la_input[58]
port 278 nsew signal input
rlabel metal2 s 199658 163200 199714 164400 6 la_input[59]
port 279 nsew signal input
rlabel metal2 s 18050 163200 18106 164400 6 la_input[5]
port 280 nsew signal input
rlabel metal2 s 203062 163200 203118 164400 6 la_input[60]
port 281 nsew signal input
rlabel metal2 s 206466 163200 206522 164400 6 la_input[61]
port 282 nsew signal input
rlabel metal2 s 209778 163200 209834 164400 6 la_input[62]
port 283 nsew signal input
rlabel metal2 s 213182 163200 213238 164400 6 la_input[63]
port 284 nsew signal input
rlabel metal2 s 216494 163200 216550 164400 6 la_input[64]
port 285 nsew signal input
rlabel metal2 s 219898 163200 219954 164400 6 la_input[65]
port 286 nsew signal input
rlabel metal2 s 223210 163200 223266 164400 6 la_input[66]
port 287 nsew signal input
rlabel metal2 s 226614 163200 226670 164400 6 la_input[67]
port 288 nsew signal input
rlabel metal2 s 230018 163200 230074 164400 6 la_input[68]
port 289 nsew signal input
rlabel metal2 s 233330 163200 233386 164400 6 la_input[69]
port 290 nsew signal input
rlabel metal2 s 21362 163200 21418 164400 6 la_input[6]
port 291 nsew signal input
rlabel metal2 s 236734 163200 236790 164400 6 la_input[70]
port 292 nsew signal input
rlabel metal2 s 240046 163200 240102 164400 6 la_input[71]
port 293 nsew signal input
rlabel metal2 s 243450 163200 243506 164400 6 la_input[72]
port 294 nsew signal input
rlabel metal2 s 246762 163200 246818 164400 6 la_input[73]
port 295 nsew signal input
rlabel metal2 s 250166 163200 250222 164400 6 la_input[74]
port 296 nsew signal input
rlabel metal2 s 253570 163200 253626 164400 6 la_input[75]
port 297 nsew signal input
rlabel metal2 s 256882 163200 256938 164400 6 la_input[76]
port 298 nsew signal input
rlabel metal2 s 260286 163200 260342 164400 6 la_input[77]
port 299 nsew signal input
rlabel metal2 s 263598 163200 263654 164400 6 la_input[78]
port 300 nsew signal input
rlabel metal2 s 267002 163200 267058 164400 6 la_input[79]
port 301 nsew signal input
rlabel metal2 s 24766 163200 24822 164400 6 la_input[7]
port 302 nsew signal input
rlabel metal2 s 270314 163200 270370 164400 6 la_input[80]
port 303 nsew signal input
rlabel metal2 s 273718 163200 273774 164400 6 la_input[81]
port 304 nsew signal input
rlabel metal2 s 277122 163200 277178 164400 6 la_input[82]
port 305 nsew signal input
rlabel metal2 s 280434 163200 280490 164400 6 la_input[83]
port 306 nsew signal input
rlabel metal2 s 283838 163200 283894 164400 6 la_input[84]
port 307 nsew signal input
rlabel metal2 s 287150 163200 287206 164400 6 la_input[85]
port 308 nsew signal input
rlabel metal2 s 290554 163200 290610 164400 6 la_input[86]
port 309 nsew signal input
rlabel metal2 s 293866 163200 293922 164400 6 la_input[87]
port 310 nsew signal input
rlabel metal2 s 297270 163200 297326 164400 6 la_input[88]
port 311 nsew signal input
rlabel metal2 s 300674 163200 300730 164400 6 la_input[89]
port 312 nsew signal input
rlabel metal2 s 28078 163200 28134 164400 6 la_input[8]
port 313 nsew signal input
rlabel metal2 s 303986 163200 304042 164400 6 la_input[90]
port 314 nsew signal input
rlabel metal2 s 307390 163200 307446 164400 6 la_input[91]
port 315 nsew signal input
rlabel metal2 s 310702 163200 310758 164400 6 la_input[92]
port 316 nsew signal input
rlabel metal2 s 314106 163200 314162 164400 6 la_input[93]
port 317 nsew signal input
rlabel metal2 s 317418 163200 317474 164400 6 la_input[94]
port 318 nsew signal input
rlabel metal2 s 320822 163200 320878 164400 6 la_input[95]
port 319 nsew signal input
rlabel metal2 s 324226 163200 324282 164400 6 la_input[96]
port 320 nsew signal input
rlabel metal2 s 327538 163200 327594 164400 6 la_input[97]
port 321 nsew signal input
rlabel metal2 s 330942 163200 330998 164400 6 la_input[98]
port 322 nsew signal input
rlabel metal2 s 334254 163200 334310 164400 6 la_input[99]
port 323 nsew signal input
rlabel metal2 s 31482 163200 31538 164400 6 la_input[9]
port 324 nsew signal input
rlabel metal2 s 2042 163200 2098 164400 6 la_oenb[0]
port 325 nsew signal tristate
rlabel metal2 s 338486 163200 338542 164400 6 la_oenb[100]
port 326 nsew signal tristate
rlabel metal2 s 341890 163200 341946 164400 6 la_oenb[101]
port 327 nsew signal tristate
rlabel metal2 s 345202 163200 345258 164400 6 la_oenb[102]
port 328 nsew signal tristate
rlabel metal2 s 348606 163200 348662 164400 6 la_oenb[103]
port 329 nsew signal tristate
rlabel metal2 s 351918 163200 351974 164400 6 la_oenb[104]
port 330 nsew signal tristate
rlabel metal2 s 355322 163200 355378 164400 6 la_oenb[105]
port 331 nsew signal tristate
rlabel metal2 s 358634 163200 358690 164400 6 la_oenb[106]
port 332 nsew signal tristate
rlabel metal2 s 362038 163200 362094 164400 6 la_oenb[107]
port 333 nsew signal tristate
rlabel metal2 s 365442 163200 365498 164400 6 la_oenb[108]
port 334 nsew signal tristate
rlabel metal2 s 368754 163200 368810 164400 6 la_oenb[109]
port 335 nsew signal tristate
rlabel metal2 s 35714 163200 35770 164400 6 la_oenb[10]
port 336 nsew signal tristate
rlabel metal2 s 372158 163200 372214 164400 6 la_oenb[110]
port 337 nsew signal tristate
rlabel metal2 s 375470 163200 375526 164400 6 la_oenb[111]
port 338 nsew signal tristate
rlabel metal2 s 378874 163200 378930 164400 6 la_oenb[112]
port 339 nsew signal tristate
rlabel metal2 s 382186 163200 382242 164400 6 la_oenb[113]
port 340 nsew signal tristate
rlabel metal2 s 385590 163200 385646 164400 6 la_oenb[114]
port 341 nsew signal tristate
rlabel metal2 s 388994 163200 389050 164400 6 la_oenb[115]
port 342 nsew signal tristate
rlabel metal2 s 392306 163200 392362 164400 6 la_oenb[116]
port 343 nsew signal tristate
rlabel metal2 s 395710 163200 395766 164400 6 la_oenb[117]
port 344 nsew signal tristate
rlabel metal2 s 399022 163200 399078 164400 6 la_oenb[118]
port 345 nsew signal tristate
rlabel metal2 s 402426 163200 402482 164400 6 la_oenb[119]
port 346 nsew signal tristate
rlabel metal2 s 39026 163200 39082 164400 6 la_oenb[11]
port 347 nsew signal tristate
rlabel metal2 s 405738 163200 405794 164400 6 la_oenb[120]
port 348 nsew signal tristate
rlabel metal2 s 409142 163200 409198 164400 6 la_oenb[121]
port 349 nsew signal tristate
rlabel metal2 s 412546 163200 412602 164400 6 la_oenb[122]
port 350 nsew signal tristate
rlabel metal2 s 415858 163200 415914 164400 6 la_oenb[123]
port 351 nsew signal tristate
rlabel metal2 s 419262 163200 419318 164400 6 la_oenb[124]
port 352 nsew signal tristate
rlabel metal2 s 422574 163200 422630 164400 6 la_oenb[125]
port 353 nsew signal tristate
rlabel metal2 s 425978 163200 426034 164400 6 la_oenb[126]
port 354 nsew signal tristate
rlabel metal2 s 429290 163200 429346 164400 6 la_oenb[127]
port 355 nsew signal tristate
rlabel metal2 s 42430 163200 42486 164400 6 la_oenb[12]
port 356 nsew signal tristate
rlabel metal2 s 45742 163200 45798 164400 6 la_oenb[13]
port 357 nsew signal tristate
rlabel metal2 s 49146 163200 49202 164400 6 la_oenb[14]
port 358 nsew signal tristate
rlabel metal2 s 52458 163200 52514 164400 6 la_oenb[15]
port 359 nsew signal tristate
rlabel metal2 s 55862 163200 55918 164400 6 la_oenb[16]
port 360 nsew signal tristate
rlabel metal2 s 59266 163200 59322 164400 6 la_oenb[17]
port 361 nsew signal tristate
rlabel metal2 s 62578 163200 62634 164400 6 la_oenb[18]
port 362 nsew signal tristate
rlabel metal2 s 65982 163200 66038 164400 6 la_oenb[19]
port 363 nsew signal tristate
rlabel metal2 s 5354 163200 5410 164400 6 la_oenb[1]
port 364 nsew signal tristate
rlabel metal2 s 69294 163200 69350 164400 6 la_oenb[20]
port 365 nsew signal tristate
rlabel metal2 s 72698 163200 72754 164400 6 la_oenb[21]
port 366 nsew signal tristate
rlabel metal2 s 76010 163200 76066 164400 6 la_oenb[22]
port 367 nsew signal tristate
rlabel metal2 s 79414 163200 79470 164400 6 la_oenb[23]
port 368 nsew signal tristate
rlabel metal2 s 82818 163200 82874 164400 6 la_oenb[24]
port 369 nsew signal tristate
rlabel metal2 s 86130 163200 86186 164400 6 la_oenb[25]
port 370 nsew signal tristate
rlabel metal2 s 89534 163200 89590 164400 6 la_oenb[26]
port 371 nsew signal tristate
rlabel metal2 s 92846 163200 92902 164400 6 la_oenb[27]
port 372 nsew signal tristate
rlabel metal2 s 96250 163200 96306 164400 6 la_oenb[28]
port 373 nsew signal tristate
rlabel metal2 s 99562 163200 99618 164400 6 la_oenb[29]
port 374 nsew signal tristate
rlabel metal2 s 8758 163200 8814 164400 6 la_oenb[2]
port 375 nsew signal tristate
rlabel metal2 s 102966 163200 103022 164400 6 la_oenb[30]
port 376 nsew signal tristate
rlabel metal2 s 106370 163200 106426 164400 6 la_oenb[31]
port 377 nsew signal tristate
rlabel metal2 s 109682 163200 109738 164400 6 la_oenb[32]
port 378 nsew signal tristate
rlabel metal2 s 113086 163200 113142 164400 6 la_oenb[33]
port 379 nsew signal tristate
rlabel metal2 s 116398 163200 116454 164400 6 la_oenb[34]
port 380 nsew signal tristate
rlabel metal2 s 119802 163200 119858 164400 6 la_oenb[35]
port 381 nsew signal tristate
rlabel metal2 s 123114 163200 123170 164400 6 la_oenb[36]
port 382 nsew signal tristate
rlabel metal2 s 126518 163200 126574 164400 6 la_oenb[37]
port 383 nsew signal tristate
rlabel metal2 s 129922 163200 129978 164400 6 la_oenb[38]
port 384 nsew signal tristate
rlabel metal2 s 133234 163200 133290 164400 6 la_oenb[39]
port 385 nsew signal tristate
rlabel metal2 s 12162 163200 12218 164400 6 la_oenb[3]
port 386 nsew signal tristate
rlabel metal2 s 136638 163200 136694 164400 6 la_oenb[40]
port 387 nsew signal tristate
rlabel metal2 s 139950 163200 140006 164400 6 la_oenb[41]
port 388 nsew signal tristate
rlabel metal2 s 143354 163200 143410 164400 6 la_oenb[42]
port 389 nsew signal tristate
rlabel metal2 s 146666 163200 146722 164400 6 la_oenb[43]
port 390 nsew signal tristate
rlabel metal2 s 150070 163200 150126 164400 6 la_oenb[44]
port 391 nsew signal tristate
rlabel metal2 s 153474 163200 153530 164400 6 la_oenb[45]
port 392 nsew signal tristate
rlabel metal2 s 156786 163200 156842 164400 6 la_oenb[46]
port 393 nsew signal tristate
rlabel metal2 s 160190 163200 160246 164400 6 la_oenb[47]
port 394 nsew signal tristate
rlabel metal2 s 163502 163200 163558 164400 6 la_oenb[48]
port 395 nsew signal tristate
rlabel metal2 s 166906 163200 166962 164400 6 la_oenb[49]
port 396 nsew signal tristate
rlabel metal2 s 15474 163200 15530 164400 6 la_oenb[4]
port 397 nsew signal tristate
rlabel metal2 s 170218 163200 170274 164400 6 la_oenb[50]
port 398 nsew signal tristate
rlabel metal2 s 173622 163200 173678 164400 6 la_oenb[51]
port 399 nsew signal tristate
rlabel metal2 s 177026 163200 177082 164400 6 la_oenb[52]
port 400 nsew signal tristate
rlabel metal2 s 180338 163200 180394 164400 6 la_oenb[53]
port 401 nsew signal tristate
rlabel metal2 s 183742 163200 183798 164400 6 la_oenb[54]
port 402 nsew signal tristate
rlabel metal2 s 187054 163200 187110 164400 6 la_oenb[55]
port 403 nsew signal tristate
rlabel metal2 s 190458 163200 190514 164400 6 la_oenb[56]
port 404 nsew signal tristate
rlabel metal2 s 193770 163200 193826 164400 6 la_oenb[57]
port 405 nsew signal tristate
rlabel metal2 s 197174 163200 197230 164400 6 la_oenb[58]
port 406 nsew signal tristate
rlabel metal2 s 200578 163200 200634 164400 6 la_oenb[59]
port 407 nsew signal tristate
rlabel metal2 s 18878 163200 18934 164400 6 la_oenb[5]
port 408 nsew signal tristate
rlabel metal2 s 203890 163200 203946 164400 6 la_oenb[60]
port 409 nsew signal tristate
rlabel metal2 s 207294 163200 207350 164400 6 la_oenb[61]
port 410 nsew signal tristate
rlabel metal2 s 210606 163200 210662 164400 6 la_oenb[62]
port 411 nsew signal tristate
rlabel metal2 s 214010 163200 214066 164400 6 la_oenb[63]
port 412 nsew signal tristate
rlabel metal2 s 217322 163200 217378 164400 6 la_oenb[64]
port 413 nsew signal tristate
rlabel metal2 s 220726 163200 220782 164400 6 la_oenb[65]
port 414 nsew signal tristate
rlabel metal2 s 224130 163200 224186 164400 6 la_oenb[66]
port 415 nsew signal tristate
rlabel metal2 s 227442 163200 227498 164400 6 la_oenb[67]
port 416 nsew signal tristate
rlabel metal2 s 230846 163200 230902 164400 6 la_oenb[68]
port 417 nsew signal tristate
rlabel metal2 s 234158 163200 234214 164400 6 la_oenb[69]
port 418 nsew signal tristate
rlabel metal2 s 22190 163200 22246 164400 6 la_oenb[6]
port 419 nsew signal tristate
rlabel metal2 s 237562 163200 237618 164400 6 la_oenb[70]
port 420 nsew signal tristate
rlabel metal2 s 240874 163200 240930 164400 6 la_oenb[71]
port 421 nsew signal tristate
rlabel metal2 s 244278 163200 244334 164400 6 la_oenb[72]
port 422 nsew signal tristate
rlabel metal2 s 247682 163200 247738 164400 6 la_oenb[73]
port 423 nsew signal tristate
rlabel metal2 s 250994 163200 251050 164400 6 la_oenb[74]
port 424 nsew signal tristate
rlabel metal2 s 254398 163200 254454 164400 6 la_oenb[75]
port 425 nsew signal tristate
rlabel metal2 s 257710 163200 257766 164400 6 la_oenb[76]
port 426 nsew signal tristate
rlabel metal2 s 261114 163200 261170 164400 6 la_oenb[77]
port 427 nsew signal tristate
rlabel metal2 s 264426 163200 264482 164400 6 la_oenb[78]
port 428 nsew signal tristate
rlabel metal2 s 267830 163200 267886 164400 6 la_oenb[79]
port 429 nsew signal tristate
rlabel metal2 s 25594 163200 25650 164400 6 la_oenb[7]
port 430 nsew signal tristate
rlabel metal2 s 271234 163200 271290 164400 6 la_oenb[80]
port 431 nsew signal tristate
rlabel metal2 s 274546 163200 274602 164400 6 la_oenb[81]
port 432 nsew signal tristate
rlabel metal2 s 277950 163200 278006 164400 6 la_oenb[82]
port 433 nsew signal tristate
rlabel metal2 s 281262 163200 281318 164400 6 la_oenb[83]
port 434 nsew signal tristate
rlabel metal2 s 284666 163200 284722 164400 6 la_oenb[84]
port 435 nsew signal tristate
rlabel metal2 s 287978 163200 288034 164400 6 la_oenb[85]
port 436 nsew signal tristate
rlabel metal2 s 291382 163200 291438 164400 6 la_oenb[86]
port 437 nsew signal tristate
rlabel metal2 s 294786 163200 294842 164400 6 la_oenb[87]
port 438 nsew signal tristate
rlabel metal2 s 298098 163200 298154 164400 6 la_oenb[88]
port 439 nsew signal tristate
rlabel metal2 s 301502 163200 301558 164400 6 la_oenb[89]
port 440 nsew signal tristate
rlabel metal2 s 28906 163200 28962 164400 6 la_oenb[8]
port 441 nsew signal tristate
rlabel metal2 s 304814 163200 304870 164400 6 la_oenb[90]
port 442 nsew signal tristate
rlabel metal2 s 308218 163200 308274 164400 6 la_oenb[91]
port 443 nsew signal tristate
rlabel metal2 s 311530 163200 311586 164400 6 la_oenb[92]
port 444 nsew signal tristate
rlabel metal2 s 314934 163200 314990 164400 6 la_oenb[93]
port 445 nsew signal tristate
rlabel metal2 s 318338 163200 318394 164400 6 la_oenb[94]
port 446 nsew signal tristate
rlabel metal2 s 321650 163200 321706 164400 6 la_oenb[95]
port 447 nsew signal tristate
rlabel metal2 s 325054 163200 325110 164400 6 la_oenb[96]
port 448 nsew signal tristate
rlabel metal2 s 328366 163200 328422 164400 6 la_oenb[97]
port 449 nsew signal tristate
rlabel metal2 s 331770 163200 331826 164400 6 la_oenb[98]
port 450 nsew signal tristate
rlabel metal2 s 335082 163200 335138 164400 6 la_oenb[99]
port 451 nsew signal tristate
rlabel metal2 s 32310 163200 32366 164400 6 la_oenb[9]
port 452 nsew signal tristate
rlabel metal2 s 2870 163200 2926 164400 6 la_output[0]
port 453 nsew signal tristate
rlabel metal2 s 339314 163200 339370 164400 6 la_output[100]
port 454 nsew signal tristate
rlabel metal2 s 342718 163200 342774 164400 6 la_output[101]
port 455 nsew signal tristate
rlabel metal2 s 346030 163200 346086 164400 6 la_output[102]
port 456 nsew signal tristate
rlabel metal2 s 349434 163200 349490 164400 6 la_output[103]
port 457 nsew signal tristate
rlabel metal2 s 352746 163200 352802 164400 6 la_output[104]
port 458 nsew signal tristate
rlabel metal2 s 356150 163200 356206 164400 6 la_output[105]
port 459 nsew signal tristate
rlabel metal2 s 359554 163200 359610 164400 6 la_output[106]
port 460 nsew signal tristate
rlabel metal2 s 362866 163200 362922 164400 6 la_output[107]
port 461 nsew signal tristate
rlabel metal2 s 366270 163200 366326 164400 6 la_output[108]
port 462 nsew signal tristate
rlabel metal2 s 369582 163200 369638 164400 6 la_output[109]
port 463 nsew signal tristate
rlabel metal2 s 36542 163200 36598 164400 6 la_output[10]
port 464 nsew signal tristate
rlabel metal2 s 372986 163200 373042 164400 6 la_output[110]
port 465 nsew signal tristate
rlabel metal2 s 376298 163200 376354 164400 6 la_output[111]
port 466 nsew signal tristate
rlabel metal2 s 379702 163200 379758 164400 6 la_output[112]
port 467 nsew signal tristate
rlabel metal2 s 383106 163200 383162 164400 6 la_output[113]
port 468 nsew signal tristate
rlabel metal2 s 386418 163200 386474 164400 6 la_output[114]
port 469 nsew signal tristate
rlabel metal2 s 389822 163200 389878 164400 6 la_output[115]
port 470 nsew signal tristate
rlabel metal2 s 393134 163200 393190 164400 6 la_output[116]
port 471 nsew signal tristate
rlabel metal2 s 396538 163200 396594 164400 6 la_output[117]
port 472 nsew signal tristate
rlabel metal2 s 399850 163200 399906 164400 6 la_output[118]
port 473 nsew signal tristate
rlabel metal2 s 403254 163200 403310 164400 6 la_output[119]
port 474 nsew signal tristate
rlabel metal2 s 39854 163200 39910 164400 6 la_output[11]
port 475 nsew signal tristate
rlabel metal2 s 406658 163200 406714 164400 6 la_output[120]
port 476 nsew signal tristate
rlabel metal2 s 409970 163200 410026 164400 6 la_output[121]
port 477 nsew signal tristate
rlabel metal2 s 413374 163200 413430 164400 6 la_output[122]
port 478 nsew signal tristate
rlabel metal2 s 416686 163200 416742 164400 6 la_output[123]
port 479 nsew signal tristate
rlabel metal2 s 420090 163200 420146 164400 6 la_output[124]
port 480 nsew signal tristate
rlabel metal2 s 423402 163200 423458 164400 6 la_output[125]
port 481 nsew signal tristate
rlabel metal2 s 426806 163200 426862 164400 6 la_output[126]
port 482 nsew signal tristate
rlabel metal2 s 430210 163200 430266 164400 6 la_output[127]
port 483 nsew signal tristate
rlabel metal2 s 43258 163200 43314 164400 6 la_output[12]
port 484 nsew signal tristate
rlabel metal2 s 46570 163200 46626 164400 6 la_output[13]
port 485 nsew signal tristate
rlabel metal2 s 49974 163200 50030 164400 6 la_output[14]
port 486 nsew signal tristate
rlabel metal2 s 53378 163200 53434 164400 6 la_output[15]
port 487 nsew signal tristate
rlabel metal2 s 56690 163200 56746 164400 6 la_output[16]
port 488 nsew signal tristate
rlabel metal2 s 60094 163200 60150 164400 6 la_output[17]
port 489 nsew signal tristate
rlabel metal2 s 63406 163200 63462 164400 6 la_output[18]
port 490 nsew signal tristate
rlabel metal2 s 66810 163200 66866 164400 6 la_output[19]
port 491 nsew signal tristate
rlabel metal2 s 6274 163200 6330 164400 6 la_output[1]
port 492 nsew signal tristate
rlabel metal2 s 70122 163200 70178 164400 6 la_output[20]
port 493 nsew signal tristate
rlabel metal2 s 73526 163200 73582 164400 6 la_output[21]
port 494 nsew signal tristate
rlabel metal2 s 76930 163200 76986 164400 6 la_output[22]
port 495 nsew signal tristate
rlabel metal2 s 80242 163200 80298 164400 6 la_output[23]
port 496 nsew signal tristate
rlabel metal2 s 83646 163200 83702 164400 6 la_output[24]
port 497 nsew signal tristate
rlabel metal2 s 86958 163200 87014 164400 6 la_output[25]
port 498 nsew signal tristate
rlabel metal2 s 90362 163200 90418 164400 6 la_output[26]
port 499 nsew signal tristate
rlabel metal2 s 93674 163200 93730 164400 6 la_output[27]
port 500 nsew signal tristate
rlabel metal2 s 97078 163200 97134 164400 6 la_output[28]
port 501 nsew signal tristate
rlabel metal2 s 100482 163200 100538 164400 6 la_output[29]
port 502 nsew signal tristate
rlabel metal2 s 9586 163200 9642 164400 6 la_output[2]
port 503 nsew signal tristate
rlabel metal2 s 103794 163200 103850 164400 6 la_output[30]
port 504 nsew signal tristate
rlabel metal2 s 107198 163200 107254 164400 6 la_output[31]
port 505 nsew signal tristate
rlabel metal2 s 110510 163200 110566 164400 6 la_output[32]
port 506 nsew signal tristate
rlabel metal2 s 113914 163200 113970 164400 6 la_output[33]
port 507 nsew signal tristate
rlabel metal2 s 117226 163200 117282 164400 6 la_output[34]
port 508 nsew signal tristate
rlabel metal2 s 120630 163200 120686 164400 6 la_output[35]
port 509 nsew signal tristate
rlabel metal2 s 124034 163200 124090 164400 6 la_output[36]
port 510 nsew signal tristate
rlabel metal2 s 127346 163200 127402 164400 6 la_output[37]
port 511 nsew signal tristate
rlabel metal2 s 130750 163200 130806 164400 6 la_output[38]
port 512 nsew signal tristate
rlabel metal2 s 134062 163200 134118 164400 6 la_output[39]
port 513 nsew signal tristate
rlabel metal2 s 12990 163200 13046 164400 6 la_output[3]
port 514 nsew signal tristate
rlabel metal2 s 137466 163200 137522 164400 6 la_output[40]
port 515 nsew signal tristate
rlabel metal2 s 140778 163200 140834 164400 6 la_output[41]
port 516 nsew signal tristate
rlabel metal2 s 144182 163200 144238 164400 6 la_output[42]
port 517 nsew signal tristate
rlabel metal2 s 147586 163200 147642 164400 6 la_output[43]
port 518 nsew signal tristate
rlabel metal2 s 150898 163200 150954 164400 6 la_output[44]
port 519 nsew signal tristate
rlabel metal2 s 154302 163200 154358 164400 6 la_output[45]
port 520 nsew signal tristate
rlabel metal2 s 157614 163200 157670 164400 6 la_output[46]
port 521 nsew signal tristate
rlabel metal2 s 161018 163200 161074 164400 6 la_output[47]
port 522 nsew signal tristate
rlabel metal2 s 164330 163200 164386 164400 6 la_output[48]
port 523 nsew signal tristate
rlabel metal2 s 167734 163200 167790 164400 6 la_output[49]
port 524 nsew signal tristate
rlabel metal2 s 16302 163200 16358 164400 6 la_output[4]
port 525 nsew signal tristate
rlabel metal2 s 171138 163200 171194 164400 6 la_output[50]
port 526 nsew signal tristate
rlabel metal2 s 174450 163200 174506 164400 6 la_output[51]
port 527 nsew signal tristate
rlabel metal2 s 177854 163200 177910 164400 6 la_output[52]
port 528 nsew signal tristate
rlabel metal2 s 181166 163200 181222 164400 6 la_output[53]
port 529 nsew signal tristate
rlabel metal2 s 184570 163200 184626 164400 6 la_output[54]
port 530 nsew signal tristate
rlabel metal2 s 187882 163200 187938 164400 6 la_output[55]
port 531 nsew signal tristate
rlabel metal2 s 191286 163200 191342 164400 6 la_output[56]
port 532 nsew signal tristate
rlabel metal2 s 194690 163200 194746 164400 6 la_output[57]
port 533 nsew signal tristate
rlabel metal2 s 198002 163200 198058 164400 6 la_output[58]
port 534 nsew signal tristate
rlabel metal2 s 201406 163200 201462 164400 6 la_output[59]
port 535 nsew signal tristate
rlabel metal2 s 19706 163200 19762 164400 6 la_output[5]
port 536 nsew signal tristate
rlabel metal2 s 204718 163200 204774 164400 6 la_output[60]
port 537 nsew signal tristate
rlabel metal2 s 208122 163200 208178 164400 6 la_output[61]
port 538 nsew signal tristate
rlabel metal2 s 211434 163200 211490 164400 6 la_output[62]
port 539 nsew signal tristate
rlabel metal2 s 214838 163200 214894 164400 6 la_output[63]
port 540 nsew signal tristate
rlabel metal2 s 218242 163200 218298 164400 6 la_output[64]
port 541 nsew signal tristate
rlabel metal2 s 221554 163200 221610 164400 6 la_output[65]
port 542 nsew signal tristate
rlabel metal2 s 224958 163200 225014 164400 6 la_output[66]
port 543 nsew signal tristate
rlabel metal2 s 228270 163200 228326 164400 6 la_output[67]
port 544 nsew signal tristate
rlabel metal2 s 231674 163200 231730 164400 6 la_output[68]
port 545 nsew signal tristate
rlabel metal2 s 234986 163200 235042 164400 6 la_output[69]
port 546 nsew signal tristate
rlabel metal2 s 23018 163200 23074 164400 6 la_output[6]
port 547 nsew signal tristate
rlabel metal2 s 238390 163200 238446 164400 6 la_output[70]
port 548 nsew signal tristate
rlabel metal2 s 241794 163200 241850 164400 6 la_output[71]
port 549 nsew signal tristate
rlabel metal2 s 245106 163200 245162 164400 6 la_output[72]
port 550 nsew signal tristate
rlabel metal2 s 248510 163200 248566 164400 6 la_output[73]
port 551 nsew signal tristate
rlabel metal2 s 251822 163200 251878 164400 6 la_output[74]
port 552 nsew signal tristate
rlabel metal2 s 255226 163200 255282 164400 6 la_output[75]
port 553 nsew signal tristate
rlabel metal2 s 258538 163200 258594 164400 6 la_output[76]
port 554 nsew signal tristate
rlabel metal2 s 261942 163200 261998 164400 6 la_output[77]
port 555 nsew signal tristate
rlabel metal2 s 265346 163200 265402 164400 6 la_output[78]
port 556 nsew signal tristate
rlabel metal2 s 268658 163200 268714 164400 6 la_output[79]
port 557 nsew signal tristate
rlabel metal2 s 26422 163200 26478 164400 6 la_output[7]
port 558 nsew signal tristate
rlabel metal2 s 272062 163200 272118 164400 6 la_output[80]
port 559 nsew signal tristate
rlabel metal2 s 275374 163200 275430 164400 6 la_output[81]
port 560 nsew signal tristate
rlabel metal2 s 278778 163200 278834 164400 6 la_output[82]
port 561 nsew signal tristate
rlabel metal2 s 282090 163200 282146 164400 6 la_output[83]
port 562 nsew signal tristate
rlabel metal2 s 285494 163200 285550 164400 6 la_output[84]
port 563 nsew signal tristate
rlabel metal2 s 288898 163200 288954 164400 6 la_output[85]
port 564 nsew signal tristate
rlabel metal2 s 292210 163200 292266 164400 6 la_output[86]
port 565 nsew signal tristate
rlabel metal2 s 295614 163200 295670 164400 6 la_output[87]
port 566 nsew signal tristate
rlabel metal2 s 298926 163200 298982 164400 6 la_output[88]
port 567 nsew signal tristate
rlabel metal2 s 302330 163200 302386 164400 6 la_output[89]
port 568 nsew signal tristate
rlabel metal2 s 29826 163200 29882 164400 6 la_output[8]
port 569 nsew signal tristate
rlabel metal2 s 305642 163200 305698 164400 6 la_output[90]
port 570 nsew signal tristate
rlabel metal2 s 309046 163200 309102 164400 6 la_output[91]
port 571 nsew signal tristate
rlabel metal2 s 312450 163200 312506 164400 6 la_output[92]
port 572 nsew signal tristate
rlabel metal2 s 315762 163200 315818 164400 6 la_output[93]
port 573 nsew signal tristate
rlabel metal2 s 319166 163200 319222 164400 6 la_output[94]
port 574 nsew signal tristate
rlabel metal2 s 322478 163200 322534 164400 6 la_output[95]
port 575 nsew signal tristate
rlabel metal2 s 325882 163200 325938 164400 6 la_output[96]
port 576 nsew signal tristate
rlabel metal2 s 329194 163200 329250 164400 6 la_output[97]
port 577 nsew signal tristate
rlabel metal2 s 332598 163200 332654 164400 6 la_output[98]
port 578 nsew signal tristate
rlabel metal2 s 336002 163200 336058 164400 6 la_output[99]
port 579 nsew signal tristate
rlabel metal2 s 33138 163200 33194 164400 6 la_output[9]
port 580 nsew signal tristate
rlabel metal2 s 431038 163200 431094 164400 6 mprj_ack_i
port 581 nsew signal input
rlabel metal2 s 435178 163200 435234 164400 6 mprj_adr_o[0]
port 582 nsew signal tristate
rlabel metal2 s 463790 163200 463846 164400 6 mprj_adr_o[10]
port 583 nsew signal tristate
rlabel metal2 s 466366 163200 466422 164400 6 mprj_adr_o[11]
port 584 nsew signal tristate
rlabel metal2 s 468850 163200 468906 164400 6 mprj_adr_o[12]
port 585 nsew signal tristate
rlabel metal2 s 471426 163200 471482 164400 6 mprj_adr_o[13]
port 586 nsew signal tristate
rlabel metal2 s 473910 163200 473966 164400 6 mprj_adr_o[14]
port 587 nsew signal tristate
rlabel metal2 s 476394 163200 476450 164400 6 mprj_adr_o[15]
port 588 nsew signal tristate
rlabel metal2 s 478970 163200 479026 164400 6 mprj_adr_o[16]
port 589 nsew signal tristate
rlabel metal2 s 481454 163200 481510 164400 6 mprj_adr_o[17]
port 590 nsew signal tristate
rlabel metal2 s 484030 163200 484086 164400 6 mprj_adr_o[18]
port 591 nsew signal tristate
rlabel metal2 s 486514 163200 486570 164400 6 mprj_adr_o[19]
port 592 nsew signal tristate
rlabel metal2 s 438582 163200 438638 164400 6 mprj_adr_o[1]
port 593 nsew signal tristate
rlabel metal2 s 489090 163200 489146 164400 6 mprj_adr_o[20]
port 594 nsew signal tristate
rlabel metal2 s 491574 163200 491630 164400 6 mprj_adr_o[21]
port 595 nsew signal tristate
rlabel metal2 s 494058 163200 494114 164400 6 mprj_adr_o[22]
port 596 nsew signal tristate
rlabel metal2 s 496634 163200 496690 164400 6 mprj_adr_o[23]
port 597 nsew signal tristate
rlabel metal2 s 499118 163200 499174 164400 6 mprj_adr_o[24]
port 598 nsew signal tristate
rlabel metal2 s 501694 163200 501750 164400 6 mprj_adr_o[25]
port 599 nsew signal tristate
rlabel metal2 s 504178 163200 504234 164400 6 mprj_adr_o[26]
port 600 nsew signal tristate
rlabel metal2 s 506754 163200 506810 164400 6 mprj_adr_o[27]
port 601 nsew signal tristate
rlabel metal2 s 509238 163200 509294 164400 6 mprj_adr_o[28]
port 602 nsew signal tristate
rlabel metal2 s 511722 163200 511778 164400 6 mprj_adr_o[29]
port 603 nsew signal tristate
rlabel metal2 s 441986 163200 442042 164400 6 mprj_adr_o[2]
port 604 nsew signal tristate
rlabel metal2 s 514298 163200 514354 164400 6 mprj_adr_o[30]
port 605 nsew signal tristate
rlabel metal2 s 516782 163200 516838 164400 6 mprj_adr_o[31]
port 606 nsew signal tristate
rlabel metal2 s 445298 163200 445354 164400 6 mprj_adr_o[3]
port 607 nsew signal tristate
rlabel metal2 s 448702 163200 448758 164400 6 mprj_adr_o[4]
port 608 nsew signal tristate
rlabel metal2 s 451186 163200 451242 164400 6 mprj_adr_o[5]
port 609 nsew signal tristate
rlabel metal2 s 453762 163200 453818 164400 6 mprj_adr_o[6]
port 610 nsew signal tristate
rlabel metal2 s 456246 163200 456302 164400 6 mprj_adr_o[7]
port 611 nsew signal tristate
rlabel metal2 s 458730 163200 458786 164400 6 mprj_adr_o[8]
port 612 nsew signal tristate
rlabel metal2 s 461306 163200 461362 164400 6 mprj_adr_o[9]
port 613 nsew signal tristate
rlabel metal2 s 431866 163200 431922 164400 6 mprj_cyc_o
port 614 nsew signal tristate
rlabel metal2 s 436098 163200 436154 164400 6 mprj_dat_i[0]
port 615 nsew signal input
rlabel metal2 s 464618 163200 464674 164400 6 mprj_dat_i[10]
port 616 nsew signal input
rlabel metal2 s 467194 163200 467250 164400 6 mprj_dat_i[11]
port 617 nsew signal input
rlabel metal2 s 469678 163200 469734 164400 6 mprj_dat_i[12]
port 618 nsew signal input
rlabel metal2 s 472254 163200 472310 164400 6 mprj_dat_i[13]
port 619 nsew signal input
rlabel metal2 s 474738 163200 474794 164400 6 mprj_dat_i[14]
port 620 nsew signal input
rlabel metal2 s 477314 163200 477370 164400 6 mprj_dat_i[15]
port 621 nsew signal input
rlabel metal2 s 479798 163200 479854 164400 6 mprj_dat_i[16]
port 622 nsew signal input
rlabel metal2 s 482282 163200 482338 164400 6 mprj_dat_i[17]
port 623 nsew signal input
rlabel metal2 s 484858 163200 484914 164400 6 mprj_dat_i[18]
port 624 nsew signal input
rlabel metal2 s 487342 163200 487398 164400 6 mprj_dat_i[19]
port 625 nsew signal input
rlabel metal2 s 439410 163200 439466 164400 6 mprj_dat_i[1]
port 626 nsew signal input
rlabel metal2 s 489918 163200 489974 164400 6 mprj_dat_i[20]
port 627 nsew signal input
rlabel metal2 s 492402 163200 492458 164400 6 mprj_dat_i[21]
port 628 nsew signal input
rlabel metal2 s 494978 163200 495034 164400 6 mprj_dat_i[22]
port 629 nsew signal input
rlabel metal2 s 497462 163200 497518 164400 6 mprj_dat_i[23]
port 630 nsew signal input
rlabel metal2 s 499946 163200 500002 164400 6 mprj_dat_i[24]
port 631 nsew signal input
rlabel metal2 s 502522 163200 502578 164400 6 mprj_dat_i[25]
port 632 nsew signal input
rlabel metal2 s 505006 163200 505062 164400 6 mprj_dat_i[26]
port 633 nsew signal input
rlabel metal2 s 507582 163200 507638 164400 6 mprj_dat_i[27]
port 634 nsew signal input
rlabel metal2 s 510066 163200 510122 164400 6 mprj_dat_i[28]
port 635 nsew signal input
rlabel metal2 s 512642 163200 512698 164400 6 mprj_dat_i[29]
port 636 nsew signal input
rlabel metal2 s 442814 163200 442870 164400 6 mprj_dat_i[2]
port 637 nsew signal input
rlabel metal2 s 515126 163200 515182 164400 6 mprj_dat_i[30]
port 638 nsew signal input
rlabel metal2 s 517610 163200 517666 164400 6 mprj_dat_i[31]
port 639 nsew signal input
rlabel metal2 s 446126 163200 446182 164400 6 mprj_dat_i[3]
port 640 nsew signal input
rlabel metal2 s 449530 163200 449586 164400 6 mprj_dat_i[4]
port 641 nsew signal input
rlabel metal2 s 452014 163200 452070 164400 6 mprj_dat_i[5]
port 642 nsew signal input
rlabel metal2 s 454590 163200 454646 164400 6 mprj_dat_i[6]
port 643 nsew signal input
rlabel metal2 s 457074 163200 457130 164400 6 mprj_dat_i[7]
port 644 nsew signal input
rlabel metal2 s 459650 163200 459706 164400 6 mprj_dat_i[8]
port 645 nsew signal input
rlabel metal2 s 462134 163200 462190 164400 6 mprj_dat_i[9]
port 646 nsew signal input
rlabel metal2 s 436926 163200 436982 164400 6 mprj_dat_o[0]
port 647 nsew signal tristate
rlabel metal2 s 465538 163200 465594 164400 6 mprj_dat_o[10]
port 648 nsew signal tristate
rlabel metal2 s 468022 163200 468078 164400 6 mprj_dat_o[11]
port 649 nsew signal tristate
rlabel metal2 s 470506 163200 470562 164400 6 mprj_dat_o[12]
port 650 nsew signal tristate
rlabel metal2 s 473082 163200 473138 164400 6 mprj_dat_o[13]
port 651 nsew signal tristate
rlabel metal2 s 475566 163200 475622 164400 6 mprj_dat_o[14]
port 652 nsew signal tristate
rlabel metal2 s 478142 163200 478198 164400 6 mprj_dat_o[15]
port 653 nsew signal tristate
rlabel metal2 s 480626 163200 480682 164400 6 mprj_dat_o[16]
port 654 nsew signal tristate
rlabel metal2 s 483202 163200 483258 164400 6 mprj_dat_o[17]
port 655 nsew signal tristate
rlabel metal2 s 485686 163200 485742 164400 6 mprj_dat_o[18]
port 656 nsew signal tristate
rlabel metal2 s 488170 163200 488226 164400 6 mprj_dat_o[19]
port 657 nsew signal tristate
rlabel metal2 s 440238 163200 440294 164400 6 mprj_dat_o[1]
port 658 nsew signal tristate
rlabel metal2 s 490746 163200 490802 164400 6 mprj_dat_o[20]
port 659 nsew signal tristate
rlabel metal2 s 493230 163200 493286 164400 6 mprj_dat_o[21]
port 660 nsew signal tristate
rlabel metal2 s 495806 163200 495862 164400 6 mprj_dat_o[22]
port 661 nsew signal tristate
rlabel metal2 s 498290 163200 498346 164400 6 mprj_dat_o[23]
port 662 nsew signal tristate
rlabel metal2 s 500866 163200 500922 164400 6 mprj_dat_o[24]
port 663 nsew signal tristate
rlabel metal2 s 503350 163200 503406 164400 6 mprj_dat_o[25]
port 664 nsew signal tristate
rlabel metal2 s 505834 163200 505890 164400 6 mprj_dat_o[26]
port 665 nsew signal tristate
rlabel metal2 s 508410 163200 508466 164400 6 mprj_dat_o[27]
port 666 nsew signal tristate
rlabel metal2 s 510894 163200 510950 164400 6 mprj_dat_o[28]
port 667 nsew signal tristate
rlabel metal2 s 513470 163200 513526 164400 6 mprj_dat_o[29]
port 668 nsew signal tristate
rlabel metal2 s 443642 163200 443698 164400 6 mprj_dat_o[2]
port 669 nsew signal tristate
rlabel metal2 s 515954 163200 516010 164400 6 mprj_dat_o[30]
port 670 nsew signal tristate
rlabel metal2 s 518530 163200 518586 164400 6 mprj_dat_o[31]
port 671 nsew signal tristate
rlabel metal2 s 446954 163200 447010 164400 6 mprj_dat_o[3]
port 672 nsew signal tristate
rlabel metal2 s 450358 163200 450414 164400 6 mprj_dat_o[4]
port 673 nsew signal tristate
rlabel metal2 s 452842 163200 452898 164400 6 mprj_dat_o[5]
port 674 nsew signal tristate
rlabel metal2 s 455418 163200 455474 164400 6 mprj_dat_o[6]
port 675 nsew signal tristate
rlabel metal2 s 457902 163200 457958 164400 6 mprj_dat_o[7]
port 676 nsew signal tristate
rlabel metal2 s 460478 163200 460534 164400 6 mprj_dat_o[8]
port 677 nsew signal tristate
rlabel metal2 s 462962 163200 463018 164400 6 mprj_dat_o[9]
port 678 nsew signal tristate
rlabel metal2 s 437754 163200 437810 164400 6 mprj_sel_o[0]
port 679 nsew signal tristate
rlabel metal2 s 441066 163200 441122 164400 6 mprj_sel_o[1]
port 680 nsew signal tristate
rlabel metal2 s 444470 163200 444526 164400 6 mprj_sel_o[2]
port 681 nsew signal tristate
rlabel metal2 s 447874 163200 447930 164400 6 mprj_sel_o[3]
port 682 nsew signal tristate
rlabel metal2 s 432694 163200 432750 164400 6 mprj_stb_o
port 683 nsew signal tristate
rlabel metal2 s 433522 163200 433578 164400 6 mprj_wb_iena
port 684 nsew signal tristate
rlabel metal2 s 434350 163200 434406 164400 6 mprj_we_o
port 685 nsew signal tristate
rlabel metal3 s 523200 89360 524400 89480 6 qspi_enabled
port 686 nsew signal tristate
rlabel metal3 s 523200 83376 524400 83496 6 ser_rx
port 687 nsew signal input
rlabel metal3 s 523200 84872 524400 84992 6 ser_tx
port 688 nsew signal tristate
rlabel metal3 s 523200 80384 524400 80504 6 spi_csb
port 689 nsew signal tristate
rlabel metal3 s 523200 86368 524400 86488 6 spi_enabled
port 690 nsew signal tristate
rlabel metal3 s 523200 78888 524400 79008 6 spi_sck
port 691 nsew signal tristate
rlabel metal3 s 523200 81880 524400 82000 6 spi_sdi
port 692 nsew signal input
rlabel metal3 s 523200 77392 524400 77512 6 spi_sdo
port 693 nsew signal tristate
rlabel metal3 s 523200 75896 524400 76016 6 spi_sdoenb
port 694 nsew signal tristate
rlabel metal3 s 523200 2184 524400 2304 6 sram_ro_addr[0]
port 695 nsew signal input
rlabel metal3 s 523200 3680 524400 3800 6 sram_ro_addr[1]
port 696 nsew signal input
rlabel metal3 s 523200 5176 524400 5296 6 sram_ro_addr[2]
port 697 nsew signal input
rlabel metal3 s 523200 6672 524400 6792 6 sram_ro_addr[3]
port 698 nsew signal input
rlabel metal3 s 523200 8168 524400 8288 6 sram_ro_addr[4]
port 699 nsew signal input
rlabel metal3 s 523200 9664 524400 9784 6 sram_ro_addr[5]
port 700 nsew signal input
rlabel metal3 s 523200 11160 524400 11280 6 sram_ro_addr[6]
port 701 nsew signal input
rlabel metal3 s 523200 12656 524400 12776 6 sram_ro_addr[7]
port 702 nsew signal input
rlabel metal3 s 523200 14152 524400 14272 6 sram_ro_clk
port 703 nsew signal input
rlabel metal3 s 523200 688 524400 808 6 sram_ro_csb
port 704 nsew signal input
rlabel metal3 s 523200 15648 524400 15768 6 sram_ro_data[0]
port 705 nsew signal tristate
rlabel metal3 s 523200 30744 524400 30864 6 sram_ro_data[10]
port 706 nsew signal tristate
rlabel metal3 s 523200 32240 524400 32360 6 sram_ro_data[11]
port 707 nsew signal tristate
rlabel metal3 s 523200 33736 524400 33856 6 sram_ro_data[12]
port 708 nsew signal tristate
rlabel metal3 s 523200 35232 524400 35352 6 sram_ro_data[13]
port 709 nsew signal tristate
rlabel metal3 s 523200 36728 524400 36848 6 sram_ro_data[14]
port 710 nsew signal tristate
rlabel metal3 s 523200 38224 524400 38344 6 sram_ro_data[15]
port 711 nsew signal tristate
rlabel metal3 s 523200 39720 524400 39840 6 sram_ro_data[16]
port 712 nsew signal tristate
rlabel metal3 s 523200 41216 524400 41336 6 sram_ro_data[17]
port 713 nsew signal tristate
rlabel metal3 s 523200 42712 524400 42832 6 sram_ro_data[18]
port 714 nsew signal tristate
rlabel metal3 s 523200 44208 524400 44328 6 sram_ro_data[19]
port 715 nsew signal tristate
rlabel metal3 s 523200 17144 524400 17264 6 sram_ro_data[1]
port 716 nsew signal tristate
rlabel metal3 s 523200 45704 524400 45824 6 sram_ro_data[20]
port 717 nsew signal tristate
rlabel metal3 s 523200 47200 524400 47320 6 sram_ro_data[21]
port 718 nsew signal tristate
rlabel metal3 s 523200 48832 524400 48952 6 sram_ro_data[22]
port 719 nsew signal tristate
rlabel metal3 s 523200 50328 524400 50448 6 sram_ro_data[23]
port 720 nsew signal tristate
rlabel metal3 s 523200 51824 524400 51944 6 sram_ro_data[24]
port 721 nsew signal tristate
rlabel metal3 s 523200 53320 524400 53440 6 sram_ro_data[25]
port 722 nsew signal tristate
rlabel metal3 s 523200 54816 524400 54936 6 sram_ro_data[26]
port 723 nsew signal tristate
rlabel metal3 s 523200 56312 524400 56432 6 sram_ro_data[27]
port 724 nsew signal tristate
rlabel metal3 s 523200 57808 524400 57928 6 sram_ro_data[28]
port 725 nsew signal tristate
rlabel metal3 s 523200 59304 524400 59424 6 sram_ro_data[29]
port 726 nsew signal tristate
rlabel metal3 s 523200 18640 524400 18760 6 sram_ro_data[2]
port 727 nsew signal tristate
rlabel metal3 s 523200 60800 524400 60920 6 sram_ro_data[30]
port 728 nsew signal tristate
rlabel metal3 s 523200 62296 524400 62416 6 sram_ro_data[31]
port 729 nsew signal tristate
rlabel metal3 s 523200 20136 524400 20256 6 sram_ro_data[3]
port 730 nsew signal tristate
rlabel metal3 s 523200 21632 524400 21752 6 sram_ro_data[4]
port 731 nsew signal tristate
rlabel metal3 s 523200 23128 524400 23248 6 sram_ro_data[5]
port 732 nsew signal tristate
rlabel metal3 s 523200 24760 524400 24880 6 sram_ro_data[6]
port 733 nsew signal tristate
rlabel metal3 s 523200 26256 524400 26376 6 sram_ro_data[7]
port 734 nsew signal tristate
rlabel metal3 s 523200 27752 524400 27872 6 sram_ro_data[8]
port 735 nsew signal tristate
rlabel metal3 s 523200 29248 524400 29368 6 sram_ro_data[9]
port 736 nsew signal tristate
rlabel metal3 s 523200 69776 524400 69896 6 trap
port 737 nsew signal tristate
rlabel metal3 s 523200 87864 524400 87984 6 uart_enabled
port 738 nsew signal tristate
rlabel metal2 s 519358 163200 519414 164400 6 user_irq_ena[0]
port 739 nsew signal tristate
rlabel metal2 s 520186 163200 520242 164400 6 user_irq_ena[1]
port 740 nsew signal tristate
rlabel metal2 s 521014 163200 521070 164400 6 user_irq_ena[2]
port 741 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 524000 164000
<< end >>
