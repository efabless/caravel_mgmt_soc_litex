magic
tech sky130A
magscale 1 2
timestamp 1638213420
<< metal1 >>
rect 338408 160092 339816 160120
rect 63402 160012 63408 160064
rect 63460 160052 63466 160064
rect 146478 160052 146484 160064
rect 63460 160024 146484 160052
rect 63460 160012 63466 160024
rect 146478 160012 146484 160024
rect 146536 160012 146542 160064
rect 146754 160012 146760 160064
rect 146812 160052 146818 160064
rect 154482 160052 154488 160064
rect 146812 160024 154488 160052
rect 146812 160012 146818 160024
rect 154482 160012 154488 160024
rect 154540 160012 154546 160064
rect 156782 160012 156788 160064
rect 156840 160052 156846 160064
rect 191742 160052 191748 160064
rect 156840 160024 191748 160052
rect 156840 160012 156846 160024
rect 191742 160012 191748 160024
rect 191800 160012 191806 160064
rect 197170 160012 197176 160064
rect 197228 160052 197234 160064
rect 207106 160052 207112 160064
rect 197228 160024 207112 160052
rect 197228 160012 197234 160024
rect 207106 160012 207112 160024
rect 207164 160012 207170 160064
rect 211430 160012 211436 160064
rect 211488 160052 211494 160064
rect 280154 160052 280160 160064
rect 211488 160024 280160 160052
rect 211488 160012 211494 160024
rect 280154 160012 280160 160024
rect 280212 160012 280218 160064
rect 281258 160012 281264 160064
rect 281316 160052 281322 160064
rect 332686 160052 332692 160064
rect 281316 160024 332692 160052
rect 281316 160012 281322 160024
rect 332686 160012 332692 160024
rect 332744 160012 332750 160064
rect 335078 160012 335084 160064
rect 335136 160052 335142 160064
rect 338408 160052 338436 160092
rect 335136 160024 338436 160052
rect 335136 160012 335142 160024
rect 338482 160012 338488 160064
rect 338540 160052 338546 160064
rect 339678 160052 339684 160064
rect 338540 160024 339684 160052
rect 338540 160012 338546 160024
rect 339678 160012 339684 160024
rect 339736 160012 339742 160064
rect 339788 160052 339816 160092
rect 374362 160052 374368 160064
rect 339788 160024 374368 160052
rect 374362 160012 374368 160024
rect 374420 160012 374426 160064
rect 378870 160012 378876 160064
rect 378928 160052 378934 160064
rect 398098 160052 398104 160064
rect 378928 160024 398104 160052
rect 378928 160012 378934 160024
rect 398098 160012 398104 160024
rect 398156 160012 398162 160064
rect 409966 160012 409972 160064
rect 410024 160052 410030 160064
rect 417602 160052 417608 160064
rect 410024 160024 417608 160052
rect 410024 160012 410030 160024
rect 417602 160012 417608 160024
rect 417660 160012 417666 160064
rect 454586 160012 454592 160064
rect 454644 160052 454650 160064
rect 465442 160052 465448 160064
rect 454644 160024 465448 160052
rect 454644 160012 454650 160024
rect 465442 160012 465448 160024
rect 465500 160012 465506 160064
rect 25590 159944 25596 159996
rect 25648 159984 25654 159996
rect 109770 159984 109776 159996
rect 25648 159956 109776 159984
rect 25648 159944 25654 159956
rect 109770 159944 109776 159956
rect 109828 159944 109834 159996
rect 117222 159944 117228 159996
rect 117280 159984 117286 159996
rect 191650 159984 191656 159996
rect 117280 159956 191656 159984
rect 117280 159944 117286 159956
rect 191650 159944 191656 159956
rect 191708 159944 191714 159996
rect 197998 159944 198004 159996
rect 198056 159984 198062 159996
rect 269850 159984 269856 159996
rect 198056 159956 269856 159984
rect 198056 159944 198062 159956
rect 269850 159944 269856 159956
rect 269908 159944 269914 159996
rect 271230 159944 271236 159996
rect 271288 159984 271294 159996
rect 272518 159984 272524 159996
rect 271288 159956 272524 159984
rect 271288 159944 271294 159956
rect 272518 159944 272524 159956
rect 272576 159944 272582 159996
rect 275370 159944 275376 159996
rect 275428 159984 275434 159996
rect 328454 159984 328460 159996
rect 275428 159956 328460 159984
rect 275428 159944 275434 159956
rect 328454 159944 328460 159956
rect 328512 159944 328518 159996
rect 329190 159944 329196 159996
rect 329248 159984 329254 159996
rect 369854 159984 369860 159996
rect 329248 159956 369860 159984
rect 329248 159944 329254 159956
rect 369854 159944 369860 159956
rect 369912 159944 369918 159996
rect 374638 159944 374644 159996
rect 374696 159984 374702 159996
rect 388346 159984 388352 159996
rect 374696 159956 388352 159984
rect 374696 159944 374702 159956
rect 388346 159944 388352 159956
rect 388404 159944 388410 159996
rect 389818 159944 389824 159996
rect 389876 159984 389882 159996
rect 413922 159984 413928 159996
rect 389876 159956 413928 159984
rect 389876 159944 389882 159956
rect 413922 159944 413928 159956
rect 413980 159944 413986 159996
rect 452838 159944 452844 159996
rect 452896 159984 452902 159996
rect 464246 159984 464252 159996
rect 452896 159956 464252 159984
rect 452896 159944 452902 159956
rect 464246 159944 464252 159956
rect 464304 159944 464310 159996
rect 468018 159944 468024 159996
rect 468076 159984 468082 159996
rect 476022 159984 476028 159996
rect 468076 159956 476028 159984
rect 468076 159944 468082 159956
rect 476022 159944 476028 159956
rect 476080 159944 476086 159996
rect 76926 159876 76932 159928
rect 76984 159916 76990 159928
rect 162578 159916 162584 159928
rect 76984 159888 162584 159916
rect 76984 159876 76990 159888
rect 162578 159876 162584 159888
rect 162636 159876 162642 159928
rect 166902 159876 166908 159928
rect 166960 159916 166966 159928
rect 186406 159916 186412 159928
rect 166960 159888 186412 159916
rect 166960 159876 166966 159888
rect 186406 159876 186412 159888
rect 186464 159876 186470 159928
rect 191282 159876 191288 159928
rect 191340 159916 191346 159928
rect 264882 159916 264888 159928
rect 191340 159888 264888 159916
rect 191340 159876 191346 159888
rect 264882 159876 264888 159888
rect 264940 159876 264946 159928
rect 268654 159876 268660 159928
rect 268712 159916 268718 159928
rect 323670 159916 323676 159928
rect 268712 159888 323676 159916
rect 268712 159876 268718 159888
rect 323670 159876 323676 159888
rect 323728 159876 323734 159928
rect 328362 159876 328368 159928
rect 328420 159916 328426 159928
rect 369210 159916 369216 159928
rect 328420 159888 369216 159916
rect 328420 159876 328426 159888
rect 369210 159876 369216 159888
rect 369268 159876 369274 159928
rect 372154 159876 372160 159928
rect 372212 159916 372218 159928
rect 396258 159916 396264 159928
rect 372212 159888 396264 159916
rect 372212 159876 372218 159888
rect 396258 159876 396264 159888
rect 396316 159876 396322 159928
rect 403250 159876 403256 159928
rect 403308 159916 403314 159928
rect 416590 159916 416596 159928
rect 403308 159888 416596 159916
rect 403308 159876 403314 159888
rect 416590 159876 416596 159888
rect 416648 159876 416654 159928
rect 455414 159876 455420 159928
rect 455472 159916 455478 159928
rect 466638 159916 466644 159928
rect 455472 159888 466644 159916
rect 455472 159876 455478 159888
rect 466638 159876 466644 159888
rect 466696 159876 466702 159928
rect 467190 159876 467196 159928
rect 467248 159916 467254 159928
rect 473354 159916 473360 159928
rect 467248 159888 473360 159916
rect 467248 159876 467254 159888
rect 473354 159876 473360 159888
rect 473412 159876 473418 159928
rect 70118 159808 70124 159860
rect 70176 159848 70182 159860
rect 156414 159848 156420 159860
rect 70176 159820 156420 159848
rect 70176 159808 70182 159820
rect 156414 159808 156420 159820
rect 156472 159808 156478 159860
rect 156598 159808 156604 159860
rect 156656 159848 156662 159860
rect 160094 159848 160100 159860
rect 156656 159820 160100 159848
rect 156656 159808 156662 159820
rect 160094 159808 160100 159820
rect 160152 159808 160158 159860
rect 180702 159848 180708 159860
rect 161446 159820 180708 159848
rect 56686 159740 56692 159792
rect 56744 159780 56750 159792
rect 137278 159780 137284 159792
rect 56744 159752 137284 159780
rect 56744 159740 56750 159752
rect 137278 159740 137284 159752
rect 137336 159740 137342 159792
rect 137370 159740 137376 159792
rect 137428 159780 137434 159792
rect 139670 159780 139676 159792
rect 137428 159752 139676 159780
rect 137428 159740 137434 159752
rect 139670 159740 139676 159752
rect 139728 159740 139734 159792
rect 139946 159740 139952 159792
rect 140004 159780 140010 159792
rect 147030 159780 147036 159792
rect 140004 159752 147036 159780
rect 140004 159740 140010 159752
rect 147030 159740 147036 159752
rect 147088 159740 147094 159792
rect 153470 159740 153476 159792
rect 153528 159780 153534 159792
rect 161446 159780 161474 159820
rect 180702 159808 180708 159820
rect 180760 159808 180766 159860
rect 184566 159808 184572 159860
rect 184624 159848 184630 159860
rect 259546 159848 259552 159860
rect 184624 159820 259552 159848
rect 184624 159808 184630 159820
rect 259546 159808 259552 159820
rect 259604 159808 259610 159860
rect 261938 159808 261944 159860
rect 261996 159848 262002 159860
rect 312354 159848 312360 159860
rect 261996 159820 312360 159848
rect 261996 159808 262002 159820
rect 312354 159808 312360 159820
rect 312412 159808 312418 159860
rect 312446 159808 312452 159860
rect 312504 159848 312510 159860
rect 313366 159848 313372 159860
rect 312504 159820 313372 159848
rect 312504 159808 312510 159820
rect 313366 159808 313372 159820
rect 313424 159808 313430 159860
rect 322474 159808 322480 159860
rect 322532 159848 322538 159860
rect 364794 159848 364800 159860
rect 322532 159820 364800 159848
rect 322532 159808 322538 159820
rect 364794 159808 364800 159820
rect 364852 159808 364858 159860
rect 376294 159808 376300 159860
rect 376352 159848 376358 159860
rect 405826 159848 405832 159860
rect 376352 159820 405832 159848
rect 376352 159808 376358 159820
rect 405826 159808 405832 159820
rect 405884 159808 405890 159860
rect 449526 159808 449532 159860
rect 449584 159848 449590 159860
rect 459554 159848 459560 159860
rect 449584 159820 459560 159848
rect 449584 159808 449590 159820
rect 459554 159808 459560 159820
rect 459612 159808 459618 159860
rect 472250 159808 472256 159860
rect 472308 159848 472314 159860
rect 479058 159848 479064 159860
rect 472308 159820 479064 159848
rect 472308 159808 472314 159820
rect 479058 159808 479064 159820
rect 479116 159808 479122 159860
rect 153528 159752 161474 159780
rect 153528 159740 153534 159752
rect 177850 159740 177856 159792
rect 177908 159780 177914 159792
rect 254302 159780 254308 159792
rect 177908 159752 254308 159780
rect 177908 159740 177914 159752
rect 254302 159740 254308 159752
rect 254360 159740 254366 159792
rect 255222 159740 255228 159792
rect 255280 159780 255286 159792
rect 313458 159780 313464 159792
rect 255280 159752 313464 159780
rect 255280 159740 255286 159752
rect 313458 159740 313464 159752
rect 313516 159740 313522 159792
rect 314102 159740 314108 159792
rect 314160 159780 314166 159792
rect 357986 159780 357992 159792
rect 314160 159752 357992 159780
rect 314160 159740 314166 159752
rect 357986 159740 357992 159752
rect 358044 159740 358050 159792
rect 365438 159740 365444 159792
rect 365496 159780 365502 159792
rect 395430 159780 395436 159792
rect 365496 159752 395436 159780
rect 365496 159740 365502 159752
rect 395430 159740 395436 159752
rect 395488 159740 395494 159792
rect 396534 159740 396540 159792
rect 396592 159780 396598 159792
rect 413830 159780 413836 159792
rect 396592 159752 413836 159780
rect 396592 159740 396598 159752
rect 413830 159740 413836 159752
rect 413888 159740 413894 159792
rect 420914 159740 420920 159792
rect 420972 159780 420978 159792
rect 440418 159780 440424 159792
rect 420972 159752 440424 159780
rect 420972 159740 420978 159752
rect 440418 159740 440424 159752
rect 440476 159740 440482 159792
rect 453758 159740 453764 159792
rect 453816 159780 453822 159792
rect 464982 159780 464988 159792
rect 453816 159752 464988 159780
rect 453816 159740 453822 159752
rect 464982 159740 464988 159752
rect 465040 159740 465046 159792
rect 18874 159672 18880 159724
rect 18932 159712 18938 159724
rect 109126 159712 109132 159724
rect 18932 159684 109132 159712
rect 18932 159672 18938 159684
rect 109126 159672 109132 159684
rect 109184 159672 109190 159724
rect 113082 159672 113088 159724
rect 113140 159712 113146 159724
rect 126422 159712 126428 159724
rect 113140 159684 126428 159712
rect 113140 159672 113146 159684
rect 126422 159672 126428 159684
rect 126480 159672 126486 159724
rect 126514 159672 126520 159724
rect 126572 159712 126578 159724
rect 156506 159712 156512 159724
rect 126572 159684 156512 159712
rect 126572 159672 126578 159684
rect 156506 159672 156512 159684
rect 156564 159672 156570 159724
rect 164142 159712 164148 159724
rect 156800 159684 164148 159712
rect 49970 159604 49976 159656
rect 50028 159644 50034 159656
rect 143258 159644 143264 159656
rect 50028 159616 143264 159644
rect 50028 159604 50034 159616
rect 143258 159604 143264 159616
rect 143316 159604 143322 159656
rect 143350 159604 143356 159656
rect 143408 159644 143414 159656
rect 156598 159644 156604 159656
rect 143408 159616 156604 159644
rect 143408 159604 143414 159616
rect 156598 159604 156604 159616
rect 156656 159604 156662 159656
rect 43254 159536 43260 159588
rect 43312 159576 43318 159588
rect 136818 159576 136824 159588
rect 43312 159548 136824 159576
rect 43312 159536 43318 159548
rect 136818 159536 136824 159548
rect 136876 159536 136882 159588
rect 137278 159536 137284 159588
rect 137336 159576 137342 159588
rect 143994 159576 144000 159588
rect 137336 159548 144000 159576
rect 137336 159536 137342 159548
rect 143994 159536 144000 159548
rect 144052 159536 144058 159588
rect 144178 159536 144184 159588
rect 144236 159576 144242 159588
rect 144236 159548 147076 159576
rect 144236 159536 144242 159548
rect 36538 159468 36544 159520
rect 36596 159508 36602 159520
rect 36596 159480 126376 159508
rect 36596 159468 36602 159480
rect 32306 159400 32312 159452
rect 32364 159440 32370 159452
rect 126238 159440 126244 159452
rect 32364 159412 126244 159440
rect 32364 159400 32370 159412
rect 126238 159400 126244 159412
rect 126296 159400 126302 159452
rect 126348 159440 126376 159480
rect 126422 159468 126428 159520
rect 126480 159508 126486 159520
rect 127618 159508 127624 159520
rect 126480 159480 127624 159508
rect 126480 159468 126486 159480
rect 127618 159468 127624 159480
rect 127676 159468 127682 159520
rect 129918 159468 129924 159520
rect 129976 159508 129982 159520
rect 146754 159508 146760 159520
rect 129976 159480 146760 159508
rect 129976 159468 129982 159480
rect 146754 159468 146760 159480
rect 146812 159468 146818 159520
rect 147048 159508 147076 159548
rect 147214 159536 147220 159588
rect 147272 159576 147278 159588
rect 156800 159576 156828 159684
rect 164142 159672 164148 159684
rect 164200 159672 164206 159724
rect 167730 159672 167736 159724
rect 167788 159712 167794 159724
rect 246574 159712 246580 159724
rect 167788 159684 246580 159712
rect 167788 159672 167794 159684
rect 246574 159672 246580 159684
rect 246632 159672 246638 159724
rect 248506 159672 248512 159724
rect 248564 159712 248570 159724
rect 308122 159712 308128 159724
rect 248564 159684 308128 159712
rect 248564 159672 248570 159684
rect 308122 159672 308128 159684
rect 308180 159672 308186 159724
rect 308214 159672 308220 159724
rect 308272 159712 308278 159724
rect 308272 159684 342668 159712
rect 308272 159672 308278 159684
rect 161014 159604 161020 159656
rect 161072 159644 161078 159656
rect 241422 159644 241428 159656
rect 161072 159616 241428 159644
rect 161072 159604 161078 159616
rect 241422 159604 241428 159616
rect 241480 159604 241486 159656
rect 244274 159604 244280 159656
rect 244332 159644 244338 159656
rect 305178 159644 305184 159656
rect 244332 159616 305184 159644
rect 244332 159604 244338 159616
rect 305178 159604 305184 159616
rect 305236 159604 305242 159656
rect 309042 159604 309048 159656
rect 309100 159644 309106 159656
rect 342640 159644 342668 159684
rect 342714 159672 342720 159724
rect 342772 159712 342778 159724
rect 343818 159712 343824 159724
rect 342772 159684 343824 159712
rect 342772 159672 342778 159684
rect 343818 159672 343824 159684
rect 343876 159672 343882 159724
rect 347774 159672 347780 159724
rect 347832 159712 347838 159724
rect 378594 159712 378600 159724
rect 347832 159684 378600 159712
rect 347832 159672 347838 159684
rect 378594 159672 378600 159684
rect 378652 159672 378658 159724
rect 379698 159672 379704 159724
rect 379756 159712 379762 159724
rect 405918 159712 405924 159724
rect 379756 159684 405924 159712
rect 379756 159672 379762 159684
rect 405918 159672 405924 159684
rect 405976 159672 405982 159724
rect 414198 159672 414204 159724
rect 414256 159712 414262 159724
rect 434806 159712 434812 159724
rect 414256 159684 434812 159712
rect 414256 159672 414262 159684
rect 434806 159672 434812 159684
rect 434864 159672 434870 159724
rect 446122 159672 446128 159724
rect 446180 159712 446186 159724
rect 456794 159712 456800 159724
rect 446180 159684 456800 159712
rect 446180 159672 446186 159684
rect 456794 159672 456800 159684
rect 456852 159672 456858 159724
rect 458726 159672 458732 159724
rect 458784 159712 458790 159724
rect 465074 159712 465080 159724
rect 458784 159684 465080 159712
rect 458784 159672 458790 159684
rect 465074 159672 465080 159684
rect 465132 159672 465138 159724
rect 470502 159672 470508 159724
rect 470560 159712 470566 159724
rect 476114 159712 476120 159724
rect 470560 159684 476120 159712
rect 470560 159672 470566 159684
rect 476114 159672 476120 159684
rect 476172 159672 476178 159724
rect 478966 159672 478972 159724
rect 479024 159712 479030 159724
rect 484670 159712 484676 159724
rect 479024 159684 484676 159712
rect 479024 159672 479030 159684
rect 484670 159672 484676 159684
rect 484728 159672 484734 159724
rect 353386 159644 353392 159656
rect 309100 159616 342392 159644
rect 342640 159616 353392 159644
rect 309100 159604 309106 159616
rect 147272 159548 156828 159576
rect 147272 159536 147278 159548
rect 157610 159536 157616 159588
rect 157668 159576 157674 159588
rect 239122 159576 239128 159588
rect 157668 159548 239128 159576
rect 157668 159536 157674 159548
rect 239122 159536 239128 159548
rect 239180 159536 239186 159588
rect 250990 159536 250996 159588
rect 251048 159576 251054 159588
rect 310606 159576 310612 159588
rect 251048 159548 310612 159576
rect 251048 159536 251054 159548
rect 310606 159536 310612 159548
rect 310664 159536 310670 159588
rect 315758 159536 315764 159588
rect 315816 159576 315822 159588
rect 342254 159576 342260 159588
rect 315816 159548 342260 159576
rect 315816 159536 315822 159548
rect 342254 159536 342260 159548
rect 342312 159536 342318 159588
rect 147398 159508 147404 159520
rect 147048 159480 147404 159508
rect 147398 159468 147404 159480
rect 147456 159468 147462 159520
rect 225230 159508 225236 159520
rect 147508 159480 225236 159508
rect 129734 159440 129740 159452
rect 126348 159412 129740 159440
rect 129734 159400 129740 159412
rect 129792 159400 129798 159452
rect 130746 159400 130752 159452
rect 130804 159440 130810 159452
rect 137186 159440 137192 159452
rect 130804 159412 137192 159440
rect 130804 159400 130810 159412
rect 137186 159400 137192 159412
rect 137244 159400 137250 159452
rect 144178 159440 144184 159452
rect 137296 159412 144184 159440
rect 6270 159332 6276 159384
rect 6328 159372 6334 159384
rect 122834 159372 122840 159384
rect 6328 159344 122840 159372
rect 6328 159332 6334 159344
rect 122834 159332 122840 159344
rect 122892 159332 122898 159384
rect 123110 159332 123116 159384
rect 123168 159372 123174 159384
rect 137296 159372 137324 159412
rect 144178 159400 144184 159412
rect 144236 159400 144242 159452
rect 144362 159400 144368 159452
rect 144420 159440 144426 159452
rect 147508 159440 147536 159480
rect 225230 159468 225236 159480
rect 225288 159468 225294 159520
rect 231670 159468 231676 159520
rect 231728 159508 231734 159520
rect 295426 159508 295432 159520
rect 231728 159480 295432 159508
rect 231728 159468 231734 159480
rect 295426 159468 295432 159480
rect 295484 159468 295490 159520
rect 295610 159468 295616 159520
rect 295668 159508 295674 159520
rect 335814 159508 335820 159520
rect 295668 159480 335820 159508
rect 295668 159468 295674 159480
rect 335814 159468 335820 159480
rect 335872 159468 335878 159520
rect 335924 159480 336136 159508
rect 144420 159412 147536 159440
rect 144420 159400 144426 159412
rect 147582 159400 147588 159452
rect 147640 159440 147646 159452
rect 149330 159440 149336 159452
rect 147640 159412 149336 159440
rect 147640 159400 147646 159412
rect 149330 159400 149336 159412
rect 149388 159400 149394 159452
rect 150894 159400 150900 159452
rect 150952 159440 150958 159452
rect 233878 159440 233884 159452
rect 150952 159412 233884 159440
rect 150952 159400 150958 159412
rect 233878 159400 233884 159412
rect 233936 159400 233942 159452
rect 234982 159400 234988 159452
rect 235040 159440 235046 159452
rect 298002 159440 298008 159452
rect 235040 159412 298008 159440
rect 235040 159400 235046 159412
rect 298002 159400 298008 159412
rect 298060 159400 298066 159452
rect 301498 159400 301504 159452
rect 301556 159440 301562 159452
rect 335924 159440 335952 159480
rect 301556 159412 335952 159440
rect 336108 159440 336136 159480
rect 336182 159468 336188 159520
rect 336240 159508 336246 159520
rect 342364 159508 342392 159616
rect 353386 159604 353392 159616
rect 353444 159604 353450 159656
rect 357434 159604 357440 159656
rect 357492 159644 357498 159656
rect 363230 159644 363236 159656
rect 357492 159616 363236 159644
rect 357492 159604 357498 159616
rect 363230 159604 363236 159616
rect 363288 159604 363294 159656
rect 369578 159604 369584 159656
rect 369636 159644 369642 159656
rect 400674 159644 400680 159656
rect 369636 159616 400680 159644
rect 369636 159604 369642 159616
rect 400674 159604 400680 159616
rect 400732 159604 400738 159656
rect 407482 159604 407488 159656
rect 407540 159644 407546 159656
rect 429562 159644 429568 159656
rect 407540 159616 429568 159644
rect 407540 159604 407546 159616
rect 429562 159604 429568 159616
rect 429620 159604 429626 159656
rect 450354 159604 450360 159656
rect 450412 159644 450418 159656
rect 462222 159644 462228 159656
rect 450412 159616 462228 159644
rect 450412 159604 450418 159616
rect 462222 159604 462228 159616
rect 462280 159604 462286 159656
rect 468846 159604 468852 159656
rect 468904 159644 468910 159656
rect 474826 159644 474832 159656
rect 468904 159616 474832 159644
rect 468904 159604 468910 159616
rect 474826 159604 474832 159616
rect 474884 159604 474890 159656
rect 477310 159604 477316 159656
rect 477368 159644 477374 159656
rect 483290 159644 483296 159656
rect 477368 159616 483296 159644
rect 477368 159604 477374 159616
rect 483290 159604 483296 159616
rect 483348 159604 483354 159656
rect 342438 159536 342444 159588
rect 342496 159576 342502 159588
rect 359642 159576 359648 159588
rect 342496 159548 359648 159576
rect 342496 159536 342502 159548
rect 359642 159536 359648 159548
rect 359700 159536 359706 159588
rect 362862 159536 362868 159588
rect 362920 159576 362926 159588
rect 395246 159576 395252 159588
rect 362920 159548 395252 159576
rect 362920 159536 362926 159548
rect 395246 159536 395252 159548
rect 395304 159536 395310 159588
rect 399018 159536 399024 159588
rect 399076 159576 399082 159588
rect 408586 159576 408592 159588
rect 399076 159548 408592 159576
rect 399076 159536 399082 159548
rect 408586 159536 408592 159548
rect 408644 159536 408650 159588
rect 410794 159536 410800 159588
rect 410852 159576 410858 159588
rect 432138 159576 432144 159588
rect 410852 159548 432144 159576
rect 410852 159536 410858 159548
rect 432138 159536 432144 159548
rect 432196 159536 432202 159588
rect 451182 159536 451188 159588
rect 451240 159576 451246 159588
rect 461486 159576 461492 159588
rect 451240 159548 461492 159576
rect 451240 159536 451246 159548
rect 461486 159536 461492 159548
rect 461544 159536 461550 159588
rect 463786 159536 463792 159588
rect 463844 159576 463850 159588
rect 471514 159576 471520 159588
rect 463844 159548 471520 159576
rect 463844 159536 463850 159548
rect 471514 159536 471520 159548
rect 471572 159536 471578 159588
rect 479794 159536 479800 159588
rect 479852 159576 479858 159588
rect 484854 159576 484860 159588
rect 479852 159548 484860 159576
rect 479852 159536 479858 159548
rect 484854 159536 484860 159548
rect 484912 159536 484918 159588
rect 354766 159508 354772 159520
rect 336240 159480 341564 159508
rect 342364 159480 354772 159508
rect 336240 159468 336246 159480
rect 341426 159440 341432 159452
rect 336108 159412 341432 159440
rect 301556 159400 301562 159412
rect 341426 159400 341432 159412
rect 341484 159400 341490 159452
rect 341536 159440 341564 159480
rect 354766 159468 354772 159480
rect 354824 159468 354830 159520
rect 358630 159468 358636 159520
rect 358688 159508 358694 159520
rect 392394 159508 392400 159520
rect 358688 159480 392400 159508
rect 358688 159468 358694 159480
rect 392394 159468 392400 159480
rect 392452 159468 392458 159520
rect 424318 159468 424324 159520
rect 424376 159508 424382 159520
rect 442442 159508 442448 159520
rect 424376 159480 442448 159508
rect 424376 159468 424382 159480
rect 442442 159468 442448 159480
rect 442500 159468 442506 159520
rect 452010 159468 452016 159520
rect 452068 159508 452074 159520
rect 463602 159508 463608 159520
rect 452068 159480 463608 159508
rect 452068 159468 452074 159480
rect 463602 159468 463608 159480
rect 463660 159468 463666 159520
rect 465534 159468 465540 159520
rect 465592 159508 465598 159520
rect 472250 159508 472256 159520
rect 465592 159480 472256 159508
rect 465592 159468 465598 159480
rect 472250 159468 472256 159480
rect 472308 159468 472314 159520
rect 343450 159440 343456 159452
rect 341536 159412 343456 159440
rect 343450 159400 343456 159412
rect 343508 159400 343514 159452
rect 348786 159440 348792 159452
rect 345952 159412 348792 159440
rect 123168 159344 137324 159372
rect 123168 159332 123174 159344
rect 137462 159332 137468 159384
rect 137520 159372 137526 159384
rect 223574 159372 223580 159384
rect 137520 159344 223580 159372
rect 137520 159332 137526 159344
rect 223574 159332 223580 159344
rect 223632 159332 223638 159384
rect 224954 159332 224960 159384
rect 225012 159372 225018 159384
rect 290274 159372 290280 159384
rect 225012 159344 290280 159372
rect 225012 159332 225018 159344
rect 290274 159332 290280 159344
rect 290332 159332 290338 159384
rect 294782 159332 294788 159384
rect 294840 159372 294846 159384
rect 335998 159372 336004 159384
rect 294840 159344 336004 159372
rect 294840 159332 294846 159344
rect 335998 159332 336004 159344
rect 336056 159332 336062 159384
rect 336090 159332 336096 159384
rect 336148 159372 336154 159384
rect 342254 159372 342260 159384
rect 336148 159344 342260 159372
rect 336148 159332 336154 159344
rect 342254 159332 342260 159344
rect 342312 159332 342318 159384
rect 342346 159332 342352 159384
rect 342404 159372 342410 159384
rect 345952 159372 345980 159412
rect 348786 159400 348792 159412
rect 348844 159400 348850 159452
rect 356146 159400 356152 159452
rect 356204 159440 356210 159452
rect 390554 159440 390560 159452
rect 356204 159412 390560 159440
rect 356204 159400 356210 159412
rect 390554 159400 390560 159412
rect 390612 159400 390618 159452
rect 404078 159400 404084 159452
rect 404136 159440 404142 159452
rect 426986 159440 426992 159452
rect 404136 159412 426992 159440
rect 404136 159400 404142 159412
rect 426986 159400 426992 159412
rect 427044 159400 427050 159452
rect 427630 159400 427636 159452
rect 427688 159440 427694 159452
rect 445018 159440 445024 159452
rect 427688 159412 445024 159440
rect 427688 159400 427694 159412
rect 445018 159400 445024 159412
rect 445076 159400 445082 159452
rect 447870 159400 447876 159452
rect 447928 159440 447934 159452
rect 460106 159440 460112 159452
rect 447928 159412 460112 159440
rect 447928 159400 447934 159412
rect 460106 159400 460112 159412
rect 460164 159400 460170 159452
rect 518342 159400 518348 159452
rect 518400 159440 518406 159452
rect 523494 159440 523500 159452
rect 518400 159412 523500 159440
rect 518400 159400 518406 159412
rect 523494 159400 523500 159412
rect 523552 159400 523558 159452
rect 342404 159344 345980 159372
rect 342404 159332 342410 159344
rect 346026 159332 346032 159384
rect 346084 159372 346090 159384
rect 382734 159372 382740 159384
rect 346084 159344 382740 159372
rect 346084 159332 346090 159344
rect 382734 159332 382740 159344
rect 382792 159332 382798 159384
rect 383102 159332 383108 159384
rect 383160 159372 383166 159384
rect 411346 159372 411352 159384
rect 383160 159344 411352 159372
rect 383160 159332 383166 159344
rect 411346 159332 411352 159344
rect 411404 159332 411410 159384
rect 417510 159332 417516 159384
rect 417568 159372 417574 159384
rect 437658 159372 437664 159384
rect 417568 159344 437664 159372
rect 417568 159332 417574 159344
rect 437658 159332 437664 159344
rect 437716 159332 437722 159384
rect 448698 159332 448704 159384
rect 448756 159372 448762 159384
rect 461210 159372 461216 159384
rect 448756 159344 461216 159372
rect 448756 159332 448762 159344
rect 461210 159332 461216 159344
rect 461268 159332 461274 159384
rect 461302 159332 461308 159384
rect 461360 159372 461366 159384
rect 468018 159372 468024 159384
rect 461360 159344 468024 159372
rect 461360 159332 461366 159344
rect 468018 159332 468024 159344
rect 468076 159332 468082 159384
rect 469674 159332 469680 159384
rect 469732 159372 469738 159384
rect 477402 159372 477408 159384
rect 469732 159344 477408 159372
rect 469732 159332 469738 159344
rect 477402 159332 477408 159344
rect 477460 159332 477466 159384
rect 478138 159332 478144 159384
rect 478196 159372 478202 159384
rect 483658 159372 483664 159384
rect 478196 159344 483664 159372
rect 478196 159332 478202 159344
rect 483658 159332 483664 159344
rect 483716 159332 483722 159384
rect 517606 159332 517612 159384
rect 517664 159372 517670 159384
rect 522666 159372 522672 159384
rect 517664 159344 522672 159372
rect 517664 159332 517670 159344
rect 522666 159332 522672 159344
rect 522724 159332 522730 159384
rect 73522 159264 73528 159316
rect 73580 159304 73586 159316
rect 80054 159304 80060 159316
rect 73580 159276 80060 159304
rect 73580 159264 73586 159276
rect 80054 159264 80060 159276
rect 80112 159264 80118 159316
rect 83642 159264 83648 159316
rect 83700 159304 83706 159316
rect 166994 159304 167000 159316
rect 83700 159276 167000 159304
rect 83700 159264 83706 159276
rect 166994 159264 167000 159276
rect 167052 159264 167058 159316
rect 170214 159264 170220 159316
rect 170272 159304 170278 159316
rect 198918 159304 198924 159316
rect 170272 159276 198924 159304
rect 170272 159264 170278 159276
rect 198918 159264 198924 159276
rect 198976 159264 198982 159316
rect 201402 159264 201408 159316
rect 201460 159304 201466 159316
rect 212626 159304 212632 159316
rect 201460 159276 212632 159304
rect 201460 159264 201466 159276
rect 212626 159264 212632 159276
rect 212684 159264 212690 159316
rect 214006 159264 214012 159316
rect 214064 159304 214070 159316
rect 281994 159304 282000 159316
rect 214064 159276 282000 159304
rect 214064 159264 214070 159276
rect 281994 159264 282000 159276
rect 282052 159264 282058 159316
rect 282086 159264 282092 159316
rect 282144 159304 282150 159316
rect 333974 159304 333980 159316
rect 282144 159276 333980 159304
rect 282144 159264 282150 159276
rect 333974 159264 333980 159276
rect 334032 159264 334038 159316
rect 334250 159264 334256 159316
rect 334308 159304 334314 159316
rect 373994 159304 374000 159316
rect 334308 159276 374000 159304
rect 334308 159264 334314 159276
rect 373994 159264 374000 159276
rect 374052 159264 374058 159316
rect 388990 159264 388996 159316
rect 389048 159304 389054 159316
rect 404170 159304 404176 159316
rect 389048 159276 404176 159304
rect 389048 159264 389054 159276
rect 404170 159264 404176 159276
rect 404228 159264 404234 159316
rect 457898 159264 457904 159316
rect 457956 159304 457962 159316
rect 468110 159304 468116 159316
rect 457956 159276 468116 159304
rect 457956 159264 457962 159276
rect 468110 159264 468116 159276
rect 468168 159264 468174 159316
rect 80238 159196 80244 159248
rect 80296 159236 80302 159248
rect 91094 159236 91100 159248
rect 80296 159208 91100 159236
rect 80296 159196 80302 159208
rect 91094 159196 91100 159208
rect 91152 159196 91158 159248
rect 100478 159196 100484 159248
rect 100536 159236 100542 159248
rect 184658 159236 184664 159248
rect 100536 159208 184664 159236
rect 100536 159196 100542 159208
rect 184658 159196 184664 159208
rect 184716 159196 184722 159248
rect 187050 159196 187056 159248
rect 187108 159236 187114 159248
rect 214650 159236 214656 159248
rect 187108 159208 214656 159236
rect 187108 159196 187114 159208
rect 214650 159196 214656 159208
rect 214708 159196 214714 159248
rect 218238 159196 218244 159248
rect 218296 159236 218302 159248
rect 285122 159236 285128 159248
rect 218296 159208 285128 159236
rect 218296 159196 218302 159208
rect 285122 159196 285128 159208
rect 285180 159196 285186 159248
rect 287974 159196 287980 159248
rect 288032 159236 288038 159248
rect 338390 159236 338396 159248
rect 288032 159208 338396 159236
rect 288032 159196 288038 159208
rect 338390 159196 338396 159208
rect 338448 159196 338454 159248
rect 339310 159196 339316 159248
rect 339368 159236 339374 159248
rect 377582 159236 377588 159248
rect 339368 159208 377588 159236
rect 339368 159196 339374 159208
rect 377582 159196 377588 159208
rect 377640 159196 377646 159248
rect 385586 159196 385592 159248
rect 385644 159236 385650 159248
rect 398926 159236 398932 159248
rect 385644 159208 398932 159236
rect 385644 159196 385650 159208
rect 398926 159196 398932 159208
rect 398984 159196 398990 159248
rect 400766 159196 400772 159248
rect 400824 159236 400830 159248
rect 424502 159236 424508 159248
rect 400824 159208 424508 159236
rect 400824 159196 400830 159208
rect 424502 159196 424508 159208
rect 424560 159196 424566 159248
rect 457070 159196 457076 159248
rect 457128 159236 457134 159248
rect 467834 159236 467840 159248
rect 457128 159208 467840 159236
rect 457128 159196 457134 159208
rect 467834 159196 467840 159208
rect 467892 159196 467898 159248
rect 86954 159128 86960 159180
rect 87012 159168 87018 159180
rect 87012 159140 162992 159168
rect 87012 159128 87018 159140
rect 93670 159060 93676 159112
rect 93728 159100 93734 159112
rect 162854 159100 162860 159112
rect 93728 159072 162860 159100
rect 93728 159060 93734 159072
rect 162854 159060 162860 159072
rect 162912 159060 162918 159112
rect 162964 159100 162992 159140
rect 163038 159128 163044 159180
rect 163096 159168 163102 159180
rect 172422 159168 172428 159180
rect 163096 159140 172428 159168
rect 163096 159128 163102 159140
rect 172422 159128 172428 159140
rect 172480 159128 172486 159180
rect 193766 159128 193772 159180
rect 193824 159168 193830 159180
rect 218054 159168 218060 159180
rect 193824 159140 218060 159168
rect 193824 159128 193830 159140
rect 218054 159128 218060 159140
rect 218112 159128 218118 159180
rect 220722 159128 220728 159180
rect 220780 159168 220786 159180
rect 283190 159168 283196 159180
rect 220780 159140 283196 159168
rect 220780 159128 220786 159140
rect 283190 159128 283196 159140
rect 283248 159128 283254 159180
rect 284662 159128 284668 159180
rect 284720 159168 284726 159180
rect 285766 159168 285772 159180
rect 284720 159140 285772 159168
rect 284720 159128 284726 159140
rect 285766 159128 285772 159140
rect 285824 159128 285830 159180
rect 288158 159168 288164 159180
rect 287026 159140 288164 159168
rect 169846 159100 169852 159112
rect 162964 159072 169852 159100
rect 169846 159060 169852 159072
rect 169904 159060 169910 159112
rect 171134 159060 171140 159112
rect 171192 159100 171198 159112
rect 172698 159100 172704 159112
rect 171192 159072 172704 159100
rect 171192 159060 171198 159072
rect 172698 159060 172704 159072
rect 172756 159060 172762 159112
rect 173618 159060 173624 159112
rect 173676 159100 173682 159112
rect 197354 159100 197360 159112
rect 173676 159072 197360 159100
rect 173676 159060 173682 159072
rect 197354 159060 197360 159072
rect 197412 159060 197418 159112
rect 224126 159060 224132 159112
rect 224184 159100 224190 159112
rect 287026 159100 287054 159140
rect 288158 159128 288164 159140
rect 288216 159128 288222 159180
rect 288894 159128 288900 159180
rect 288952 159168 288958 159180
rect 339034 159168 339040 159180
rect 288952 159140 339040 159168
rect 288952 159128 288958 159140
rect 339034 159128 339040 159140
rect 339092 159128 339098 159180
rect 341426 159128 341432 159180
rect 341484 159168 341490 159180
rect 348694 159168 348700 159180
rect 341484 159140 348700 159168
rect 341484 159128 341490 159140
rect 348694 159128 348700 159140
rect 348752 159128 348758 159180
rect 348786 159128 348792 159180
rect 348844 159168 348850 159180
rect 374086 159168 374092 159180
rect 348844 159140 374092 159168
rect 348844 159128 348850 159140
rect 374086 159128 374092 159140
rect 374144 159128 374150 159180
rect 385402 159168 385408 159180
rect 377968 159140 385408 159168
rect 224184 159072 287054 159100
rect 224184 159060 224190 159072
rect 302326 159060 302332 159112
rect 302384 159100 302390 159112
rect 349246 159100 349252 159112
rect 302384 159072 349252 159100
rect 302384 159060 302390 159072
rect 349246 159060 349252 159072
rect 349304 159060 349310 159112
rect 351822 159100 351828 159112
rect 350506 159072 351828 159100
rect 107194 158992 107200 159044
rect 107252 159032 107258 159044
rect 182542 159032 182548 159044
rect 107252 159004 182548 159032
rect 107252 158992 107258 159004
rect 182542 158992 182548 159004
rect 182600 158992 182606 159044
rect 183738 158992 183744 159044
rect 183796 159032 183802 159044
rect 200482 159032 200488 159044
rect 183796 159004 200488 159032
rect 183796 158992 183802 159004
rect 200482 158992 200488 159004
rect 200540 158992 200546 159044
rect 200574 158992 200580 159044
rect 200632 159032 200638 159044
rect 224954 159032 224960 159044
rect 200632 159004 224960 159032
rect 200632 158992 200638 159004
rect 224954 158992 224960 159004
rect 225012 158992 225018 159044
rect 230842 158992 230848 159044
rect 230900 159032 230906 159044
rect 294782 159032 294788 159044
rect 230900 159004 294788 159032
rect 230900 158992 230906 159004
rect 294782 158992 294788 159004
rect 294840 158992 294846 159044
rect 298094 158992 298100 159044
rect 298152 159032 298158 159044
rect 299658 159032 299664 159044
rect 298152 159004 299664 159032
rect 298152 158992 298158 159004
rect 299658 158992 299664 159004
rect 299716 158992 299722 159044
rect 307386 158992 307392 159044
rect 307444 159032 307450 159044
rect 350506 159032 350534 159072
rect 351822 159060 351828 159072
rect 351880 159060 351886 159112
rect 351914 159060 351920 159112
rect 351972 159100 351978 159112
rect 377968 159100 377996 159140
rect 385402 159128 385408 159140
rect 385460 159128 385466 159180
rect 392302 159128 392308 159180
rect 392360 159168 392366 159180
rect 404262 159168 404268 159180
rect 392360 159140 404268 159168
rect 392360 159128 392366 159140
rect 404262 159128 404268 159140
rect 404320 159128 404326 159180
rect 456242 159128 456248 159180
rect 456300 159168 456306 159180
rect 466914 159168 466920 159180
rect 456300 159140 466920 159168
rect 456300 159128 456306 159140
rect 466914 159128 466920 159140
rect 466972 159128 466978 159180
rect 351972 159072 377996 159100
rect 351972 159060 351978 159072
rect 378042 159060 378048 159112
rect 378100 159100 378106 159112
rect 388438 159100 388444 159112
rect 378100 159072 388444 159100
rect 378100 159060 378106 159072
rect 388438 159060 388444 159072
rect 388496 159060 388502 159112
rect 395706 159060 395712 159112
rect 395764 159100 395770 159112
rect 405458 159100 405464 159112
rect 395764 159072 405464 159100
rect 395764 159060 395770 159072
rect 405458 159060 405464 159072
rect 405516 159060 405522 159112
rect 460474 159060 460480 159112
rect 460532 159100 460538 159112
rect 466546 159100 466552 159112
rect 460532 159072 466552 159100
rect 460532 159060 460538 159072
rect 466546 159060 466552 159072
rect 466604 159060 466610 159112
rect 471422 159060 471428 159112
rect 471480 159100 471486 159112
rect 478414 159100 478420 159112
rect 471480 159072 478420 159100
rect 471480 159060 471486 159072
rect 478414 159060 478420 159072
rect 478472 159060 478478 159112
rect 307444 159004 350534 159032
rect 307444 158992 307450 159004
rect 351086 158992 351092 159044
rect 351144 159032 351150 159044
rect 382366 159032 382372 159044
rect 351144 159004 382372 159032
rect 351144 158992 351150 159004
rect 382366 158992 382372 159004
rect 382424 158992 382430 159044
rect 459646 158992 459652 159044
rect 459704 159032 459710 159044
rect 466454 159032 466460 159044
rect 459704 159004 466460 159032
rect 459704 158992 459710 159004
rect 466454 158992 466460 159004
rect 466512 158992 466518 159044
rect 473906 158992 473912 159044
rect 473964 159032 473970 159044
rect 480346 159032 480352 159044
rect 473964 159004 480352 159032
rect 473964 158992 473970 159004
rect 480346 158992 480352 159004
rect 480404 158992 480410 159044
rect 480622 158992 480628 159044
rect 480680 159032 480686 159044
rect 485958 159032 485964 159044
rect 480680 159004 485964 159032
rect 480680 158992 480686 159004
rect 485958 158992 485964 159004
rect 486016 158992 486022 159044
rect 96246 158924 96252 158976
rect 96304 158964 96310 158976
rect 121638 158964 121644 158976
rect 96304 158936 121644 158964
rect 96304 158924 96310 158936
rect 121638 158924 121644 158936
rect 121696 158924 121702 158976
rect 124030 158924 124036 158976
rect 124088 158964 124094 158976
rect 193398 158964 193404 158976
rect 124088 158936 193404 158964
rect 124088 158924 124094 158936
rect 193398 158924 193404 158936
rect 193456 158924 193462 158976
rect 194686 158924 194692 158976
rect 194744 158964 194750 158976
rect 203702 158964 203708 158976
rect 194744 158936 203708 158964
rect 194744 158924 194750 158936
rect 203702 158924 203708 158936
rect 203760 158924 203766 158976
rect 207290 158924 207296 158976
rect 207348 158964 207354 158976
rect 230750 158964 230756 158976
rect 207348 158936 230756 158964
rect 207348 158924 207354 158936
rect 230750 158924 230756 158936
rect 230808 158924 230814 158976
rect 237558 158924 237564 158976
rect 237616 158964 237622 158976
rect 299474 158964 299480 158976
rect 237616 158936 299480 158964
rect 237616 158924 237622 158936
rect 299474 158924 299480 158936
rect 299532 158924 299538 158976
rect 314930 158924 314936 158976
rect 314988 158964 314994 158976
rect 357526 158964 357532 158976
rect 314988 158936 357532 158964
rect 314988 158924 314994 158936
rect 357526 158924 357532 158936
rect 357584 158924 357590 158976
rect 357802 158924 357808 158976
rect 357860 158964 357866 158976
rect 384942 158964 384948 158976
rect 357860 158936 384948 158964
rect 357860 158924 357866 158936
rect 384942 158924 384948 158936
rect 385000 158924 385006 158976
rect 409138 158924 409144 158976
rect 409196 158964 409202 158976
rect 410886 158964 410892 158976
rect 409196 158936 410892 158964
rect 409196 158924 409202 158936
rect 410886 158924 410892 158936
rect 410944 158924 410950 158976
rect 413370 158924 413376 158976
rect 413428 158964 413434 158976
rect 419718 158964 419724 158976
rect 413428 158936 419724 158964
rect 413428 158924 413434 158936
rect 419718 158924 419724 158936
rect 419776 158924 419782 158976
rect 462130 158924 462136 158976
rect 462188 158964 462194 158976
rect 467926 158964 467932 158976
rect 462188 158936 467932 158964
rect 462188 158924 462194 158936
rect 467926 158924 467932 158936
rect 467984 158924 467990 158976
rect 475562 158924 475568 158976
rect 475620 158964 475626 158976
rect 481726 158964 481732 158976
rect 475620 158936 481732 158964
rect 475620 158924 475626 158936
rect 481726 158924 481732 158936
rect 481784 158924 481790 158976
rect 506658 158924 506664 158976
rect 506716 158964 506722 158976
rect 508406 158964 508412 158976
rect 506716 158936 508412 158964
rect 506716 158924 506722 158936
rect 508406 158924 508412 158936
rect 508464 158924 508470 158976
rect 102962 158856 102968 158908
rect 103020 158896 103026 158908
rect 125502 158896 125508 158908
rect 103020 158868 125508 158896
rect 103020 158856 103026 158868
rect 125502 158856 125508 158868
rect 125560 158856 125566 158908
rect 137094 158896 137100 158908
rect 133156 158868 137100 158896
rect 109678 158788 109684 158840
rect 109736 158828 109742 158840
rect 133156 158828 133184 158868
rect 137094 158856 137100 158868
rect 137152 158856 137158 158908
rect 137186 158856 137192 158908
rect 137244 158896 137250 158908
rect 195422 158896 195428 158908
rect 137244 158868 195428 158896
rect 137244 158856 137250 158868
rect 195422 158856 195428 158868
rect 195480 158856 195486 158908
rect 208118 158856 208124 158908
rect 208176 158896 208182 158908
rect 212442 158896 212448 158908
rect 208176 158868 212448 158896
rect 208176 158856 208182 158868
rect 212442 158856 212448 158868
rect 212500 158856 212506 158908
rect 217318 158856 217324 158908
rect 217376 158896 217382 158908
rect 220722 158896 220728 158908
rect 217376 158868 220728 158896
rect 217376 158856 217382 158868
rect 220722 158856 220728 158868
rect 220780 158856 220786 158908
rect 241790 158856 241796 158908
rect 241848 158896 241854 158908
rect 303246 158896 303252 158908
rect 241848 158868 303252 158896
rect 241848 158856 241854 158868
rect 303246 158856 303252 158868
rect 303304 158856 303310 158908
rect 305638 158856 305644 158908
rect 305696 158896 305702 158908
rect 307386 158896 307392 158908
rect 305696 158868 307392 158896
rect 305696 158856 305702 158868
rect 307386 158856 307392 158868
rect 307444 158856 307450 158908
rect 310698 158856 310704 158908
rect 310756 158896 310762 158908
rect 311986 158896 311992 158908
rect 310756 158868 311992 158896
rect 310756 158856 310762 158868
rect 311986 158856 311992 158868
rect 312044 158856 312050 158908
rect 312354 158856 312360 158908
rect 312412 158896 312418 158908
rect 318794 158896 318800 158908
rect 312412 158868 318800 158896
rect 312412 158856 312418 158868
rect 318794 158856 318800 158868
rect 318852 158856 318858 158908
rect 320818 158856 320824 158908
rect 320876 158896 320882 158908
rect 320876 158868 357572 158896
rect 320876 158856 320882 158868
rect 109736 158800 133184 158828
rect 109736 158788 109742 158800
rect 133230 158788 133236 158840
rect 133288 158828 133294 158840
rect 158714 158828 158720 158840
rect 133288 158800 158720 158828
rect 133288 158788 133294 158800
rect 158714 158788 158720 158800
rect 158772 158788 158778 158840
rect 163498 158788 163504 158840
rect 163556 158828 163562 158840
rect 197262 158828 197268 158840
rect 163556 158800 197268 158828
rect 163556 158788 163562 158800
rect 197262 158788 197268 158800
rect 197320 158788 197326 158840
rect 203886 158788 203892 158840
rect 203944 158828 203950 158840
rect 213638 158828 213644 158840
rect 203944 158800 213644 158828
rect 203944 158788 203950 158800
rect 213638 158788 213644 158800
rect 213696 158788 213702 158840
rect 214834 158788 214840 158840
rect 214892 158828 214898 158840
rect 222102 158828 222108 158840
rect 214892 158800 222108 158828
rect 214892 158788 214898 158800
rect 222102 158788 222108 158800
rect 222160 158788 222166 158840
rect 238386 158788 238392 158840
rect 238444 158828 238450 158840
rect 241606 158828 241612 158840
rect 238444 158800 241612 158828
rect 238444 158788 238450 158800
rect 241606 158788 241612 158800
rect 241664 158788 241670 158840
rect 261110 158788 261116 158840
rect 261168 158828 261174 158840
rect 316310 158828 316316 158840
rect 261168 158800 316316 158828
rect 261168 158788 261174 158800
rect 316310 158788 316316 158800
rect 316368 158788 316374 158840
rect 319162 158788 319168 158840
rect 319220 158828 319226 158840
rect 319220 158800 321600 158828
rect 319220 158788 319226 158800
rect 90358 158720 90364 158772
rect 90416 158760 90422 158772
rect 92566 158760 92572 158772
rect 90416 158732 92572 158760
rect 90416 158720 90422 158732
rect 92566 158720 92572 158732
rect 92624 158720 92630 158772
rect 92842 158720 92848 158772
rect 92900 158760 92906 158772
rect 114462 158760 114468 158772
rect 92900 158732 114468 158760
rect 92900 158720 92906 158732
rect 114462 158720 114468 158732
rect 114520 158720 114526 158772
rect 119798 158720 119804 158772
rect 119856 158760 119862 158772
rect 146570 158760 146576 158772
rect 119856 158732 146576 158760
rect 119856 158720 119862 158732
rect 146570 158720 146576 158732
rect 146628 158720 146634 158772
rect 146662 158720 146668 158772
rect 146720 158760 146726 158772
rect 176654 158760 176660 158772
rect 146720 158732 176660 158760
rect 146720 158720 146726 158732
rect 176654 158720 176660 158732
rect 176712 158720 176718 158772
rect 180334 158720 180340 158772
rect 180392 158760 180398 158772
rect 204898 158760 204904 158772
rect 180392 158732 204904 158760
rect 180392 158720 180398 158732
rect 204898 158720 204904 158732
rect 204956 158720 204962 158772
rect 210602 158720 210608 158772
rect 210660 158760 210666 158772
rect 215386 158760 215392 158772
rect 210660 158732 215392 158760
rect 210660 158720 210666 158732
rect 215386 158720 215392 158732
rect 215444 158720 215450 158772
rect 221550 158720 221556 158772
rect 221608 158760 221614 158772
rect 224034 158760 224040 158772
rect 221608 158732 224040 158760
rect 221608 158720 221614 158732
rect 224034 158720 224040 158732
rect 224092 158720 224098 158772
rect 240870 158720 240876 158772
rect 240928 158760 240934 158772
rect 243354 158760 243360 158772
rect 240928 158732 243360 158760
rect 240928 158720 240934 158732
rect 243354 158720 243360 158732
rect 243412 158720 243418 158772
rect 254394 158720 254400 158772
rect 254452 158760 254458 158772
rect 255406 158760 255412 158772
rect 254452 158732 255412 158760
rect 254452 158720 254458 158732
rect 255406 158720 255412 158732
rect 255464 158720 255470 158772
rect 258534 158720 258540 158772
rect 258592 158760 258598 158772
rect 260834 158760 260840 158772
rect 258592 158732 260840 158760
rect 258592 158720 258598 158732
rect 260834 158720 260840 158732
rect 260892 158720 260898 158772
rect 264422 158720 264428 158772
rect 264480 158760 264486 158772
rect 266354 158760 266360 158772
rect 264480 158732 266360 158760
rect 264480 158720 264486 158732
rect 266354 158720 266360 158732
rect 266412 158720 266418 158772
rect 267826 158720 267832 158772
rect 267884 158760 267890 158772
rect 320266 158760 320272 158772
rect 267884 158732 320272 158760
rect 267884 158720 267890 158732
rect 320266 158720 320272 158732
rect 320324 158720 320330 158772
rect 321572 158704 321600 158800
rect 321646 158788 321652 158840
rect 321704 158828 321710 158840
rect 357434 158828 357440 158840
rect 321704 158800 357440 158828
rect 321704 158788 321710 158800
rect 357434 158788 357440 158800
rect 357492 158788 357498 158840
rect 357544 158828 357572 158868
rect 361206 158856 361212 158908
rect 361264 158896 361270 158908
rect 385126 158896 385132 158908
rect 361264 158868 385132 158896
rect 361264 158856 361270 158868
rect 385126 158856 385132 158868
rect 385184 158856 385190 158908
rect 391474 158856 391480 158908
rect 391532 158896 391538 158908
rect 394602 158896 394608 158908
rect 391532 158868 394608 158896
rect 391532 158856 391538 158868
rect 394602 158856 394608 158868
rect 394660 158856 394666 158908
rect 412542 158856 412548 158908
rect 412600 158896 412606 158908
rect 413094 158896 413100 158908
rect 412600 158868 413100 158896
rect 412600 158856 412606 158868
rect 413094 158856 413100 158868
rect 413152 158856 413158 158908
rect 420086 158856 420092 158908
rect 420144 158896 420150 158908
rect 423582 158896 423588 158908
rect 420144 158868 423588 158896
rect 420144 158856 420150 158868
rect 423582 158856 423588 158868
rect 423640 158856 423646 158908
rect 462958 158856 462964 158908
rect 463016 158896 463022 158908
rect 469214 158896 469220 158908
rect 463016 158868 469220 158896
rect 463016 158856 463022 158868
rect 469214 158856 469220 158868
rect 469272 158856 469278 158908
rect 474734 158856 474740 158908
rect 474792 158896 474798 158908
rect 481082 158896 481088 158908
rect 474792 158868 481088 158896
rect 474792 158856 474798 158868
rect 481082 158856 481088 158868
rect 481140 158856 481146 158908
rect 482278 158856 482284 158908
rect 482336 158896 482342 158908
rect 487246 158896 487252 158908
rect 482336 158868 487252 158896
rect 482336 158856 482342 158868
rect 487246 158856 487252 158868
rect 487304 158856 487310 158908
rect 507946 158856 507952 158908
rect 508004 158896 508010 158908
rect 510062 158896 510068 158908
rect 508004 158868 510068 158896
rect 508004 158856 508010 158868
rect 510062 158856 510068 158868
rect 510120 158856 510126 158908
rect 362954 158828 362960 158840
rect 357544 158800 362960 158828
rect 362954 158788 362960 158800
rect 363012 158788 363018 158840
rect 367922 158788 367928 158840
rect 367980 158828 367986 158840
rect 386322 158828 386328 158840
rect 367980 158800 373994 158828
rect 367980 158788 367986 158800
rect 327534 158720 327540 158772
rect 327592 158760 327598 158772
rect 368382 158760 368388 158772
rect 327592 158732 368388 158760
rect 327592 158720 327598 158732
rect 368382 158720 368388 158732
rect 368440 158720 368446 158772
rect 373966 158760 373994 158800
rect 374104 158800 386328 158828
rect 374104 158760 374132 158800
rect 386322 158788 386328 158800
rect 386380 158788 386386 158840
rect 389174 158828 389180 158840
rect 386984 158800 389180 158828
rect 373966 158732 374132 158760
rect 374178 158720 374184 158772
rect 374236 158760 374242 158772
rect 379422 158760 379428 158772
rect 374236 158732 379428 158760
rect 374236 158720 374242 158732
rect 379422 158720 379428 158732
rect 379480 158720 379486 158772
rect 384758 158720 384764 158772
rect 384816 158760 384822 158772
rect 386984 158760 387012 158800
rect 389174 158788 389180 158800
rect 389232 158788 389238 158840
rect 405734 158788 405740 158840
rect 405792 158828 405798 158840
rect 409230 158828 409236 158840
rect 405792 158800 409236 158828
rect 405792 158788 405798 158800
rect 409230 158788 409236 158800
rect 409288 158788 409294 158840
rect 416682 158788 416688 158840
rect 416740 158828 416746 158840
rect 419626 158828 419632 158840
rect 416740 158800 419632 158828
rect 416740 158788 416746 158800
rect 419626 158788 419632 158800
rect 419684 158788 419690 158840
rect 466362 158788 466368 158840
rect 466420 158828 466426 158840
rect 472434 158828 472440 158840
rect 466420 158800 472440 158828
rect 466420 158788 466426 158800
rect 472434 158788 472440 158800
rect 472492 158788 472498 158840
rect 476390 158788 476396 158840
rect 476448 158828 476454 158840
rect 482370 158828 482376 158840
rect 476448 158800 482376 158828
rect 476448 158788 476454 158800
rect 482370 158788 482376 158800
rect 482428 158788 482434 158840
rect 506106 158788 506112 158840
rect 506164 158828 506170 158840
rect 507578 158828 507584 158840
rect 506164 158800 507584 158828
rect 506164 158788 506170 158800
rect 507578 158788 507584 158800
rect 507636 158788 507642 158840
rect 384816 158732 387012 158760
rect 384816 158720 384822 158732
rect 388070 158720 388076 158772
rect 388128 158760 388134 158772
rect 390370 158760 390376 158772
rect 388128 158732 390376 158760
rect 388128 158720 388134 158732
rect 390370 158720 390376 158732
rect 390428 158720 390434 158772
rect 464614 158720 464620 158772
rect 464672 158760 464678 158772
rect 471238 158760 471244 158772
rect 464672 158732 471244 158760
rect 464672 158720 464678 158732
rect 471238 158720 471244 158732
rect 471296 158720 471302 158772
rect 473078 158720 473084 158772
rect 473136 158760 473142 158772
rect 479702 158760 479708 158772
rect 473136 158732 479708 158760
rect 473136 158720 473142 158732
rect 479702 158720 479708 158732
rect 479760 158720 479766 158772
rect 481450 158720 481456 158772
rect 481508 158760 481514 158772
rect 486142 158760 486148 158772
rect 481508 158732 486148 158760
rect 481508 158720 481514 158732
rect 486142 158720 486148 158732
rect 486200 158720 486206 158772
rect 505370 158720 505376 158772
rect 505428 158760 505434 158772
rect 506750 158760 506756 158772
rect 505428 158732 506756 158760
rect 505428 158720 505434 158732
rect 506750 158720 506756 158732
rect 506808 158720 506814 158772
rect 509326 158720 509332 158772
rect 509384 158760 509390 158772
rect 511718 158760 511724 158772
rect 509384 158732 511724 158760
rect 509384 158720 509390 158732
rect 511718 158720 511724 158732
rect 511776 158720 511782 158772
rect 514938 158720 514944 158772
rect 514996 158760 515002 158772
rect 518526 158760 518532 158772
rect 514996 158732 518532 158760
rect 514996 158720 515002 158732
rect 518526 158720 518532 158732
rect 518584 158720 518590 158772
rect 81066 158652 81072 158704
rect 81124 158692 81130 158704
rect 180886 158692 180892 158704
rect 81124 158664 180892 158692
rect 81124 158652 81130 158664
rect 180886 158652 180892 158664
rect 180944 158652 180950 158704
rect 181990 158652 181996 158704
rect 182048 158692 182054 158704
rect 257522 158692 257528 158704
rect 182048 158664 257528 158692
rect 182048 158652 182054 158664
rect 257522 158652 257528 158664
rect 257580 158652 257586 158704
rect 321554 158652 321560 158704
rect 321612 158652 321618 158704
rect 67634 158584 67640 158636
rect 67692 158624 67698 158636
rect 170214 158624 170220 158636
rect 67692 158596 170220 158624
rect 67692 158584 67698 158596
rect 170214 158584 170220 158596
rect 170272 158584 170278 158636
rect 171962 158584 171968 158636
rect 172020 158624 172026 158636
rect 249794 158624 249800 158636
rect 172020 158596 249800 158624
rect 172020 158584 172026 158596
rect 249794 158584 249800 158596
rect 249852 158584 249858 158636
rect 74350 158516 74356 158568
rect 74408 158556 74414 158568
rect 175366 158556 175372 158568
rect 74408 158528 175372 158556
rect 74408 158516 74414 158528
rect 175366 158516 175372 158528
rect 175424 158516 175430 158568
rect 178678 158516 178684 158568
rect 178736 158556 178742 158568
rect 255590 158556 255596 158568
rect 178736 158528 255596 158556
rect 178736 158516 178742 158528
rect 255590 158516 255596 158528
rect 255648 158516 255654 158568
rect 71038 158448 71044 158500
rect 71096 158488 71102 158500
rect 172790 158488 172796 158500
rect 71096 158460 172796 158488
rect 71096 158448 71102 158460
rect 172790 158448 172796 158460
rect 172848 158448 172854 158500
rect 175274 158448 175280 158500
rect 175332 158488 175338 158500
rect 252554 158488 252560 158500
rect 175332 158460 252560 158488
rect 175332 158448 175338 158460
rect 252554 158448 252560 158460
rect 252612 158448 252618 158500
rect 60918 158380 60924 158432
rect 60976 158420 60982 158432
rect 165062 158420 165068 158432
rect 60976 158392 165068 158420
rect 60976 158380 60982 158392
rect 165062 158380 165068 158392
rect 165120 158380 165126 158432
rect 165246 158380 165252 158432
rect 165304 158420 165310 158432
rect 244642 158420 244648 158432
rect 165304 158392 244648 158420
rect 165304 158380 165310 158392
rect 244642 158380 244648 158392
rect 244700 158380 244706 158432
rect 64230 158312 64236 158364
rect 64288 158352 64294 158364
rect 167546 158352 167552 158364
rect 64288 158324 167552 158352
rect 64288 158312 64294 158324
rect 167546 158312 167552 158324
rect 167604 158312 167610 158364
rect 168558 158312 168564 158364
rect 168616 158352 168622 158364
rect 247126 158352 247132 158364
rect 168616 158324 247132 158352
rect 168616 158312 168622 158324
rect 247126 158312 247132 158324
rect 247184 158312 247190 158364
rect 54202 158244 54208 158296
rect 54260 158284 54266 158296
rect 160278 158284 160284 158296
rect 54260 158256 160284 158284
rect 54260 158244 54266 158256
rect 160278 158244 160284 158256
rect 160336 158244 160342 158296
rect 161842 158244 161848 158296
rect 161900 158284 161906 158296
rect 242066 158284 242072 158296
rect 161900 158256 242072 158284
rect 161900 158244 161906 158256
rect 242066 158244 242072 158256
rect 242124 158244 242130 158296
rect 50798 158176 50804 158228
rect 50856 158216 50862 158228
rect 157334 158216 157340 158228
rect 50856 158188 157340 158216
rect 50856 158176 50862 158188
rect 157334 158176 157340 158188
rect 157392 158176 157398 158228
rect 158438 158176 158444 158228
rect 158496 158216 158502 158228
rect 239674 158216 239680 158228
rect 158496 158188 239680 158216
rect 158496 158176 158502 158188
rect 239674 158176 239680 158188
rect 239732 158176 239738 158228
rect 256878 158176 256884 158228
rect 256936 158216 256942 158228
rect 314746 158216 314752 158228
rect 256936 158188 314752 158216
rect 256936 158176 256942 158188
rect 314746 158176 314752 158188
rect 314804 158176 314810 158228
rect 47486 158108 47492 158160
rect 47544 158148 47550 158160
rect 154758 158148 154764 158160
rect 47544 158120 154764 158148
rect 47544 158108 47550 158120
rect 154758 158108 154764 158120
rect 154816 158108 154822 158160
rect 155126 158108 155132 158160
rect 155184 158148 155190 158160
rect 237374 158148 237380 158160
rect 155184 158120 237380 158148
rect 155184 158108 155190 158120
rect 237374 158108 237380 158120
rect 237432 158108 237438 158160
rect 246758 158108 246764 158160
rect 246816 158148 246822 158160
rect 306926 158148 306932 158160
rect 246816 158120 306932 158148
rect 246816 158108 246822 158120
rect 306926 158108 306932 158120
rect 306984 158108 306990 158160
rect 37366 158040 37372 158092
rect 37424 158080 37430 158092
rect 146754 158080 146760 158092
rect 37424 158052 146760 158080
rect 37424 158040 37430 158052
rect 146754 158040 146760 158052
rect 146812 158040 146818 158092
rect 148410 158040 148416 158092
rect 148468 158080 148474 158092
rect 231946 158080 231952 158092
rect 148468 158052 231952 158080
rect 148468 158040 148474 158052
rect 231946 158040 231952 158052
rect 232004 158040 232010 158092
rect 243446 158040 243452 158092
rect 243504 158080 243510 158092
rect 304350 158080 304356 158092
rect 243504 158052 304356 158080
rect 243504 158040 243510 158052
rect 304350 158040 304356 158052
rect 304408 158040 304414 158092
rect 382 157972 388 158024
rect 440 158012 446 158024
rect 118878 158012 118884 158024
rect 440 157984 118884 158012
rect 440 157972 446 157984
rect 118878 157972 118884 157984
rect 118936 157972 118942 158024
rect 131574 157972 131580 158024
rect 131632 158012 131638 158024
rect 218974 158012 218980 158024
rect 131632 157984 218980 158012
rect 131632 157972 131638 157984
rect 218974 157972 218980 157984
rect 219032 157972 219038 158024
rect 236730 157972 236736 158024
rect 236788 158012 236794 158024
rect 299566 158012 299572 158024
rect 236788 157984 299572 158012
rect 236788 157972 236794 157984
rect 299566 157972 299572 157984
rect 299624 157972 299630 158024
rect 77754 157904 77760 157956
rect 77812 157944 77818 157956
rect 77812 157916 176056 157944
rect 77812 157904 77818 157916
rect 84470 157836 84476 157888
rect 84528 157876 84534 157888
rect 175918 157876 175924 157888
rect 84528 157848 175924 157876
rect 84528 157836 84534 157848
rect 175918 157836 175924 157848
rect 175976 157836 175982 157888
rect 176028 157876 176056 157916
rect 176194 157904 176200 157956
rect 176252 157944 176258 157956
rect 183002 157944 183008 157956
rect 176252 157916 183008 157944
rect 176252 157904 176258 157916
rect 183002 157904 183008 157916
rect 183060 157904 183066 157956
rect 185394 157904 185400 157956
rect 185452 157944 185458 157956
rect 260098 157944 260104 157956
rect 185452 157916 260104 157944
rect 185452 157904 185458 157916
rect 260098 157904 260104 157916
rect 260156 157904 260162 157956
rect 178034 157876 178040 157888
rect 176028 157848 178040 157876
rect 178034 157836 178040 157848
rect 178092 157836 178098 157888
rect 180702 157836 180708 157888
rect 180760 157876 180766 157888
rect 181346 157876 181352 157888
rect 180760 157848 181352 157876
rect 180760 157836 180766 157848
rect 181346 157836 181352 157848
rect 181404 157836 181410 157888
rect 181530 157836 181536 157888
rect 181588 157876 181594 157888
rect 188154 157876 188160 157888
rect 181588 157848 188160 157876
rect 181588 157836 181594 157848
rect 188154 157836 188160 157848
rect 188212 157836 188218 157888
rect 188798 157836 188804 157888
rect 188856 157876 188862 157888
rect 262674 157876 262680 157888
rect 188856 157848 262680 157876
rect 188856 157836 188862 157848
rect 262674 157836 262680 157848
rect 262732 157836 262738 157888
rect 87782 157768 87788 157820
rect 87840 157808 87846 157820
rect 87840 157780 181300 157808
rect 87840 157768 87846 157780
rect 91186 157700 91192 157752
rect 91244 157740 91250 157752
rect 181070 157740 181076 157752
rect 91244 157712 181076 157740
rect 91244 157700 91250 157712
rect 181070 157700 181076 157712
rect 181128 157700 181134 157752
rect 94590 157632 94596 157684
rect 94648 157672 94654 157684
rect 181162 157672 181168 157684
rect 94648 157644 181168 157672
rect 94648 157632 94654 157644
rect 181162 157632 181168 157644
rect 181220 157632 181226 157684
rect 181272 157672 181300 157780
rect 181806 157768 181812 157820
rect 181864 157808 181870 157820
rect 190638 157808 190644 157820
rect 181864 157780 190644 157808
rect 181864 157768 181870 157780
rect 190638 157768 190644 157780
rect 190696 157768 190702 157820
rect 195514 157768 195520 157820
rect 195572 157808 195578 157820
rect 267734 157808 267740 157820
rect 195572 157780 267740 157808
rect 195572 157768 195578 157780
rect 267734 157768 267740 157780
rect 267792 157768 267798 157820
rect 181714 157700 181720 157752
rect 181772 157740 181778 157752
rect 181772 157712 186314 157740
rect 181772 157700 181778 157712
rect 185578 157672 185584 157684
rect 181272 157644 185584 157672
rect 185578 157632 185584 157644
rect 185636 157632 185642 157684
rect 186286 157672 186314 157712
rect 190454 157700 190460 157752
rect 190512 157740 190518 157752
rect 264054 157740 264060 157752
rect 190512 157712 264060 157740
rect 190512 157700 190518 157712
rect 264054 157700 264060 157712
rect 264112 157700 264118 157752
rect 236086 157672 236092 157684
rect 186286 157644 236092 157672
rect 236086 157632 236092 157644
rect 236144 157632 236150 157684
rect 97902 157564 97908 157616
rect 97960 157604 97966 157616
rect 193214 157604 193220 157616
rect 97960 157576 193220 157604
rect 97960 157564 97966 157576
rect 193214 157564 193220 157576
rect 193272 157564 193278 157616
rect 197354 157564 197360 157616
rect 197412 157604 197418 157616
rect 251266 157604 251272 157616
rect 197412 157576 251272 157604
rect 197412 157564 197418 157576
rect 251266 157564 251272 157576
rect 251324 157564 251330 157616
rect 111334 157496 111340 157548
rect 111392 157536 111398 157548
rect 203426 157536 203432 157548
rect 111392 157508 203432 157536
rect 111392 157496 111398 157508
rect 203426 157496 203432 157508
rect 203484 157496 203490 157548
rect 204898 157496 204904 157548
rect 204956 157536 204962 157548
rect 255866 157536 255872 157548
rect 204956 157508 255872 157536
rect 204956 157496 204962 157508
rect 255866 157496 255872 157508
rect 255924 157496 255930 157548
rect 114738 157428 114744 157480
rect 114796 157468 114802 157480
rect 206186 157468 206192 157480
rect 114796 157440 206192 157468
rect 114796 157428 114802 157440
rect 206186 157428 206192 157440
rect 206244 157428 206250 157480
rect 141694 157360 141700 157412
rect 141752 157400 141758 157412
rect 226702 157400 226708 157412
rect 141752 157372 226708 157400
rect 141752 157360 141758 157372
rect 226702 157360 226708 157372
rect 226760 157360 226766 157412
rect 49142 157292 49148 157344
rect 49200 157332 49206 157344
rect 156046 157332 156052 157344
rect 49200 157304 156052 157332
rect 49200 157292 49206 157304
rect 156046 157292 156052 157304
rect 156104 157292 156110 157344
rect 158714 157292 158720 157344
rect 158772 157332 158778 157344
rect 214466 157332 214472 157344
rect 158772 157304 214472 157332
rect 158772 157292 158778 157304
rect 214466 157292 214472 157304
rect 214524 157292 214530 157344
rect 214558 157292 214564 157344
rect 214616 157332 214622 157344
rect 221366 157332 221372 157344
rect 214616 157304 221372 157332
rect 214616 157292 214622 157304
rect 221366 157292 221372 157304
rect 221424 157292 221430 157344
rect 224218 157292 224224 157344
rect 224276 157332 224282 157344
rect 281626 157332 281632 157344
rect 224276 157304 281632 157332
rect 224276 157292 224282 157304
rect 281626 157292 281632 157304
rect 281684 157292 281690 157344
rect 45738 157224 45744 157276
rect 45796 157264 45802 157276
rect 153562 157264 153568 157276
rect 45796 157236 153568 157264
rect 45796 157224 45802 157236
rect 153562 157224 153568 157236
rect 153620 157224 153626 157276
rect 164142 157224 164148 157276
rect 164200 157264 164206 157276
rect 166258 157264 166264 157276
rect 164200 157236 166264 157264
rect 164200 157224 164206 157236
rect 166258 157224 166264 157236
rect 166316 157224 166322 157276
rect 192110 157224 192116 157276
rect 192168 157264 192174 157276
rect 265158 157264 265164 157276
rect 192168 157236 265164 157264
rect 192168 157224 192174 157236
rect 265158 157224 265164 157236
rect 265216 157224 265222 157276
rect 283834 157224 283840 157276
rect 283892 157264 283898 157276
rect 335446 157264 335452 157276
rect 283892 157236 335452 157264
rect 283892 157224 283898 157236
rect 335446 157224 335452 157236
rect 335504 157224 335510 157276
rect 39022 157156 39028 157208
rect 39080 157196 39086 157208
rect 148226 157196 148232 157208
rect 39080 157168 148232 157196
rect 39080 157156 39086 157168
rect 148226 157156 148232 157168
rect 148284 157156 148290 157208
rect 150066 157156 150072 157208
rect 150124 157196 150130 157208
rect 233510 157196 233516 157208
rect 150124 157168 233516 157196
rect 150124 157156 150130 157168
rect 233510 157156 233516 157168
rect 233568 157156 233574 157208
rect 290550 157156 290556 157208
rect 290608 157196 290614 157208
rect 340046 157196 340052 157208
rect 290608 157168 340052 157196
rect 290608 157156 290614 157168
rect 340046 157156 340052 157168
rect 340104 157156 340110 157208
rect 42426 157088 42432 157140
rect 42484 157128 42490 157140
rect 150894 157128 150900 157140
rect 42484 157100 150900 157128
rect 42484 157088 42490 157100
rect 150894 157088 150900 157100
rect 150952 157088 150958 157140
rect 156506 157088 156512 157140
rect 156564 157128 156570 157140
rect 158898 157128 158904 157140
rect 156564 157100 158904 157128
rect 156564 157088 156570 157100
rect 158898 157088 158904 157100
rect 158956 157088 158962 157140
rect 160094 157088 160100 157140
rect 160152 157128 160158 157140
rect 165890 157128 165896 157140
rect 160152 157100 165896 157128
rect 160152 157088 160158 157100
rect 165890 157088 165896 157100
rect 165948 157088 165954 157140
rect 165982 157088 165988 157140
rect 166040 157128 166046 157140
rect 171594 157128 171600 157140
rect 166040 157100 171600 157128
rect 166040 157088 166046 157100
rect 171594 157088 171600 157100
rect 171652 157088 171658 157140
rect 177022 157088 177028 157140
rect 177080 157128 177086 157140
rect 254026 157128 254032 157140
rect 177080 157100 254032 157128
rect 177080 157088 177086 157100
rect 254026 157088 254032 157100
rect 254084 157088 254090 157140
rect 287146 157088 287152 157140
rect 287204 157128 287210 157140
rect 338114 157128 338120 157140
rect 287204 157100 338120 157128
rect 287204 157088 287210 157100
rect 338114 157088 338120 157100
rect 338172 157088 338178 157140
rect 35710 157020 35716 157072
rect 35768 157060 35774 157072
rect 145926 157060 145932 157072
rect 35768 157032 145932 157060
rect 35768 157020 35774 157032
rect 145926 157020 145932 157032
rect 145984 157020 145990 157072
rect 151722 157020 151728 157072
rect 151780 157060 151786 157072
rect 234798 157060 234804 157072
rect 151780 157032 234804 157060
rect 151780 157020 151786 157032
rect 234798 157020 234804 157032
rect 234856 157020 234862 157072
rect 280430 157020 280436 157072
rect 280488 157060 280494 157072
rect 332870 157060 332876 157072
rect 280488 157032 332876 157060
rect 280488 157020 280494 157032
rect 332870 157020 332876 157032
rect 332928 157020 332934 157072
rect 24762 156952 24768 157004
rect 24820 156992 24826 157004
rect 137370 156992 137376 157004
rect 24820 156964 137376 156992
rect 24820 156952 24826 156964
rect 137370 156952 137376 156964
rect 137428 156952 137434 157004
rect 138290 156952 138296 157004
rect 138348 156992 138354 157004
rect 224126 156992 224132 157004
rect 138348 156964 224132 156992
rect 138348 156952 138354 156964
rect 224126 156952 224132 156964
rect 224184 156952 224190 157004
rect 273714 156952 273720 157004
rect 273772 156992 273778 157004
rect 327534 156992 327540 157004
rect 273772 156964 327540 156992
rect 273772 156952 273778 156964
rect 327534 156952 327540 156964
rect 327592 156952 327598 157004
rect 18046 156884 18052 156936
rect 18104 156924 18110 156936
rect 132494 156924 132500 156936
rect 18104 156896 132500 156924
rect 18104 156884 18110 156896
rect 132494 156884 132500 156896
rect 132552 156884 132558 156936
rect 134886 156884 134892 156936
rect 134944 156924 134950 156936
rect 214558 156924 214564 156936
rect 134944 156896 214564 156924
rect 134944 156884 134950 156896
rect 214558 156884 214564 156896
rect 214616 156884 214622 156936
rect 224954 156884 224960 156936
rect 225012 156924 225018 156936
rect 272058 156924 272064 156936
rect 225012 156896 272064 156924
rect 225012 156884 225018 156896
rect 272058 156884 272064 156896
rect 272116 156884 272122 156936
rect 277118 156884 277124 156936
rect 277176 156924 277182 156936
rect 330018 156924 330024 156936
rect 277176 156896 330024 156924
rect 277176 156884 277182 156896
rect 330018 156884 330024 156896
rect 330076 156884 330082 156936
rect 21358 156816 21364 156868
rect 21416 156856 21422 156868
rect 135254 156856 135260 156868
rect 21416 156828 135260 156856
rect 21416 156816 21422 156828
rect 135254 156816 135260 156828
rect 135312 156816 135318 156868
rect 135806 156816 135812 156868
rect 135864 156856 135870 156868
rect 222378 156856 222384 156868
rect 135864 156828 222384 156856
rect 135864 156816 135870 156828
rect 222378 156816 222384 156828
rect 222436 156816 222442 156868
rect 226610 156816 226616 156868
rect 226668 156856 226674 156868
rect 291562 156856 291568 156868
rect 226668 156828 291568 156856
rect 226668 156816 226674 156828
rect 291562 156816 291568 156828
rect 291620 156816 291626 156868
rect 300670 156816 300676 156868
rect 300728 156856 300734 156868
rect 348050 156856 348056 156868
rect 300728 156828 348056 156856
rect 300728 156816 300734 156828
rect 348050 156816 348056 156828
rect 348108 156816 348114 156868
rect 14642 156748 14648 156800
rect 14700 156788 14706 156800
rect 129826 156788 129832 156800
rect 14700 156760 129832 156788
rect 14700 156748 14706 156760
rect 129826 156748 129832 156760
rect 129884 156748 129890 156800
rect 139118 156748 139124 156800
rect 139176 156788 139182 156800
rect 225138 156788 225144 156800
rect 139176 156760 225144 156788
rect 139176 156748 139182 156760
rect 225138 156748 225144 156760
rect 225196 156748 225202 156800
rect 230014 156748 230020 156800
rect 230072 156788 230078 156800
rect 294046 156788 294052 156800
rect 230072 156760 294052 156788
rect 230072 156748 230078 156760
rect 294046 156748 294052 156760
rect 294104 156748 294110 156800
rect 297266 156748 297272 156800
rect 297324 156788 297330 156800
rect 345566 156788 345572 156800
rect 297324 156760 345572 156788
rect 297324 156748 297330 156760
rect 345566 156748 345572 156760
rect 345624 156748 345630 156800
rect 11238 156680 11244 156732
rect 11296 156720 11302 156732
rect 127158 156720 127164 156732
rect 11296 156692 127164 156720
rect 11296 156680 11302 156692
rect 127158 156680 127164 156692
rect 127216 156680 127222 156732
rect 128170 156680 128176 156732
rect 128228 156720 128234 156732
rect 216674 156720 216680 156732
rect 128228 156692 216680 156720
rect 128228 156680 128234 156692
rect 216674 156680 216680 156692
rect 216732 156680 216738 156732
rect 223206 156680 223212 156732
rect 223264 156720 223270 156732
rect 288986 156720 288992 156732
rect 223264 156692 288992 156720
rect 223264 156680 223270 156692
rect 288986 156680 288992 156692
rect 289044 156680 289050 156732
rect 293862 156680 293868 156732
rect 293920 156720 293926 156732
rect 342806 156720 342812 156732
rect 293920 156692 342812 156720
rect 293920 156680 293926 156692
rect 342806 156680 342812 156692
rect 342864 156680 342870 156732
rect 2038 156612 2044 156664
rect 2096 156652 2102 156664
rect 120166 156652 120172 156664
rect 2096 156624 120172 156652
rect 2096 156612 2102 156624
rect 120166 156612 120172 156624
rect 120224 156612 120230 156664
rect 124858 156612 124864 156664
rect 124916 156652 124922 156664
rect 213914 156652 213920 156664
rect 124916 156624 213920 156652
rect 124916 156612 124922 156624
rect 213914 156612 213920 156624
rect 213972 156612 213978 156664
rect 216490 156612 216496 156664
rect 216548 156652 216554 156664
rect 283098 156652 283104 156664
rect 216548 156624 283104 156652
rect 216548 156612 216554 156624
rect 283098 156612 283104 156624
rect 283156 156612 283162 156664
rect 52454 156544 52460 156596
rect 52512 156584 52518 156596
rect 158806 156584 158812 156596
rect 52512 156556 158812 156584
rect 52512 156544 52518 156556
rect 158806 156544 158812 156556
rect 158864 156544 158870 156596
rect 158898 156544 158904 156596
rect 158956 156584 158962 156596
rect 200758 156584 200764 156596
rect 158956 156556 200764 156584
rect 158956 156544 158962 156556
rect 200758 156544 200764 156556
rect 200816 156544 200822 156596
rect 200942 156544 200948 156596
rect 201000 156584 201006 156596
rect 270494 156584 270500 156596
rect 201000 156556 270500 156584
rect 201000 156544 201006 156556
rect 270494 156544 270500 156556
rect 270552 156544 270558 156596
rect 59262 156476 59268 156528
rect 59320 156516 59326 156528
rect 163774 156516 163780 156528
rect 59320 156488 163780 156516
rect 59320 156476 59326 156488
rect 163774 156476 163780 156488
rect 163832 156476 163838 156528
rect 165890 156476 165896 156528
rect 165948 156516 165954 156528
rect 165948 156488 166120 156516
rect 165948 156476 165954 156488
rect 69290 156408 69296 156460
rect 69348 156448 69354 156460
rect 165982 156448 165988 156460
rect 69348 156420 165988 156448
rect 69348 156408 69354 156420
rect 165982 156408 165988 156420
rect 166040 156408 166046 156460
rect 166092 156448 166120 156488
rect 166258 156476 166264 156528
rect 166316 156516 166322 156528
rect 225506 156516 225512 156528
rect 166316 156488 225512 156516
rect 166316 156476 166322 156488
rect 225506 156476 225512 156488
rect 225564 156476 225570 156528
rect 228082 156448 228088 156460
rect 166092 156420 228088 156448
rect 228082 156408 228088 156420
rect 228140 156408 228146 156460
rect 82814 156340 82820 156392
rect 82872 156380 82878 156392
rect 181806 156380 181812 156392
rect 82872 156352 181812 156380
rect 82872 156340 82878 156352
rect 181806 156340 181812 156352
rect 181864 156340 181870 156392
rect 198826 156340 198832 156392
rect 198884 156380 198890 156392
rect 200942 156380 200948 156392
rect 198884 156352 200948 156380
rect 198884 156340 198890 156352
rect 200942 156340 200948 156352
rect 201000 156340 201006 156392
rect 209774 156340 209780 156392
rect 209832 156380 209838 156392
rect 278958 156380 278964 156392
rect 209832 156352 278964 156380
rect 209832 156340 209838 156352
rect 278958 156340 278964 156352
rect 279016 156340 279022 156392
rect 101306 156272 101312 156324
rect 101364 156312 101370 156324
rect 196158 156312 196164 156324
rect 101364 156284 196164 156312
rect 101364 156272 101370 156284
rect 196158 156272 196164 156284
rect 196216 156272 196222 156324
rect 200758 156272 200764 156324
rect 200816 156312 200822 156324
rect 200816 156284 212672 156312
rect 200816 156272 200822 156284
rect 99558 156204 99564 156256
rect 99616 156244 99622 156256
rect 194686 156244 194692 156256
rect 99616 156216 194692 156244
rect 99616 156204 99622 156216
rect 194686 156204 194692 156216
rect 194744 156204 194750 156256
rect 197998 156204 198004 156256
rect 198056 156244 198062 156256
rect 211338 156244 211344 156256
rect 198056 156216 211344 156244
rect 198056 156204 198062 156216
rect 211338 156204 211344 156216
rect 211396 156204 211402 156256
rect 108022 156136 108028 156188
rect 108080 156176 108086 156188
rect 200666 156176 200672 156188
rect 108080 156148 200672 156176
rect 108080 156136 108086 156148
rect 200666 156136 200672 156148
rect 200724 156136 200730 156188
rect 208762 156176 208768 156188
rect 201236 156148 208768 156176
rect 118142 156068 118148 156120
rect 118200 156108 118206 156120
rect 201236 156108 201264 156148
rect 208762 156136 208768 156148
rect 208820 156136 208826 156188
rect 212644 156176 212672 156284
rect 213178 156272 213184 156324
rect 213236 156312 213242 156324
rect 224218 156312 224224 156324
rect 213236 156284 224224 156312
rect 213236 156272 213242 156284
rect 224218 156272 224224 156284
rect 224276 156272 224282 156324
rect 286226 156312 286232 156324
rect 224328 156284 286232 156312
rect 214466 156204 214472 156256
rect 214524 156244 214530 156256
rect 219986 156244 219992 156256
rect 214524 156216 219992 156244
rect 214524 156204 214530 156216
rect 219986 156204 219992 156216
rect 220044 156204 220050 156256
rect 220078 156204 220084 156256
rect 220136 156244 220142 156256
rect 224328 156244 224356 156284
rect 286226 156272 286232 156284
rect 286284 156272 286290 156324
rect 266538 156244 266544 156256
rect 220136 156216 224356 156244
rect 229066 156216 266544 156244
rect 220136 156204 220142 156216
rect 215478 156176 215484 156188
rect 212644 156148 215484 156176
rect 215478 156136 215484 156148
rect 215536 156136 215542 156188
rect 218054 156136 218060 156188
rect 218112 156176 218118 156188
rect 229066 156176 229094 156216
rect 266538 156204 266544 156216
rect 266596 156204 266602 156256
rect 218112 156148 229094 156176
rect 218112 156136 218118 156148
rect 230750 156136 230756 156188
rect 230808 156176 230814 156188
rect 276750 156176 276756 156188
rect 230808 156148 276756 156176
rect 230808 156136 230814 156148
rect 276750 156136 276756 156148
rect 276808 156136 276814 156188
rect 118200 156080 201264 156108
rect 118200 156068 118206 156080
rect 203058 156068 203064 156120
rect 203116 156108 203122 156120
rect 273530 156108 273536 156120
rect 203116 156080 273536 156108
rect 203116 156068 203122 156080
rect 273530 156068 273536 156080
rect 273588 156068 273594 156120
rect 121454 156000 121460 156052
rect 121512 156040 121518 156052
rect 197998 156040 198004 156052
rect 121512 156012 198004 156040
rect 121512 156000 121518 156012
rect 197998 156000 198004 156012
rect 198056 156000 198062 156052
rect 202230 156000 202236 156052
rect 202288 156040 202294 156052
rect 273346 156040 273352 156052
rect 202288 156012 273352 156040
rect 202288 156000 202294 156012
rect 273346 156000 273352 156012
rect 273404 156000 273410 156052
rect 145006 155932 145012 155984
rect 145064 155972 145070 155984
rect 229278 155972 229284 155984
rect 145064 155944 229284 155972
rect 145064 155932 145070 155944
rect 229278 155932 229284 155944
rect 229336 155932 229342 155984
rect 66806 155864 66812 155916
rect 66864 155904 66870 155916
rect 82906 155904 82912 155916
rect 66864 155876 82912 155904
rect 66864 155864 66870 155876
rect 82906 155864 82912 155876
rect 82964 155864 82970 155916
rect 92014 155864 92020 155916
rect 92072 155904 92078 155916
rect 92072 155876 186544 155904
rect 92072 155864 92078 155876
rect 60090 155796 60096 155848
rect 60148 155836 60154 155848
rect 78766 155836 78772 155848
rect 60148 155808 78772 155836
rect 60148 155796 60154 155808
rect 78766 155796 78772 155808
rect 78824 155796 78830 155848
rect 88702 155796 88708 155848
rect 88760 155836 88766 155848
rect 186406 155836 186412 155848
rect 88760 155808 186412 155836
rect 88760 155796 88766 155808
rect 186406 155796 186412 155808
rect 186464 155796 186470 155848
rect 186516 155836 186544 155876
rect 186590 155864 186596 155916
rect 186648 155904 186654 155916
rect 194042 155904 194048 155916
rect 186648 155876 194048 155904
rect 186648 155864 186654 155876
rect 194042 155864 194048 155876
rect 194100 155864 194106 155916
rect 196342 155864 196348 155916
rect 196400 155904 196406 155916
rect 268470 155904 268476 155916
rect 196400 155876 268476 155904
rect 196400 155864 196406 155876
rect 268470 155864 268476 155876
rect 268528 155864 268534 155916
rect 296438 155864 296444 155916
rect 296496 155904 296502 155916
rect 345198 155904 345204 155916
rect 296496 155876 345204 155904
rect 296496 155864 296502 155876
rect 345198 155864 345204 155876
rect 345256 155864 345262 155916
rect 189074 155836 189080 155848
rect 186516 155808 189080 155836
rect 189074 155796 189080 155808
rect 189132 155796 189138 155848
rect 192938 155796 192944 155848
rect 192996 155836 193002 155848
rect 265894 155836 265900 155848
rect 192996 155808 265900 155836
rect 192996 155796 193002 155808
rect 265894 155796 265900 155808
rect 265952 155796 265958 155848
rect 293034 155796 293040 155848
rect 293092 155836 293098 155848
rect 342346 155836 342352 155848
rect 293092 155808 342352 155836
rect 293092 155796 293098 155808
rect 342346 155796 342352 155808
rect 342404 155796 342410 155848
rect 12158 155728 12164 155780
rect 12216 155768 12222 155780
rect 110322 155768 110328 155780
rect 12216 155740 110328 155768
rect 12216 155728 12222 155740
rect 110322 155728 110328 155740
rect 110380 155728 110386 155780
rect 112254 155728 112260 155780
rect 112312 155768 112318 155780
rect 204346 155768 204352 155780
rect 112312 155740 204352 155768
rect 112312 155728 112318 155740
rect 204346 155728 204352 155740
rect 204404 155728 204410 155780
rect 206462 155728 206468 155780
rect 206520 155768 206526 155780
rect 276106 155768 276112 155780
rect 206520 155740 276112 155768
rect 206520 155728 206526 155740
rect 276106 155728 276112 155740
rect 276164 155728 276170 155780
rect 289722 155728 289728 155780
rect 289780 155768 289786 155780
rect 339586 155768 339592 155780
rect 289780 155740 339592 155768
rect 289780 155728 289786 155740
rect 339586 155728 339592 155740
rect 339644 155728 339650 155780
rect 46566 155660 46572 155712
rect 46624 155700 46630 155712
rect 75086 155700 75092 155712
rect 46624 155672 75092 155700
rect 46624 155660 46630 155672
rect 75086 155660 75092 155672
rect 75144 155660 75150 155712
rect 81894 155660 81900 155712
rect 81952 155700 81958 155712
rect 181162 155700 181168 155712
rect 81952 155672 181168 155700
rect 81952 155660 81958 155672
rect 181162 155660 181168 155672
rect 181220 155660 181226 155712
rect 186222 155660 186228 155712
rect 186280 155700 186286 155712
rect 260926 155700 260932 155712
rect 186280 155672 260932 155700
rect 186280 155660 186286 155672
rect 260926 155660 260932 155672
rect 260984 155660 260990 155712
rect 270310 155660 270316 155712
rect 270368 155700 270374 155712
rect 324958 155700 324964 155712
rect 270368 155672 324964 155700
rect 270368 155660 270374 155672
rect 324958 155660 324964 155672
rect 325016 155660 325022 155712
rect 340966 155660 340972 155712
rect 341024 155700 341030 155712
rect 378686 155700 378692 155712
rect 341024 155672 378692 155700
rect 341024 155660 341030 155672
rect 378686 155660 378692 155672
rect 378744 155660 378750 155712
rect 53374 155592 53380 155644
rect 53432 155632 53438 155644
rect 66622 155632 66628 155644
rect 53432 155604 66628 155632
rect 53432 155592 53438 155604
rect 66622 155592 66628 155604
rect 66680 155592 66686 155644
rect 71866 155592 71872 155644
rect 71924 155632 71930 155644
rect 173526 155632 173532 155644
rect 71924 155604 173532 155632
rect 71924 155592 71930 155604
rect 173526 155592 173532 155604
rect 173584 155592 173590 155644
rect 176286 155592 176292 155644
rect 176344 155632 176350 155644
rect 253014 155632 253020 155644
rect 176344 155604 253020 155632
rect 176344 155592 176350 155604
rect 253014 155592 253020 155604
rect 253072 155592 253078 155644
rect 266998 155592 267004 155644
rect 267056 155632 267062 155644
rect 322106 155632 322112 155644
rect 267056 155604 322112 155632
rect 267056 155592 267062 155604
rect 322106 155592 322112 155604
rect 322164 155592 322170 155644
rect 344370 155592 344376 155644
rect 344428 155632 344434 155644
rect 381446 155632 381452 155644
rect 344428 155604 381452 155632
rect 344428 155592 344434 155604
rect 381446 155592 381452 155604
rect 381504 155592 381510 155644
rect 39850 155524 39856 155576
rect 39908 155564 39914 155576
rect 68922 155564 68928 155576
rect 39908 155536 68928 155564
rect 39908 155524 39914 155536
rect 68922 155524 68928 155536
rect 68980 155524 68986 155576
rect 75178 155524 75184 155576
rect 75236 155564 75242 155576
rect 176010 155564 176016 155576
rect 75236 155536 176016 155564
rect 75236 155524 75242 155536
rect 176010 155524 176016 155536
rect 176068 155524 176074 155576
rect 179506 155524 179512 155576
rect 179564 155564 179570 155576
rect 255682 155564 255688 155576
rect 179564 155536 255688 155564
rect 179564 155524 179570 155536
rect 255682 155524 255688 155536
rect 255740 155524 255746 155576
rect 263594 155524 263600 155576
rect 263652 155564 263658 155576
rect 320174 155564 320180 155576
rect 263652 155536 320180 155564
rect 263652 155524 263658 155536
rect 320174 155524 320180 155536
rect 320232 155524 320238 155576
rect 337654 155524 337660 155576
rect 337712 155564 337718 155576
rect 376294 155564 376300 155576
rect 337712 155536 376300 155564
rect 337712 155524 337718 155536
rect 376294 155524 376300 155536
rect 376352 155524 376358 155576
rect 65150 155456 65156 155508
rect 65208 155496 65214 155508
rect 168558 155496 168564 155508
rect 65208 155468 168564 155496
rect 65208 155456 65214 155468
rect 168558 155456 168564 155468
rect 168616 155456 168622 155508
rect 169386 155456 169392 155508
rect 169444 155496 169450 155508
rect 247862 155496 247868 155508
rect 169444 155468 247868 155496
rect 169444 155456 169450 155468
rect 247862 155456 247868 155468
rect 247920 155456 247926 155508
rect 260282 155456 260288 155508
rect 260340 155496 260346 155508
rect 317598 155496 317604 155508
rect 260340 155468 317604 155496
rect 260340 155456 260346 155468
rect 317598 155456 317604 155468
rect 317656 155456 317662 155508
rect 333422 155456 333428 155508
rect 333480 155496 333486 155508
rect 373074 155496 373080 155508
rect 333480 155468 373080 155496
rect 333480 155456 333486 155468
rect 373074 155456 373080 155468
rect 373132 155456 373138 155508
rect 7926 155388 7932 155440
rect 7984 155428 7990 155440
rect 124582 155428 124588 155440
rect 7984 155400 124588 155428
rect 7984 155388 7990 155400
rect 124582 155388 124588 155400
rect 124640 155388 124646 155440
rect 145834 155388 145840 155440
rect 145892 155428 145898 155440
rect 230014 155428 230020 155440
rect 145892 155400 230020 155428
rect 145892 155388 145898 155400
rect 230014 155388 230020 155400
rect 230072 155388 230078 155440
rect 253566 155388 253572 155440
rect 253624 155428 253630 155440
rect 312078 155428 312084 155440
rect 253624 155400 312084 155428
rect 253624 155388 253630 155400
rect 312078 155388 312084 155400
rect 312136 155388 312142 155440
rect 330110 155388 330116 155440
rect 330168 155428 330174 155440
rect 370498 155428 370504 155440
rect 330168 155400 370504 155428
rect 330168 155388 330174 155400
rect 370498 155388 370504 155400
rect 370556 155388 370562 155440
rect 8754 155320 8760 155372
rect 8812 155360 8818 155372
rect 125778 155360 125784 155372
rect 8812 155332 125784 155360
rect 8812 155320 8818 155332
rect 125778 155320 125784 155332
rect 125836 155320 125842 155372
rect 142522 155320 142528 155372
rect 142580 155360 142586 155372
rect 227898 155360 227904 155372
rect 142580 155332 227904 155360
rect 142580 155320 142586 155332
rect 227898 155320 227904 155332
rect 227956 155320 227962 155372
rect 250162 155320 250168 155372
rect 250220 155360 250226 155372
rect 309502 155360 309508 155372
rect 250220 155332 309508 155360
rect 250220 155320 250226 155332
rect 309502 155320 309508 155332
rect 309560 155320 309566 155372
rect 319990 155320 319996 155372
rect 320048 155360 320054 155372
rect 363138 155360 363144 155372
rect 320048 155332 363144 155360
rect 320048 155320 320054 155332
rect 363138 155320 363144 155332
rect 363196 155320 363202 155372
rect 4522 155252 4528 155304
rect 4580 155292 4586 155304
rect 122006 155292 122012 155304
rect 4580 155264 122012 155292
rect 4580 155252 4586 155264
rect 122006 155252 122012 155264
rect 122064 155252 122070 155304
rect 128998 155252 129004 155304
rect 129056 155292 129062 155304
rect 217042 155292 217048 155304
rect 129056 155264 217048 155292
rect 129056 155252 129062 155264
rect 217042 155252 217048 155264
rect 217100 155252 217106 155304
rect 233326 155252 233332 155304
rect 233384 155292 233390 155304
rect 296806 155292 296812 155304
rect 233384 155264 296812 155292
rect 233384 155252 233390 155264
rect 296806 155252 296812 155264
rect 296864 155252 296870 155304
rect 299750 155252 299756 155304
rect 299808 155292 299814 155304
rect 347958 155292 347964 155304
rect 299808 155264 347964 155292
rect 299808 155252 299814 155264
rect 347958 155252 347964 155264
rect 348016 155252 348022 155304
rect 373810 155252 373816 155304
rect 373868 155292 373874 155304
rect 403526 155292 403532 155304
rect 373868 155264 403532 155292
rect 373868 155252 373874 155264
rect 403526 155252 403532 155264
rect 403584 155252 403590 155304
rect 5350 155184 5356 155236
rect 5408 155224 5414 155236
rect 122926 155224 122932 155236
rect 5408 155196 122932 155224
rect 5408 155184 5414 155196
rect 122926 155184 122932 155196
rect 122984 155184 122990 155236
rect 125686 155184 125692 155236
rect 125744 155224 125750 155236
rect 214466 155224 214472 155236
rect 125744 155196 214472 155224
rect 125744 155184 125750 155196
rect 214466 155184 214472 155196
rect 214524 155184 214530 155236
rect 240042 155184 240048 155236
rect 240100 155224 240106 155236
rect 302510 155224 302516 155236
rect 240100 155196 302516 155224
rect 240100 155184 240106 155196
rect 302510 155184 302516 155196
rect 302568 155184 302574 155236
rect 306558 155184 306564 155236
rect 306616 155224 306622 155236
rect 352466 155224 352472 155236
rect 306616 155196 352472 155224
rect 306616 155184 306622 155196
rect 352466 155184 352472 155196
rect 352524 155184 352530 155236
rect 370406 155184 370412 155236
rect 370464 155224 370470 155236
rect 401778 155224 401784 155236
rect 370464 155196 401784 155224
rect 370464 155184 370470 155196
rect 401778 155184 401784 155196
rect 401836 155184 401842 155236
rect 89530 155116 89536 155168
rect 89588 155156 89594 155168
rect 186958 155156 186964 155168
rect 89588 155128 186964 155156
rect 89588 155116 89594 155128
rect 186958 155116 186964 155128
rect 187016 155116 187022 155168
rect 189626 155116 189632 155168
rect 189684 155156 189690 155168
rect 263686 155156 263692 155168
rect 189684 155128 263692 155156
rect 189684 155116 189690 155128
rect 263686 155116 263692 155128
rect 263744 155116 263750 155168
rect 95418 155048 95424 155100
rect 95476 155088 95482 155100
rect 95476 155060 186452 155088
rect 95476 155048 95482 155060
rect 98730 154980 98736 155032
rect 98788 155020 98794 155032
rect 186314 155020 186320 155032
rect 98788 154992 186320 155020
rect 98788 154980 98794 154992
rect 186314 154980 186320 154992
rect 186372 154980 186378 155032
rect 186424 155020 186452 155060
rect 186774 155048 186780 155100
rect 186832 155088 186838 155100
rect 186832 155060 195974 155088
rect 186832 155048 186838 155060
rect 191466 155020 191472 155032
rect 186424 154992 191472 155020
rect 191466 154980 191472 154992
rect 191524 154980 191530 155032
rect 195946 155020 195974 155060
rect 199654 155048 199660 155100
rect 199712 155088 199718 155100
rect 271046 155088 271052 155100
rect 199712 155060 271052 155088
rect 199712 155048 199718 155060
rect 271046 155048 271052 155060
rect 271104 155048 271110 155100
rect 303154 155048 303160 155100
rect 303212 155088 303218 155100
rect 349982 155088 349988 155100
rect 303212 155060 349988 155088
rect 303212 155048 303218 155060
rect 349982 155048 349988 155060
rect 350040 155048 350046 155100
rect 200206 155020 200212 155032
rect 195946 154992 200212 155020
rect 200206 154980 200212 154992
rect 200264 154980 200270 155032
rect 207106 154980 207112 155032
rect 207164 155020 207170 155032
rect 269298 155020 269304 155032
rect 207164 154992 269304 155020
rect 207164 154980 207170 154992
rect 269298 154980 269304 154992
rect 269356 154980 269362 155032
rect 15470 154912 15476 154964
rect 15528 154952 15534 154964
rect 109034 154952 109040 154964
rect 15528 154924 109040 154952
rect 15528 154912 15534 154924
rect 109034 154912 109040 154924
rect 109092 154912 109098 154964
rect 122282 154912 122288 154964
rect 122340 154952 122346 154964
rect 211982 154952 211988 154964
rect 122340 154924 211988 154952
rect 122340 154912 122346 154924
rect 211982 154912 211988 154924
rect 212040 154912 212046 154964
rect 214650 154912 214656 154964
rect 214708 154952 214714 154964
rect 261478 154952 261484 154964
rect 214708 154924 261484 154952
rect 214708 154912 214714 154924
rect 261478 154912 261484 154924
rect 261536 154912 261542 154964
rect 106366 154844 106372 154896
rect 106424 154884 106430 154896
rect 186590 154884 186596 154896
rect 106424 154856 186596 154884
rect 106424 154844 106430 154856
rect 186590 154844 186596 154856
rect 186648 154844 186654 154896
rect 186682 154844 186688 154896
rect 186740 154884 186746 154896
rect 245838 154884 245844 154896
rect 186740 154856 245844 154884
rect 186740 154844 186746 154856
rect 245838 154844 245844 154856
rect 245896 154844 245902 154896
rect 110506 154776 110512 154828
rect 110564 154816 110570 154828
rect 139302 154816 139308 154828
rect 110564 154788 139308 154816
rect 110564 154776 110570 154788
rect 139302 154776 139308 154788
rect 139360 154776 139366 154828
rect 149238 154776 149244 154828
rect 149296 154816 149302 154828
rect 232498 154816 232504 154828
rect 149296 154788 232504 154816
rect 149296 154776 149302 154788
rect 232498 154776 232504 154788
rect 232556 154776 232562 154828
rect 109126 154708 109132 154760
rect 109184 154748 109190 154760
rect 132954 154748 132960 154760
rect 109184 154720 132960 154748
rect 109184 154708 109190 154720
rect 132954 154708 132960 154720
rect 133012 154708 133018 154760
rect 155954 154708 155960 154760
rect 156012 154748 156018 154760
rect 237650 154748 237656 154760
rect 156012 154720 237656 154748
rect 156012 154708 156018 154720
rect 237650 154708 237656 154720
rect 237708 154708 237714 154760
rect 156322 154640 156328 154692
rect 156380 154680 156386 154692
rect 156380 154652 156828 154680
rect 156380 154640 156386 154652
rect 118602 154572 118608 154624
rect 118660 154612 118666 154624
rect 119706 154612 119712 154624
rect 118660 154584 119712 154612
rect 118660 154572 118666 154584
rect 119706 154572 119712 154584
rect 119764 154572 119770 154624
rect 154482 154572 154488 154624
rect 154540 154612 154546 154624
rect 156690 154612 156696 154624
rect 154540 154584 155080 154612
rect 154540 154572 154546 154584
rect 51074 154504 51080 154556
rect 51132 154544 51138 154556
rect 154942 154544 154948 154556
rect 51132 154516 154948 154544
rect 51132 154504 51138 154516
rect 154942 154504 154948 154516
rect 155000 154504 155006 154556
rect 155052 154544 155080 154584
rect 156524 154584 156696 154612
rect 156524 154544 156552 154584
rect 156690 154572 156696 154584
rect 156748 154572 156754 154624
rect 155052 154516 156552 154544
rect 156800 154544 156828 154652
rect 162670 154640 162676 154692
rect 162728 154680 162734 154692
rect 242894 154680 242900 154692
rect 162728 154652 242900 154680
rect 162728 154640 162734 154652
rect 242894 154640 242900 154652
rect 242952 154640 242958 154692
rect 159358 154572 159364 154624
rect 159416 154612 159422 154624
rect 240226 154612 240232 154624
rect 159416 154584 240232 154612
rect 159416 154572 159422 154584
rect 240226 154572 240232 154584
rect 240284 154572 240290 154624
rect 283282 154612 283288 154624
rect 280080 154584 280476 154612
rect 212718 154544 212724 154556
rect 156800 154516 212724 154544
rect 212718 154504 212724 154516
rect 212776 154504 212782 154556
rect 218330 154504 218336 154556
rect 218388 154544 218394 154556
rect 280080 154544 280108 154584
rect 218388 154516 280108 154544
rect 218388 154504 218394 154516
rect 44174 154436 44180 154488
rect 44232 154476 44238 154488
rect 142890 154476 142896 154488
rect 44232 154448 142896 154476
rect 44232 154436 44238 154448
rect 142890 154436 142896 154448
rect 142948 154436 142954 154488
rect 142982 154436 142988 154488
rect 143040 154476 143046 154488
rect 191098 154476 191104 154488
rect 143040 154448 191104 154476
rect 143040 154436 143046 154448
rect 191098 154436 191104 154448
rect 191156 154436 191162 154488
rect 202414 154476 202420 154488
rect 191208 154448 202420 154476
rect 114462 154368 114468 154420
rect 114520 154408 114526 154420
rect 118602 154408 118608 154420
rect 114520 154380 118608 154408
rect 114520 154368 114526 154380
rect 118602 154368 118608 154380
rect 118660 154368 118666 154420
rect 118694 154368 118700 154420
rect 118752 154408 118758 154420
rect 119614 154408 119620 154420
rect 118752 154380 119620 154408
rect 118752 154368 118758 154380
rect 119614 154368 119620 154380
rect 119672 154368 119678 154420
rect 119706 154368 119712 154420
rect 119764 154408 119770 154420
rect 189534 154408 189540 154420
rect 119764 154380 189540 154408
rect 119764 154368 119770 154380
rect 189534 154368 189540 154380
rect 189592 154368 189598 154420
rect 191006 154368 191012 154420
rect 191064 154408 191070 154420
rect 191208 154408 191236 154448
rect 202414 154436 202420 154448
rect 202472 154436 202478 154488
rect 215294 154436 215300 154488
rect 215352 154476 215358 154488
rect 280246 154476 280252 154488
rect 215352 154448 280252 154476
rect 215352 154436 215358 154448
rect 280246 154436 280252 154448
rect 280304 154436 280310 154488
rect 280448 154476 280476 154584
rect 282840 154584 283288 154612
rect 280614 154504 280620 154556
rect 280672 154544 280678 154556
rect 282840 154544 282868 154584
rect 283282 154572 283288 154584
rect 283340 154572 283346 154624
rect 285582 154544 285588 154556
rect 280672 154516 282868 154544
rect 283116 154516 285588 154544
rect 280672 154504 280678 154516
rect 283116 154476 283144 154516
rect 285582 154504 285588 154516
rect 285640 154504 285646 154556
rect 285674 154504 285680 154556
rect 285732 154544 285738 154556
rect 337194 154544 337200 154556
rect 285732 154516 337200 154544
rect 285732 154504 285738 154516
rect 337194 154504 337200 154516
rect 337252 154504 337258 154556
rect 353662 154504 353668 154556
rect 353720 154544 353726 154556
rect 388622 154544 388628 154556
rect 353720 154516 388628 154544
rect 353720 154504 353726 154516
rect 388622 154504 388628 154516
rect 388680 154504 388686 154556
rect 280448 154448 283144 154476
rect 283374 154436 283380 154488
rect 283432 154476 283438 154488
rect 334618 154476 334624 154488
rect 283432 154448 334624 154476
rect 283432 154436 283438 154448
rect 334618 154436 334624 154448
rect 334676 154436 334682 154488
rect 349522 154436 349528 154488
rect 349580 154476 349586 154488
rect 386046 154476 386052 154488
rect 349580 154448 386052 154476
rect 349580 154436 349586 154448
rect 386046 154436 386052 154448
rect 386104 154436 386110 154488
rect 390646 154436 390652 154488
rect 390704 154476 390710 154488
rect 416866 154476 416872 154488
rect 390704 154448 416872 154476
rect 390704 154436 390710 154448
rect 416866 154436 416872 154448
rect 416924 154436 416930 154488
rect 191064 154380 191236 154408
rect 191064 154368 191070 154380
rect 191282 154368 191288 154420
rect 191340 154408 191346 154420
rect 201770 154408 201776 154420
rect 191340 154380 201776 154408
rect 191340 154368 191346 154380
rect 201770 154368 201776 154380
rect 201828 154368 201834 154420
rect 204990 154368 204996 154420
rect 205048 154408 205054 154420
rect 275554 154408 275560 154420
rect 205048 154380 275560 154408
rect 205048 154368 205054 154380
rect 275554 154368 275560 154380
rect 275612 154368 275618 154420
rect 276198 154368 276204 154420
rect 276256 154408 276262 154420
rect 329926 154408 329932 154420
rect 276256 154380 329932 154408
rect 276256 154368 276262 154380
rect 329926 154368 329932 154380
rect 329984 154368 329990 154420
rect 346394 154368 346400 154420
rect 346452 154408 346458 154420
rect 383746 154408 383752 154420
rect 346452 154380 383752 154408
rect 346452 154368 346458 154380
rect 383746 154368 383752 154380
rect 383804 154368 383810 154420
rect 393314 154368 393320 154420
rect 393372 154408 393378 154420
rect 419534 154408 419540 154420
rect 393372 154380 419540 154408
rect 393372 154368 393378 154380
rect 419534 154368 419540 154380
rect 419592 154368 419598 154420
rect 34514 154300 34520 154352
rect 34572 154340 34578 154352
rect 137922 154340 137928 154352
rect 34572 154312 137928 154340
rect 34572 154300 34578 154312
rect 137922 154300 137928 154312
rect 137980 154300 137986 154352
rect 138106 154300 138112 154352
rect 138164 154340 138170 154352
rect 139486 154340 139492 154352
rect 138164 154312 139492 154340
rect 138164 154300 138170 154312
rect 139486 154300 139492 154312
rect 139544 154300 139550 154352
rect 139670 154300 139676 154352
rect 139728 154340 139734 154352
rect 139728 154312 142844 154340
rect 139728 154300 139734 154312
rect 37918 154232 37924 154284
rect 37976 154272 37982 154284
rect 142816 154272 142844 154312
rect 143074 154300 143080 154352
rect 143132 154340 143138 154352
rect 205082 154340 205088 154352
rect 143132 154312 205088 154340
rect 143132 154300 143138 154312
rect 205082 154300 205088 154312
rect 205140 154300 205146 154352
rect 208394 154300 208400 154352
rect 208452 154340 208458 154352
rect 278130 154340 278136 154352
rect 208452 154312 278136 154340
rect 208452 154300 208458 154312
rect 278130 154300 278136 154312
rect 278188 154300 278194 154352
rect 278866 154300 278872 154352
rect 278924 154340 278930 154352
rect 332134 154340 332140 154352
rect 278924 154312 332140 154340
rect 278924 154300 278930 154312
rect 332134 154300 332140 154312
rect 332192 154300 332198 154352
rect 339494 154300 339500 154352
rect 339552 154340 339558 154352
rect 378318 154340 378324 154352
rect 339552 154312 378324 154340
rect 339552 154300 339558 154312
rect 378318 154300 378324 154312
rect 378376 154300 378382 154352
rect 397362 154300 397368 154352
rect 397420 154340 397426 154352
rect 422478 154340 422484 154352
rect 397420 154312 422484 154340
rect 397420 154300 397426 154312
rect 422478 154300 422484 154312
rect 422536 154300 422542 154352
rect 145374 154272 145380 154284
rect 37976 154244 142752 154272
rect 142816 154244 145380 154272
rect 37976 154232 37982 154244
rect 27246 154164 27252 154216
rect 27304 154204 27310 154216
rect 137002 154204 137008 154216
rect 27304 154176 137008 154204
rect 27304 154164 27310 154176
rect 137002 154164 137008 154176
rect 137060 154164 137066 154216
rect 137112 154176 142568 154204
rect 23474 154096 23480 154148
rect 23532 154136 23538 154148
rect 136910 154136 136916 154148
rect 23532 154108 136916 154136
rect 23532 154096 23538 154108
rect 136910 154096 136916 154108
rect 136968 154096 136974 154148
rect 13814 154028 13820 154080
rect 13872 154068 13878 154080
rect 129182 154068 129188 154080
rect 13872 154040 129188 154068
rect 13872 154028 13878 154040
rect 129182 154028 129188 154040
rect 129240 154028 129246 154080
rect 137112 154068 137140 154176
rect 142430 154136 142436 154148
rect 129384 154040 137140 154068
rect 137204 154108 142436 154136
rect 9674 153960 9680 154012
rect 9732 154000 9738 154012
rect 126606 154000 126612 154012
rect 9732 153972 126612 154000
rect 9732 153960 9738 153972
rect 126606 153960 126612 153972
rect 126664 153960 126670 154012
rect 127618 153960 127624 154012
rect 127676 154000 127682 154012
rect 129274 154000 129280 154012
rect 127676 153972 129280 154000
rect 127676 153960 127682 153972
rect 129274 153960 129280 153972
rect 129332 153960 129338 154012
rect 7098 153892 7104 153944
rect 7156 153932 7162 153944
rect 124214 153932 124220 153944
rect 7156 153904 124220 153932
rect 7156 153892 7162 153904
rect 124214 153892 124220 153904
rect 124272 153892 124278 153944
rect 125502 153892 125508 153944
rect 125560 153932 125566 153944
rect 129384 153932 129412 154040
rect 129458 153960 129464 154012
rect 129516 154000 129522 154012
rect 137204 154000 137232 154108
rect 142430 154096 142436 154108
rect 142488 154096 142494 154148
rect 142540 154136 142568 154176
rect 142724 154136 142752 154244
rect 145374 154232 145380 154244
rect 145432 154232 145438 154284
rect 146938 154232 146944 154284
rect 146996 154272 147002 154284
rect 147950 154272 147956 154284
rect 146996 154244 147956 154272
rect 146996 154232 147002 154244
rect 147950 154232 147956 154244
rect 148008 154232 148014 154284
rect 148042 154232 148048 154284
rect 148100 154272 148106 154284
rect 156322 154272 156328 154284
rect 148100 154244 156328 154272
rect 148100 154232 148106 154244
rect 156322 154232 156328 154244
rect 156380 154232 156386 154284
rect 156782 154272 156788 154284
rect 156432 154244 156788 154272
rect 142890 154164 142896 154216
rect 142948 154204 142954 154216
rect 153286 154204 153292 154216
rect 142948 154176 153292 154204
rect 142948 154164 142954 154176
rect 153286 154164 153292 154176
rect 153344 154164 153350 154216
rect 156432 154204 156460 154244
rect 156782 154232 156788 154244
rect 156840 154232 156846 154284
rect 163222 154272 163228 154284
rect 161446 154244 163228 154272
rect 153396 154176 156460 154204
rect 147858 154136 147864 154148
rect 142540 154108 142660 154136
rect 142724 154108 147864 154136
rect 137278 154028 137284 154080
rect 137336 154068 137342 154080
rect 138014 154068 138020 154080
rect 137336 154040 138020 154068
rect 137336 154028 137342 154040
rect 138014 154028 138020 154040
rect 138072 154028 138078 154080
rect 142632 154068 142660 154108
rect 147858 154096 147864 154108
rect 147916 154096 147922 154148
rect 147950 154096 147956 154148
rect 148008 154136 148014 154148
rect 148008 154108 151814 154136
rect 148008 154096 148014 154108
rect 142982 154068 142988 154080
rect 142632 154040 142988 154068
rect 142982 154028 142988 154040
rect 143040 154028 143046 154080
rect 143442 154028 143448 154080
rect 143500 154068 143506 154080
rect 150434 154068 150440 154080
rect 143500 154040 150440 154068
rect 143500 154028 143506 154040
rect 150434 154028 150440 154040
rect 150492 154028 150498 154080
rect 151786 154068 151814 154108
rect 151906 154096 151912 154148
rect 151964 154136 151970 154148
rect 153396 154136 153424 154176
rect 156506 154164 156512 154216
rect 156564 154204 156570 154216
rect 161446 154204 161474 154244
rect 163222 154232 163228 154244
rect 163280 154232 163286 154284
rect 176654 154232 176660 154284
rect 176712 154272 176718 154284
rect 179506 154272 179512 154284
rect 176712 154244 179512 154272
rect 176712 154232 176718 154244
rect 179506 154232 179512 154244
rect 179564 154232 179570 154284
rect 182174 154232 182180 154284
rect 182232 154272 182238 154284
rect 258258 154272 258264 154284
rect 182232 154244 258264 154272
rect 182232 154232 182238 154244
rect 258258 154232 258264 154244
rect 258316 154232 258322 154284
rect 262214 154232 262220 154284
rect 262272 154272 262278 154284
rect 319254 154272 319260 154284
rect 262272 154244 319260 154272
rect 262272 154232 262278 154244
rect 319254 154232 319260 154244
rect 319312 154232 319318 154284
rect 343542 154232 343548 154284
rect 343600 154272 343606 154284
rect 380986 154272 380992 154284
rect 343600 154244 380992 154272
rect 343600 154232 343606 154244
rect 380986 154232 380992 154244
rect 381044 154232 381050 154284
rect 386506 154232 386512 154284
rect 386564 154272 386570 154284
rect 414198 154272 414204 154284
rect 386564 154244 414204 154272
rect 386564 154232 386570 154244
rect 414198 154232 414204 154244
rect 414256 154232 414262 154284
rect 156564 154176 161474 154204
rect 156564 154164 156570 154176
rect 162670 154164 162676 154216
rect 162728 154204 162734 154216
rect 165798 154204 165804 154216
rect 162728 154176 165804 154204
rect 162728 154164 162734 154176
rect 165798 154164 165804 154176
rect 165856 154164 165862 154216
rect 172514 154164 172520 154216
rect 172572 154204 172578 154216
rect 250530 154204 250536 154216
rect 172572 154176 250536 154204
rect 172572 154164 172578 154176
rect 250530 154164 250536 154176
rect 250588 154164 250594 154216
rect 255314 154164 255320 154216
rect 255372 154204 255378 154216
rect 314102 154204 314108 154216
rect 255372 154176 314108 154204
rect 255372 154164 255378 154176
rect 314102 154164 314108 154176
rect 314160 154164 314166 154216
rect 336826 154164 336832 154216
rect 336884 154204 336890 154216
rect 375742 154204 375748 154216
rect 336884 154176 375748 154204
rect 336884 154164 336890 154176
rect 375742 154164 375748 154176
rect 375800 154164 375806 154216
rect 383654 154164 383660 154216
rect 383712 154204 383718 154216
rect 411714 154204 411720 154216
rect 383712 154176 411720 154204
rect 383712 154164 383718 154176
rect 411714 154164 411720 154176
rect 411772 154164 411778 154216
rect 151964 154108 153424 154136
rect 151964 154096 151970 154108
rect 154942 154096 154948 154148
rect 155000 154136 155006 154148
rect 158070 154136 158076 154148
rect 155000 154108 158076 154136
rect 155000 154096 155006 154108
rect 158070 154096 158076 154108
rect 158128 154096 158134 154148
rect 160186 154096 160192 154148
rect 160244 154136 160250 154148
rect 160244 154108 162900 154136
rect 160244 154096 160250 154108
rect 162762 154068 162768 154080
rect 151786 154040 162768 154068
rect 162762 154028 162768 154040
rect 162820 154028 162826 154080
rect 162872 154068 162900 154108
rect 165614 154096 165620 154148
rect 165672 154136 165678 154148
rect 245654 154136 245660 154148
rect 165672 154108 245660 154136
rect 165672 154096 165678 154108
rect 245654 154096 245660 154108
rect 245712 154096 245718 154148
rect 245930 154096 245936 154148
rect 245988 154136 245994 154148
rect 306374 154136 306380 154148
rect 245988 154108 306380 154136
rect 245988 154096 245994 154108
rect 306374 154096 306380 154108
rect 306432 154096 306438 154148
rect 326706 154096 326712 154148
rect 326764 154136 326770 154148
rect 368014 154136 368020 154148
rect 326764 154108 368020 154136
rect 326764 154096 326770 154108
rect 368014 154096 368020 154108
rect 368072 154096 368078 154148
rect 376846 154096 376852 154148
rect 376904 154136 376910 154148
rect 406562 154136 406568 154148
rect 376904 154108 406568 154136
rect 376904 154096 376910 154108
rect 406562 154096 406568 154108
rect 406620 154096 406626 154148
rect 240962 154068 240968 154080
rect 162872 154040 240968 154068
rect 240962 154028 240968 154040
rect 241020 154028 241026 154080
rect 248598 154028 248604 154080
rect 248656 154068 248662 154080
rect 309226 154068 309232 154080
rect 248656 154040 309232 154068
rect 248656 154028 248662 154040
rect 309226 154028 309232 154040
rect 309284 154028 309290 154080
rect 323302 154028 323308 154080
rect 323360 154068 323366 154080
rect 365806 154068 365812 154080
rect 323360 154040 365812 154068
rect 323360 154028 323366 154040
rect 365806 154028 365812 154040
rect 365864 154028 365870 154080
rect 380158 154028 380164 154080
rect 380216 154068 380222 154080
rect 409138 154068 409144 154080
rect 380216 154040 409144 154068
rect 380216 154028 380222 154040
rect 409138 154028 409144 154040
rect 409196 154028 409202 154080
rect 219710 154000 219716 154012
rect 129516 153972 137232 154000
rect 137388 153972 138428 154000
rect 129516 153960 129522 153972
rect 125560 153904 129412 153932
rect 125560 153892 125566 153904
rect 132402 153892 132408 153944
rect 132460 153932 132466 153944
rect 137388 153932 137416 153972
rect 132460 153904 137416 153932
rect 132460 153892 132466 153904
rect 137462 153892 137468 153944
rect 137520 153932 137526 153944
rect 138400 153932 138428 153972
rect 143184 153972 219716 154000
rect 143184 153932 143212 153972
rect 219710 153960 219716 153972
rect 219768 153960 219774 154012
rect 222470 153960 222476 154012
rect 222528 154000 222534 154012
rect 288434 154000 288440 154012
rect 222528 153972 288440 154000
rect 222528 153960 222534 153972
rect 288434 153960 288440 153972
rect 288492 153960 288498 154012
rect 316034 153960 316040 154012
rect 316092 154000 316098 154012
rect 360378 154000 360384 154012
rect 316092 153972 360384 154000
rect 316092 153960 316098 153972
rect 360378 153960 360384 153972
rect 360436 153960 360442 154012
rect 367094 153960 367100 154012
rect 367152 154000 367158 154012
rect 398834 154000 398840 154012
rect 367152 153972 398840 154000
rect 367152 153960 367158 153972
rect 398834 153960 398840 153972
rect 398892 153960 398898 154012
rect 137520 153904 138336 153932
rect 138400 153904 143212 153932
rect 137520 153892 137526 153904
rect 474 153824 480 153876
rect 532 153864 538 153876
rect 119522 153864 119528 153876
rect 532 153836 119528 153864
rect 532 153824 538 153836
rect 119522 153824 119528 153836
rect 119580 153824 119586 153876
rect 119614 153824 119620 153876
rect 119672 153864 119678 153876
rect 138198 153864 138204 153876
rect 119672 153836 138204 153864
rect 119672 153824 119678 153836
rect 138198 153824 138204 153836
rect 138256 153824 138262 153876
rect 138308 153864 138336 153904
rect 143534 153892 143540 153944
rect 143592 153932 143598 153944
rect 145282 153932 145288 153944
rect 143592 153904 145288 153932
rect 143592 153892 143598 153904
rect 145282 153892 145288 153904
rect 145340 153892 145346 153944
rect 145374 153892 145380 153944
rect 145432 153932 145438 153944
rect 222930 153932 222936 153944
rect 145432 153904 222936 153932
rect 145432 153892 145438 153904
rect 222930 153892 222936 153904
rect 222988 153892 222994 153944
rect 225046 153892 225052 153944
rect 225104 153932 225110 153944
rect 291286 153932 291292 153944
rect 225104 153904 291292 153932
rect 225104 153892 225110 153904
rect 291286 153892 291292 153904
rect 291344 153892 291350 153944
rect 313274 153892 313280 153944
rect 313332 153932 313338 153944
rect 357802 153932 357808 153944
rect 313332 153904 357808 153932
rect 313332 153892 313338 153904
rect 357802 153892 357808 153904
rect 357860 153892 357866 153944
rect 363046 153892 363052 153944
rect 363104 153932 363110 153944
rect 396350 153932 396356 153944
rect 363104 153904 396356 153932
rect 363104 153892 363110 153904
rect 396350 153892 396356 153904
rect 396408 153892 396414 153944
rect 401594 153892 401600 153944
rect 401652 153932 401658 153944
rect 425330 153932 425336 153944
rect 401652 153904 425336 153932
rect 401652 153892 401658 153904
rect 425330 153892 425336 153904
rect 425388 153892 425394 153944
rect 138308 153836 156460 153864
rect 48314 153756 48320 153808
rect 48372 153796 48378 153808
rect 155494 153796 155500 153808
rect 48372 153768 155500 153796
rect 48372 153756 48378 153768
rect 155494 153756 155500 153768
rect 155552 153756 155558 153808
rect 156432 153796 156460 153836
rect 156782 153824 156788 153876
rect 156840 153864 156846 153876
rect 235166 153864 235172 153876
rect 156840 153836 235172 153864
rect 156840 153824 156846 153836
rect 235166 153824 235172 153836
rect 235224 153824 235230 153876
rect 241882 153824 241888 153876
rect 241940 153864 241946 153876
rect 303798 153864 303804 153876
rect 241940 153836 303804 153864
rect 241940 153824 241946 153836
rect 303798 153824 303804 153836
rect 303856 153824 303862 153876
rect 309134 153824 309140 153876
rect 309192 153864 309198 153876
rect 355226 153864 355232 153876
rect 309192 153836 355232 153864
rect 309192 153824 309198 153836
rect 355226 153824 355232 153836
rect 355284 153824 355290 153876
rect 356238 153824 356244 153876
rect 356296 153864 356302 153876
rect 391198 153864 391204 153876
rect 356296 153836 391204 153864
rect 356296 153824 356302 153836
rect 391198 153824 391204 153836
rect 391256 153824 391262 153876
rect 397454 153824 397460 153876
rect 397512 153864 397518 153876
rect 422662 153864 422668 153876
rect 397512 153836 422668 153864
rect 397512 153824 397518 153836
rect 422662 153824 422668 153836
rect 422720 153824 422726 153876
rect 191006 153796 191012 153808
rect 156432 153768 191012 153796
rect 191006 153756 191012 153768
rect 191064 153756 191070 153808
rect 191098 153756 191104 153808
rect 191156 153796 191162 153808
rect 197354 153796 197360 153808
rect 191156 153768 197360 153796
rect 191156 153756 191162 153768
rect 197354 153756 197360 153768
rect 197412 153756 197418 153808
rect 197446 153756 197452 153808
rect 197504 153796 197510 153808
rect 199286 153796 199292 153808
rect 197504 153768 199292 153796
rect 197504 153756 197510 153768
rect 199286 153756 199292 153768
rect 199344 153756 199350 153808
rect 210142 153796 210148 153808
rect 200408 153768 210148 153796
rect 61102 153688 61108 153740
rect 61160 153728 61166 153740
rect 162670 153728 162676 153740
rect 61160 153700 162676 153728
rect 61160 153688 61166 153700
rect 162670 153688 162676 153700
rect 162728 153688 162734 153740
rect 162762 153688 162768 153740
rect 162820 153728 162826 153740
rect 200408 153728 200436 153768
rect 210142 153756 210148 153768
rect 210200 153756 210206 153808
rect 231854 153756 231860 153808
rect 231912 153796 231918 153808
rect 296162 153796 296168 153808
rect 231912 153768 296168 153796
rect 231912 153756 231918 153768
rect 296162 153756 296168 153768
rect 296220 153756 296226 153808
rect 360470 153756 360476 153808
rect 360528 153796 360534 153808
rect 393774 153796 393780 153808
rect 360528 153768 393780 153796
rect 360528 153756 360534 153768
rect 393774 153756 393780 153768
rect 393832 153756 393838 153808
rect 427814 153756 427820 153808
rect 427872 153796 427878 153808
rect 432690 153796 432696 153808
rect 427872 153768 432696 153796
rect 427872 153756 427878 153768
rect 432690 153756 432696 153768
rect 432748 153756 432754 153808
rect 162820 153700 200436 153728
rect 162820 153688 162826 153700
rect 200482 153688 200488 153740
rect 200540 153728 200546 153740
rect 209774 153728 209780 153740
rect 200540 153700 209780 153728
rect 200540 153688 200546 153700
rect 209774 153688 209780 153700
rect 209832 153688 209838 153740
rect 235074 153688 235080 153740
rect 235132 153728 235138 153740
rect 298738 153728 298744 153740
rect 235132 153700 298744 153728
rect 235132 153688 235138 153700
rect 298738 153688 298744 153700
rect 298796 153688 298802 153740
rect 57974 153620 57980 153672
rect 58032 153660 58038 153672
rect 156506 153660 156512 153672
rect 58032 153632 156512 153660
rect 58032 153620 58038 153632
rect 156506 153620 156512 153632
rect 156564 153620 156570 153672
rect 156690 153620 156696 153672
rect 156748 153660 156754 153672
rect 218054 153660 218060 153672
rect 156748 153632 218060 153660
rect 156748 153620 156754 153632
rect 218054 153620 218060 153632
rect 218112 153620 218118 153672
rect 229094 153620 229100 153672
rect 229152 153660 229158 153672
rect 293586 153660 293592 153672
rect 229152 153632 293592 153660
rect 229152 153620 229158 153632
rect 293586 153620 293592 153632
rect 293644 153620 293650 153672
rect 78674 153552 78680 153604
rect 78732 153592 78738 153604
rect 179414 153592 179420 153604
rect 78732 153564 179420 153592
rect 78732 153552 78738 153564
rect 179414 153552 179420 153564
rect 179472 153552 179478 153604
rect 179506 153552 179512 153604
rect 179564 153592 179570 153604
rect 230658 153592 230664 153604
rect 179564 153564 230664 153592
rect 179564 153552 179570 153564
rect 230658 153552 230664 153564
rect 230716 153552 230722 153604
rect 238846 153552 238852 153604
rect 238904 153592 238910 153604
rect 301314 153592 301320 153604
rect 238904 153564 301320 153592
rect 238904 153552 238910 153564
rect 301314 153552 301320 153564
rect 301372 153552 301378 153604
rect 102134 153484 102140 153536
rect 102192 153524 102198 153536
rect 196618 153524 196624 153536
rect 102192 153496 196624 153524
rect 102192 153484 102198 153496
rect 196618 153484 196624 153496
rect 196676 153484 196682 153536
rect 198918 153484 198924 153536
rect 198976 153524 198982 153536
rect 248598 153524 248604 153536
rect 198976 153496 248604 153524
rect 198976 153484 198982 153496
rect 248598 153484 248604 153496
rect 248656 153484 248662 153536
rect 252646 153484 252652 153536
rect 252704 153524 252710 153536
rect 311526 153524 311532 153536
rect 252704 153496 311532 153524
rect 252704 153484 252710 153496
rect 311526 153484 311532 153496
rect 311584 153484 311590 153536
rect 104894 153416 104900 153468
rect 104952 153456 104958 153468
rect 199194 153456 199200 153468
rect 104952 153428 199200 153456
rect 104952 153416 104958 153428
rect 199194 153416 199200 153428
rect 199252 153416 199258 153468
rect 199286 153416 199292 153468
rect 199344 153456 199350 153468
rect 199344 153428 200528 153456
rect 199344 153416 199350 153428
rect 108298 153348 108304 153400
rect 108356 153388 108362 153400
rect 191282 153388 191288 153400
rect 108356 153360 191288 153388
rect 108356 153348 108362 153360
rect 191282 153348 191288 153360
rect 191340 153348 191346 153400
rect 191742 153348 191748 153400
rect 191800 153388 191806 153400
rect 200114 153388 200120 153400
rect 191800 153360 200120 153388
rect 191800 153348 191806 153360
rect 200114 153348 200120 153360
rect 200172 153348 200178 153400
rect 115934 153280 115940 153332
rect 115992 153320 115998 153332
rect 200500 153320 200528 153428
rect 200574 153416 200580 153468
rect 200632 153456 200638 153468
rect 258902 153456 258908 153468
rect 200632 153428 258908 153456
rect 200632 153416 200638 153428
rect 258902 153416 258908 153428
rect 258960 153416 258966 153468
rect 265434 153416 265440 153468
rect 265492 153456 265498 153468
rect 321830 153456 321836 153468
rect 265492 153428 321836 153456
rect 265492 153416 265498 153428
rect 321830 153416 321836 153428
rect 321888 153416 321894 153468
rect 243446 153388 243452 153400
rect 200776 153360 243452 153388
rect 200776 153320 200804 153360
rect 243446 153348 243452 153360
rect 243504 153348 243510 153400
rect 259454 153348 259460 153400
rect 259512 153388 259518 153400
rect 316770 153388 316776 153400
rect 259512 153360 316776 153388
rect 259512 153348 259518 153360
rect 316770 153348 316776 153360
rect 316828 153348 316834 153400
rect 441614 153348 441620 153400
rect 441672 153388 441678 153400
rect 441672 153360 441936 153388
rect 441672 153348 441678 153360
rect 115992 153292 200436 153320
rect 200500 153292 200804 153320
rect 115992 153280 115998 153292
rect 41598 153212 41604 153264
rect 41656 153252 41662 153264
rect 138106 153252 138112 153264
rect 41656 153224 138112 153252
rect 41656 153212 41662 153224
rect 138106 153212 138112 153224
rect 138164 153212 138170 153264
rect 138198 153212 138204 153264
rect 138256 153252 138262 153264
rect 200298 153252 200304 153264
rect 138256 153224 200304 153252
rect 138256 153212 138262 153224
rect 200298 153212 200304 153224
rect 200356 153212 200362 153264
rect 200408 153252 200436 153292
rect 200850 153280 200856 153332
rect 200908 153320 200914 153332
rect 238386 153320 238392 153332
rect 200908 153292 238392 153320
rect 200908 153280 200914 153292
rect 238386 153280 238392 153292
rect 238444 153280 238450 153332
rect 272886 153280 272892 153332
rect 272944 153320 272950 153332
rect 327074 153320 327080 153332
rect 272944 153292 327080 153320
rect 272944 153280 272950 153292
rect 327074 153280 327080 153292
rect 327132 153280 327138 153332
rect 207566 153252 207572 153264
rect 200408 153224 207572 153252
rect 207566 153212 207572 153224
rect 207624 153212 207630 153264
rect 269206 153212 269212 153264
rect 269264 153252 269270 153264
rect 324406 153252 324412 153264
rect 269264 153224 324412 153252
rect 269264 153212 269270 153224
rect 324406 153212 324412 153224
rect 324464 153212 324470 153264
rect 423582 153212 423588 153264
rect 423640 153252 423646 153264
rect 427998 153252 428004 153264
rect 423640 153224 428004 153252
rect 423640 153212 423646 153224
rect 427998 153212 428004 153224
rect 428056 153212 428062 153264
rect 23290 153144 23296 153196
rect 23348 153184 23354 153196
rect 110966 153184 110972 153196
rect 23348 153156 110972 153184
rect 23348 153144 23354 153156
rect 110966 153144 110972 153156
rect 111024 153144 111030 153196
rect 113174 153144 113180 153196
rect 113232 153184 113238 153196
rect 205634 153184 205640 153196
rect 113232 153156 205640 153184
rect 113232 153144 113238 153156
rect 205634 153144 205640 153156
rect 205692 153144 205698 153196
rect 215386 153144 215392 153196
rect 215444 153184 215450 153196
rect 279418 153184 279424 153196
rect 215444 153156 279424 153184
rect 215444 153144 215450 153156
rect 279418 153144 279424 153156
rect 279476 153144 279482 153196
rect 285490 153144 285496 153196
rect 285548 153184 285554 153196
rect 336734 153184 336740 153196
rect 285548 153156 336740 153184
rect 285548 153144 285554 153156
rect 336734 153144 336740 153156
rect 336792 153144 336798 153196
rect 339678 153144 339684 153196
rect 339736 153184 339742 153196
rect 377030 153184 377036 153196
rect 339736 153156 377036 153184
rect 339736 153144 339742 153156
rect 377030 153144 377036 153156
rect 377088 153144 377094 153196
rect 385402 153144 385408 153196
rect 385460 153184 385466 153196
rect 387334 153184 387340 153196
rect 385460 153156 387340 153184
rect 385460 153144 385466 153156
rect 387334 153144 387340 153156
rect 387392 153144 387398 153196
rect 389174 153144 389180 153196
rect 389232 153184 389238 153196
rect 412634 153184 412640 153196
rect 389232 153156 412640 153184
rect 389232 153144 389238 153156
rect 412634 153144 412640 153156
rect 412692 153144 412698 153196
rect 413094 153144 413100 153196
rect 413152 153184 413158 153196
rect 433426 153184 433432 153196
rect 413152 153156 433432 153184
rect 413152 153144 413158 153156
rect 433426 153144 433432 153156
rect 433484 153144 433490 153196
rect 433518 153144 433524 153196
rect 433576 153184 433582 153196
rect 441798 153184 441804 153196
rect 433576 153156 441804 153184
rect 433576 153144 433582 153156
rect 441798 153144 441804 153156
rect 441856 153144 441862 153196
rect 441908 153184 441936 153360
rect 442920 153224 444052 153252
rect 442920 153184 442948 153224
rect 441908 153156 442948 153184
rect 442994 153144 443000 153196
rect 443052 153184 443058 153196
rect 443914 153184 443920 153196
rect 443052 153156 443920 153184
rect 443052 153144 443058 153156
rect 443914 153144 443920 153156
rect 443972 153144 443978 153196
rect 444024 153184 444052 153224
rect 450262 153184 450268 153196
rect 444024 153156 450268 153184
rect 450262 153144 450268 153156
rect 450320 153144 450326 153196
rect 456794 153144 456800 153196
rect 456852 153184 456858 153196
rect 459186 153184 459192 153196
rect 456852 153156 459192 153184
rect 456852 153144 456858 153156
rect 459186 153144 459192 153156
rect 459244 153144 459250 153196
rect 461486 153144 461492 153196
rect 461544 153184 461550 153196
rect 463050 153184 463056 153196
rect 461544 153156 463056 153184
rect 461544 153144 461550 153156
rect 463050 153144 463056 153156
rect 463108 153144 463114 153196
rect 466454 153144 466460 153196
rect 466512 153184 466518 153196
rect 469490 153184 469496 153196
rect 466512 153156 469496 153184
rect 466512 153144 466518 153156
rect 469490 153144 469496 153156
rect 469548 153144 469554 153196
rect 471238 153144 471244 153196
rect 471296 153184 471302 153196
rect 473538 153184 473544 153196
rect 471296 153156 473544 153184
rect 471296 153144 471302 153156
rect 473538 153144 473544 153156
rect 473596 153144 473602 153196
rect 474826 153144 474832 153196
rect 474884 153184 474890 153196
rect 476574 153184 476580 153196
rect 474884 153156 476580 153184
rect 474884 153144 474890 153156
rect 476574 153144 476580 153156
rect 476632 153144 476638 153196
rect 485682 153144 485688 153196
rect 485740 153184 485746 153196
rect 489362 153184 489368 153196
rect 485740 153156 489368 153184
rect 485740 153144 485746 153156
rect 489362 153144 489368 153156
rect 489420 153144 489426 153196
rect 490742 153144 490748 153196
rect 490800 153184 490806 153196
rect 493226 153184 493232 153196
rect 490800 153156 493232 153184
rect 490800 153144 490806 153156
rect 493226 153144 493232 153156
rect 493284 153144 493290 153196
rect 494146 153144 494152 153196
rect 494204 153184 494210 153196
rect 496446 153184 496452 153196
rect 494204 153156 496452 153184
rect 494204 153144 494210 153156
rect 496446 153144 496452 153156
rect 496504 153144 496510 153196
rect 496630 153144 496636 153196
rect 496688 153184 496694 153196
rect 497734 153184 497740 153196
rect 496688 153156 497740 153184
rect 496688 153144 496694 153156
rect 497734 153144 497740 153156
rect 497792 153144 497798 153196
rect 512546 153144 512552 153196
rect 512604 153184 512610 153196
rect 514846 153184 514852 153196
rect 512604 153156 514852 153184
rect 512604 153144 512610 153156
rect 514846 153144 514852 153156
rect 514904 153144 514910 153196
rect 80054 153076 80060 153128
rect 80112 153116 80118 153128
rect 174814 153116 174820 153128
rect 80112 153088 174820 153116
rect 80112 153076 80118 153088
rect 174814 153076 174820 153088
rect 174872 153076 174878 153128
rect 180794 153076 180800 153128
rect 180852 153116 180858 153128
rect 256970 153116 256976 153128
rect 180852 153088 256976 153116
rect 180852 153076 180858 153088
rect 256970 153076 256976 153088
rect 257028 153076 257034 153128
rect 264974 153076 264980 153128
rect 265032 153116 265038 153128
rect 321186 153116 321192 153128
rect 265032 153088 321192 153116
rect 265032 153076 265038 153088
rect 321186 153076 321192 153088
rect 321244 153076 321250 153128
rect 324314 153076 324320 153128
rect 324372 153116 324378 153128
rect 366726 153116 366732 153128
rect 324372 153088 366732 153116
rect 324372 153076 324378 153088
rect 366726 153076 366732 153088
rect 366784 153076 366790 153128
rect 382182 153076 382188 153128
rect 382240 153116 382246 153128
rect 410426 153116 410432 153128
rect 382240 153088 410432 153116
rect 382240 153076 382246 153088
rect 410426 153076 410432 153088
rect 410484 153076 410490 153128
rect 414290 153076 414296 153128
rect 414348 153116 414354 153128
rect 414348 153088 430620 153116
rect 414348 153076 414354 153088
rect 103514 153008 103520 153060
rect 103572 153048 103578 153060
rect 197906 153048 197912 153060
rect 103572 153020 197912 153048
rect 103572 153008 103578 153020
rect 197906 153008 197912 153020
rect 197964 153008 197970 153060
rect 203702 153008 203708 153060
rect 203760 153048 203766 153060
rect 267274 153048 267280 153060
rect 203760 153020 267280 153048
rect 203760 153008 203766 153020
rect 267274 153008 267280 153020
rect 267332 153008 267338 153060
rect 272150 153008 272156 153060
rect 272208 153048 272214 153060
rect 326338 153048 326344 153060
rect 272208 153020 326344 153048
rect 272208 153008 272214 153020
rect 326338 153008 326344 153020
rect 326396 153008 326402 153060
rect 330938 153008 330944 153060
rect 330996 153048 331002 153060
rect 371234 153048 371240 153060
rect 330996 153020 371240 153048
rect 330996 153008 331002 153020
rect 371234 153008 371240 153020
rect 371292 153008 371298 153060
rect 372614 153008 372620 153060
rect 372672 153048 372678 153060
rect 403342 153048 403348 153060
rect 372672 153020 403348 153048
rect 372672 153008 372678 153020
rect 403342 153008 403348 153020
rect 403400 153008 403406 153060
rect 404354 153008 404360 153060
rect 404412 153048 404418 153060
rect 427906 153048 427912 153060
rect 404412 153020 427912 153048
rect 404412 153008 404418 153020
rect 427906 153008 427912 153020
rect 427964 153008 427970 153060
rect 430592 153048 430620 153088
rect 430666 153076 430672 153128
rect 430724 153116 430730 153128
rect 436278 153116 436284 153128
rect 430724 153088 436284 153116
rect 430724 153076 430730 153088
rect 436278 153076 436284 153088
rect 436336 153076 436342 153128
rect 436922 153076 436928 153128
rect 436980 153116 436986 153128
rect 452194 153116 452200 153128
rect 436980 153088 452200 153116
rect 436980 153076 436986 153088
rect 452194 153076 452200 153088
rect 452252 153076 452258 153128
rect 466546 153076 466552 153128
rect 466604 153116 466610 153128
rect 470134 153116 470140 153128
rect 466604 153088 470140 153116
rect 466604 153076 466610 153088
rect 470134 153076 470140 153088
rect 470192 153076 470198 153128
rect 471514 153076 471520 153128
rect 471572 153116 471578 153128
rect 472710 153116 472716 153128
rect 471572 153088 472716 153116
rect 471572 153076 471578 153088
rect 472710 153076 472716 153088
rect 472768 153076 472774 153128
rect 473354 153076 473360 153128
rect 473412 153116 473418 153128
rect 475286 153116 475292 153128
rect 473412 153088 475292 153116
rect 473412 153076 473418 153088
rect 475286 153076 475292 153088
rect 475344 153076 475350 153128
rect 476114 153076 476120 153128
rect 476172 153116 476178 153128
rect 477862 153116 477868 153128
rect 476172 153088 477868 153116
rect 476172 153076 476178 153088
rect 477862 153076 477868 153088
rect 477920 153076 477926 153128
rect 484026 153076 484032 153128
rect 484084 153116 484090 153128
rect 488074 153116 488080 153128
rect 484084 153088 488080 153116
rect 484084 153076 484090 153088
rect 488074 153076 488080 153088
rect 488132 153076 488138 153128
rect 489914 153076 489920 153128
rect 489972 153116 489978 153128
rect 492766 153116 492772 153128
rect 489972 153088 492772 153116
rect 489972 153076 489978 153088
rect 492766 153076 492772 153088
rect 492824 153076 492830 153128
rect 494054 153076 494060 153128
rect 494112 153116 494118 153128
rect 495802 153116 495808 153128
rect 494112 153088 495808 153116
rect 494112 153076 494118 153088
rect 495802 153076 495808 153088
rect 495860 153076 495866 153128
rect 496814 153076 496820 153128
rect 496872 153116 496878 153128
rect 498378 153116 498384 153128
rect 496872 153088 498384 153116
rect 496872 153076 496878 153088
rect 498378 153076 498384 153088
rect 498436 153076 498442 153128
rect 511258 153076 511264 153128
rect 511316 153116 511322 153128
rect 513466 153116 513472 153128
rect 511316 153088 513472 153116
rect 511316 153076 511322 153088
rect 513466 153076 513472 153088
rect 513524 153076 513530 153128
rect 514478 153076 514484 153128
rect 514536 153116 514542 153128
rect 517422 153116 517428 153128
rect 514536 153088 517428 153116
rect 514536 153076 514542 153088
rect 517422 153076 517428 153088
rect 517480 153076 517486 153128
rect 431862 153048 431868 153060
rect 430592 153020 431868 153048
rect 431862 153008 431868 153020
rect 431920 153008 431926 153060
rect 431954 153008 431960 153060
rect 432012 153048 432018 153060
rect 448974 153048 448980 153060
rect 432012 153020 448980 153048
rect 432012 153008 432018 153020
rect 448974 153008 448980 153020
rect 449032 153008 449038 153060
rect 465074 153008 465080 153060
rect 465132 153048 465138 153060
rect 468846 153048 468852 153060
rect 465132 153020 468852 153048
rect 465132 153008 465138 153020
rect 468846 153008 468852 153020
rect 468904 153008 468910 153060
rect 472434 153008 472440 153060
rect 472492 153048 472498 153060
rect 474734 153048 474740 153060
rect 472492 153020 474740 153048
rect 472492 153008 472498 153020
rect 474734 153008 474740 153020
rect 474792 153008 474798 153060
rect 484486 153008 484492 153060
rect 484544 153048 484550 153060
rect 488718 153048 488724 153060
rect 484544 153020 488724 153048
rect 484544 153008 484550 153020
rect 488718 153008 488724 153020
rect 488776 153008 488782 153060
rect 492674 153008 492680 153060
rect 492732 153048 492738 153060
rect 495434 153048 495440 153060
rect 492732 153020 495440 153048
rect 492732 153008 492738 153020
rect 495434 153008 495440 153020
rect 495492 153008 495498 153060
rect 495526 153008 495532 153060
rect 495584 153048 495590 153060
rect 497090 153048 497096 153060
rect 495584 153020 497096 153048
rect 495584 153008 495590 153020
rect 497090 153008 497096 153020
rect 497148 153008 497154 153060
rect 511718 153008 511724 153060
rect 511776 153048 511782 153060
rect 514294 153048 514300 153060
rect 511776 153020 514300 153048
rect 511776 153008 511782 153020
rect 514294 153008 514300 153020
rect 514352 153008 514358 153060
rect 92566 152940 92572 152992
rect 92624 152980 92630 152992
rect 187694 152980 187700 152992
rect 92624 152952 187700 152980
rect 92624 152940 92630 152952
rect 187694 152940 187700 152952
rect 187752 152940 187758 152992
rect 195422 152940 195428 152992
rect 195480 152980 195486 152992
rect 218422 152980 218428 152992
rect 195480 152952 218428 152980
rect 195480 152940 195486 152952
rect 218422 152940 218428 152952
rect 218480 152940 218486 152992
rect 225230 152940 225236 152992
rect 225288 152980 225294 152992
rect 228726 152980 228732 152992
rect 225288 152952 228732 152980
rect 225288 152940 225294 152952
rect 228726 152940 228732 152952
rect 228784 152940 228790 152992
rect 228818 152940 228824 152992
rect 228876 152980 228882 152992
rect 284570 152980 284576 152992
rect 228876 152952 284576 152980
rect 228876 152940 228882 152952
rect 284570 152940 284576 152952
rect 284628 152940 284634 152992
rect 288158 152940 288164 152992
rect 288216 152980 288222 152992
rect 289906 152980 289912 152992
rect 288216 152952 289912 152980
rect 288216 152940 288222 152952
rect 289906 152940 289912 152952
rect 289964 152940 289970 152992
rect 291378 152940 291384 152992
rect 291436 152980 291442 152992
rect 341058 152980 341064 152992
rect 291436 152952 341064 152980
rect 291436 152940 291442 152952
rect 341058 152940 341064 152952
rect 341116 152940 341122 152992
rect 342254 152940 342260 152992
rect 342312 152980 342318 152992
rect 344278 152980 344284 152992
rect 342312 152952 344284 152980
rect 342312 152940 342318 152952
rect 344278 152940 344284 152952
rect 344336 152940 344342 152992
rect 345290 152940 345296 152992
rect 345348 152980 345354 152992
rect 382274 152980 382280 152992
rect 345348 152952 382280 152980
rect 345348 152940 345354 152952
rect 382274 152940 382280 152952
rect 382332 152940 382338 152992
rect 382366 152940 382372 152992
rect 382424 152980 382430 152992
rect 386690 152980 386696 152992
rect 382424 152952 386696 152980
rect 382424 152940 382430 152952
rect 386690 152940 386696 152952
rect 386748 152940 386754 152992
rect 390370 152940 390376 152992
rect 390428 152980 390434 152992
rect 414934 152980 414940 152992
rect 390428 152952 414940 152980
rect 390428 152940 390434 152952
rect 414934 152940 414940 152952
rect 414992 152940 414998 152992
rect 418154 152940 418160 152992
rect 418212 152980 418218 152992
rect 432874 152980 432880 152992
rect 418212 152952 432880 152980
rect 418212 152940 418218 152952
rect 432874 152940 432880 152952
rect 432932 152940 432938 152992
rect 438854 152940 438860 152992
rect 438912 152980 438918 152992
rect 454218 152980 454224 152992
rect 438912 152952 454224 152980
rect 438912 152940 438918 152952
rect 454218 152940 454224 152952
rect 454276 152940 454282 152992
rect 472250 152940 472256 152992
rect 472308 152980 472314 152992
rect 473998 152980 474004 152992
rect 472308 152952 474004 152980
rect 472308 152940 472314 152952
rect 473998 152940 474004 152952
rect 474056 152940 474062 152992
rect 483198 152940 483204 152992
rect 483256 152980 483262 152992
rect 487522 152980 487528 152992
rect 483256 152952 487528 152980
rect 483256 152940 483262 152952
rect 487522 152940 487528 152952
rect 487580 152940 487586 152992
rect 491294 152940 491300 152992
rect 491352 152980 491358 152992
rect 494054 152980 494060 152992
rect 491352 152952 494060 152980
rect 491352 152940 491358 152952
rect 494054 152940 494060 152952
rect 494112 152940 494118 152992
rect 513190 152940 513196 152992
rect 513248 152980 513254 152992
rect 515950 152980 515956 152992
rect 513248 152952 515956 152980
rect 513248 152940 513254 152952
rect 515950 152940 515956 152952
rect 516008 152940 516014 152992
rect 71406 152872 71412 152924
rect 71464 152912 71470 152924
rect 92474 152912 92480 152924
rect 71464 152884 92480 152912
rect 71464 152872 71470 152884
rect 92474 152872 92480 152884
rect 92532 152872 92538 152924
rect 96614 152872 96620 152924
rect 96672 152912 96678 152924
rect 192754 152912 192760 152924
rect 96672 152884 192760 152912
rect 96672 152872 96678 152884
rect 192754 152872 192760 152884
rect 192812 152872 192818 152924
rect 212442 152872 212448 152924
rect 212500 152912 212506 152924
rect 277486 152912 277492 152924
rect 212500 152884 277492 152912
rect 212500 152872 212506 152884
rect 277486 152872 277492 152884
rect 277544 152872 277550 152924
rect 278774 152872 278780 152924
rect 278832 152912 278838 152924
rect 331490 152912 331496 152924
rect 278832 152884 331496 152912
rect 278832 152872 278838 152884
rect 331490 152872 331496 152884
rect 331548 152872 331554 152924
rect 332594 152872 332600 152924
rect 332652 152912 332658 152924
rect 372614 152912 372620 152924
rect 332652 152884 372620 152912
rect 332652 152872 332658 152884
rect 372614 152872 372620 152884
rect 372672 152872 372678 152924
rect 375466 152872 375472 152924
rect 375524 152912 375530 152924
rect 405274 152912 405280 152924
rect 375524 152884 405280 152912
rect 375524 152872 375530 152884
rect 405274 152872 405280 152884
rect 405332 152872 405338 152924
rect 405918 152872 405924 152924
rect 405976 152912 405982 152924
rect 408494 152912 408500 152924
rect 405976 152884 408500 152912
rect 405976 152872 405982 152884
rect 408494 152872 408500 152884
rect 408552 152872 408558 152924
rect 411254 152872 411260 152924
rect 411312 152912 411318 152924
rect 432598 152912 432604 152924
rect 411312 152884 432604 152912
rect 411312 152872 411318 152884
rect 432598 152872 432604 152884
rect 432656 152872 432662 152924
rect 434346 152872 434352 152924
rect 434404 152912 434410 152924
rect 441614 152912 441620 152924
rect 434404 152884 441620 152912
rect 434404 152872 434410 152884
rect 441614 152872 441620 152884
rect 441672 152872 441678 152924
rect 441706 152872 441712 152924
rect 441764 152912 441770 152924
rect 447870 152912 447876 152924
rect 441764 152884 447876 152912
rect 441764 152872 441770 152884
rect 447870 152872 447876 152884
rect 447928 152872 447934 152924
rect 491662 152872 491668 152924
rect 491720 152912 491726 152924
rect 494514 152912 494520 152924
rect 491720 152884 494520 152912
rect 491720 152872 491726 152884
rect 494514 152872 494520 152884
rect 494572 152872 494578 152924
rect 513834 152872 513840 152924
rect 513892 152912 513898 152924
rect 516134 152912 516140 152924
rect 513892 152884 516140 152912
rect 513892 152872 513898 152884
rect 516134 152872 516140 152884
rect 516192 152872 516198 152924
rect 33134 152804 33140 152856
rect 33192 152844 33198 152856
rect 138290 152844 138296 152856
rect 33192 152816 138296 152844
rect 33192 152804 33198 152816
rect 138290 152804 138296 152816
rect 138348 152804 138354 152856
rect 138566 152804 138572 152856
rect 138624 152844 138630 152856
rect 141418 152844 141424 152856
rect 138624 152816 141424 152844
rect 138624 152804 138630 152816
rect 141418 152804 141424 152816
rect 141476 152804 141482 152856
rect 146478 152804 146484 152856
rect 146536 152844 146542 152856
rect 167086 152844 167092 152856
rect 146536 152816 167092 152844
rect 146536 152804 146542 152816
rect 167086 152804 167092 152816
rect 167144 152804 167150 152856
rect 173894 152804 173900 152856
rect 173952 152844 173958 152856
rect 251818 152844 251824 152856
rect 173952 152816 251824 152844
rect 173952 152804 173958 152816
rect 251818 152804 251824 152816
rect 251876 152804 251882 152856
rect 255406 152804 255412 152856
rect 255464 152844 255470 152856
rect 312814 152844 312820 152856
rect 255464 152816 312820 152844
rect 255464 152804 255470 152816
rect 312814 152804 312820 152816
rect 312872 152804 312878 152856
rect 316310 152804 316316 152856
rect 316368 152844 316374 152856
rect 317966 152844 317972 152856
rect 316368 152816 317972 152844
rect 316368 152804 316374 152816
rect 317966 152804 317972 152816
rect 318024 152804 318030 152856
rect 361022 152844 361028 152856
rect 318076 152816 361028 152844
rect 26418 152736 26424 152788
rect 26476 152776 26482 152788
rect 138842 152776 138848 152788
rect 26476 152748 138848 152776
rect 26476 152736 26482 152748
rect 138842 152736 138848 152748
rect 138900 152736 138906 152788
rect 140866 152736 140872 152788
rect 140924 152776 140930 152788
rect 143994 152776 144000 152788
rect 140924 152748 144000 152776
rect 140924 152736 140930 152748
rect 143994 152736 144000 152748
rect 144052 152736 144058 152788
rect 144086 152736 144092 152788
rect 144144 152776 144150 152788
rect 161934 152776 161940 152788
rect 144144 152748 161940 152776
rect 144144 152736 144150 152748
rect 161934 152736 161940 152748
rect 161992 152736 161998 152788
rect 164326 152736 164332 152788
rect 164384 152776 164390 152788
rect 244274 152776 244280 152788
rect 164384 152748 244280 152776
rect 164384 152736 164390 152748
rect 244274 152736 244280 152748
rect 244332 152736 244338 152788
rect 257706 152736 257712 152788
rect 257764 152776 257770 152788
rect 315390 152776 315396 152788
rect 257764 152748 315396 152776
rect 257764 152736 257770 152748
rect 315390 152736 315396 152748
rect 315448 152736 315454 152788
rect 317414 152736 317420 152788
rect 317472 152776 317478 152788
rect 318076 152776 318104 152816
rect 361022 152804 361028 152816
rect 361080 152804 361086 152856
rect 361574 152804 361580 152856
rect 361632 152844 361638 152856
rect 395062 152844 395068 152856
rect 361632 152816 395068 152844
rect 361632 152804 361638 152816
rect 395062 152804 395068 152816
rect 395120 152804 395126 152856
rect 395430 152804 395436 152856
rect 395488 152844 395494 152856
rect 397546 152844 397552 152856
rect 395488 152816 397552 152844
rect 395488 152804 395494 152816
rect 397546 152804 397552 152816
rect 397604 152804 397610 152856
rect 406654 152804 406660 152856
rect 406712 152844 406718 152856
rect 429194 152844 429200 152856
rect 406712 152816 429200 152844
rect 406712 152804 406718 152816
rect 429194 152804 429200 152816
rect 429252 152804 429258 152856
rect 429378 152804 429384 152856
rect 429436 152844 429442 152856
rect 447134 152844 447140 152856
rect 429436 152816 447140 152844
rect 429436 152804 429442 152816
rect 447134 152804 447140 152816
rect 447192 152804 447198 152856
rect 317472 152748 318104 152776
rect 317472 152736 317478 152748
rect 320266 152736 320272 152788
rect 320324 152776 320330 152788
rect 323118 152776 323124 152788
rect 320324 152748 323124 152776
rect 320324 152736 320330 152748
rect 323118 152736 323124 152748
rect 323176 152736 323182 152788
rect 324222 152736 324228 152788
rect 324280 152776 324286 152788
rect 366082 152776 366088 152788
rect 324280 152748 366088 152776
rect 324280 152736 324286 152748
rect 366082 152736 366088 152748
rect 366140 152736 366146 152788
rect 368474 152736 368480 152788
rect 368532 152776 368538 152788
rect 400214 152776 400220 152788
rect 368532 152748 400220 152776
rect 368532 152736 368538 152748
rect 400214 152736 400220 152748
rect 400272 152736 400278 152788
rect 402422 152736 402428 152788
rect 402480 152776 402486 152788
rect 425882 152776 425888 152788
rect 402480 152748 425888 152776
rect 402480 152736 402486 152748
rect 425882 152736 425888 152748
rect 425940 152736 425946 152788
rect 426434 152736 426440 152788
rect 426492 152776 426498 152788
rect 444558 152776 444564 152788
rect 426492 152748 444564 152776
rect 426492 152736 426498 152748
rect 444558 152736 444564 152748
rect 444616 152736 444622 152788
rect 446306 152736 446312 152788
rect 446364 152776 446370 152788
rect 459830 152776 459836 152788
rect 446364 152748 459836 152776
rect 446364 152736 446370 152748
rect 459830 152736 459836 152748
rect 459888 152736 459894 152788
rect 510522 152736 510528 152788
rect 510580 152776 510586 152788
rect 511994 152776 512000 152788
rect 510580 152748 512000 152776
rect 510580 152736 510586 152748
rect 511994 152736 512000 152748
rect 512052 152736 512058 152788
rect 28166 152668 28172 152720
rect 28224 152708 28230 152720
rect 140774 152708 140780 152720
rect 28224 152680 140780 152708
rect 28224 152668 28230 152680
rect 140774 152668 140780 152680
rect 140832 152668 140838 152720
rect 142798 152668 142804 152720
rect 142856 152708 142862 152720
rect 149146 152708 149152 152720
rect 142856 152680 149152 152708
rect 142856 152668 142862 152680
rect 149146 152668 149152 152680
rect 149204 152668 149210 152720
rect 149330 152668 149336 152720
rect 149388 152708 149394 152720
rect 231302 152708 231308 152720
rect 149388 152680 231308 152708
rect 149388 152668 149394 152680
rect 231302 152668 231308 152680
rect 231360 152668 231366 152720
rect 251174 152668 251180 152720
rect 251232 152708 251238 152720
rect 310882 152708 310888 152720
rect 251232 152680 310888 152708
rect 251232 152668 251238 152680
rect 310882 152668 310888 152680
rect 310940 152668 310946 152720
rect 311986 152668 311992 152720
rect 312044 152708 312050 152720
rect 356054 152708 356060 152720
rect 312044 152680 356060 152708
rect 312044 152668 312050 152680
rect 356054 152668 356060 152680
rect 356112 152668 356118 152720
rect 358814 152668 358820 152720
rect 358872 152708 358878 152720
rect 393314 152708 393320 152720
rect 358872 152680 393320 152708
rect 358872 152668 358878 152680
rect 393314 152668 393320 152680
rect 393372 152668 393378 152720
rect 394878 152668 394884 152720
rect 394936 152708 394942 152720
rect 420086 152708 420092 152720
rect 394936 152680 420092 152708
rect 394936 152668 394942 152680
rect 420086 152668 420092 152680
rect 420144 152668 420150 152720
rect 421006 152668 421012 152720
rect 421064 152708 421070 152720
rect 421064 152680 432598 152708
rect 421064 152668 421070 152680
rect 22186 152600 22192 152652
rect 22244 152640 22250 152652
rect 135622 152640 135628 152652
rect 22244 152612 135628 152640
rect 22244 152600 22250 152612
rect 135622 152600 135628 152612
rect 135680 152600 135686 152652
rect 151814 152640 151820 152652
rect 137986 152612 151820 152640
rect 19334 152532 19340 152584
rect 19392 152572 19398 152584
rect 133874 152572 133880 152584
rect 19392 152544 133880 152572
rect 19392 152532 19398 152544
rect 133874 152532 133880 152544
rect 133932 152532 133938 152584
rect 136818 152532 136824 152584
rect 136876 152572 136882 152584
rect 137986 152572 138014 152612
rect 151814 152600 151820 152612
rect 151872 152600 151878 152652
rect 153654 152600 153660 152652
rect 153712 152640 153718 152652
rect 236454 152640 236460 152652
rect 153712 152612 236460 152640
rect 153712 152600 153718 152612
rect 236454 152600 236460 152612
rect 236512 152600 236518 152652
rect 247034 152600 247040 152652
rect 247092 152640 247098 152652
rect 307754 152640 307760 152652
rect 247092 152612 307760 152640
rect 247092 152600 247098 152612
rect 307754 152600 307760 152612
rect 307812 152600 307818 152652
rect 311618 152600 311624 152652
rect 311676 152640 311682 152652
rect 320726 152640 320732 152652
rect 311676 152612 320732 152640
rect 311676 152600 311682 152612
rect 320726 152600 320732 152612
rect 320784 152600 320790 152652
rect 320818 152600 320824 152652
rect 320876 152640 320882 152652
rect 361666 152640 361672 152652
rect 320876 152612 361672 152640
rect 320876 152600 320882 152612
rect 361666 152600 361672 152612
rect 361724 152600 361730 152652
rect 364518 152600 364524 152652
rect 364576 152640 364582 152652
rect 396902 152640 396908 152652
rect 364576 152612 396908 152640
rect 364576 152600 364582 152612
rect 396902 152600 396908 152612
rect 396960 152600 396966 152652
rect 399110 152600 399116 152652
rect 399168 152640 399174 152652
rect 417418 152640 417424 152652
rect 399168 152612 417424 152640
rect 399168 152600 399174 152612
rect 417418 152600 417424 152612
rect 417476 152600 417482 152652
rect 418614 152600 418620 152652
rect 418672 152640 418678 152652
rect 427722 152640 427728 152652
rect 418672 152612 427728 152640
rect 418672 152600 418678 152612
rect 427722 152600 427728 152612
rect 427780 152600 427786 152652
rect 136876 152544 138014 152572
rect 136876 152532 136882 152544
rect 138290 152532 138296 152584
rect 138348 152572 138354 152584
rect 143994 152572 144000 152584
rect 138348 152544 144000 152572
rect 138348 152532 138354 152544
rect 143994 152532 144000 152544
rect 144052 152532 144058 152584
rect 144086 152532 144092 152584
rect 144144 152572 144150 152584
rect 226334 152572 226340 152584
rect 144144 152544 226340 152572
rect 144144 152532 144150 152544
rect 226334 152532 226340 152544
rect 226392 152532 226398 152584
rect 228818 152572 228824 152584
rect 226444 152544 228824 152572
rect 2866 152464 2872 152516
rect 2924 152504 2930 152516
rect 120810 152504 120816 152516
rect 2924 152476 120816 152504
rect 2924 152464 2930 152476
rect 120810 152464 120816 152476
rect 120868 152464 120874 152516
rect 126974 152464 126980 152516
rect 127032 152504 127038 152516
rect 215846 152504 215852 152516
rect 127032 152476 215852 152504
rect 127032 152464 127038 152476
rect 215846 152464 215852 152476
rect 215904 152464 215910 152516
rect 220722 152464 220728 152516
rect 220780 152504 220786 152516
rect 226444 152504 226472 152544
rect 228818 152532 228824 152544
rect 228876 152532 228882 152584
rect 234154 152532 234160 152584
rect 234212 152572 234218 152584
rect 297450 152572 297456 152584
rect 234212 152544 297456 152572
rect 234212 152532 234218 152544
rect 297450 152532 297456 152544
rect 297508 152532 297514 152584
rect 303614 152532 303620 152584
rect 303672 152572 303678 152584
rect 350718 152572 350724 152584
rect 303672 152544 350724 152572
rect 303672 152532 303678 152544
rect 350718 152532 350724 152544
rect 350776 152532 350782 152584
rect 351914 152532 351920 152584
rect 351972 152572 351978 152584
rect 353294 152572 353300 152584
rect 351972 152544 353300 152572
rect 351972 152532 351978 152544
rect 353294 152532 353300 152544
rect 353352 152532 353358 152584
rect 354490 152532 354496 152584
rect 354548 152572 354554 152584
rect 389266 152572 389272 152584
rect 354548 152544 389272 152572
rect 354548 152532 354554 152544
rect 389266 152532 389272 152544
rect 389324 152532 389330 152584
rect 393130 152532 393136 152584
rect 393188 152572 393194 152584
rect 418798 152572 418804 152584
rect 393188 152544 418804 152572
rect 393188 152532 393194 152544
rect 418798 152532 418804 152544
rect 418856 152532 418862 152584
rect 418890 152532 418896 152584
rect 418948 152572 418954 152584
rect 426894 152572 426900 152584
rect 418948 152544 426900 152572
rect 418948 152532 418954 152544
rect 426894 152532 426900 152544
rect 426952 152532 426958 152584
rect 220780 152476 226472 152504
rect 220780 152464 220786 152476
rect 227714 152464 227720 152516
rect 227772 152504 227778 152516
rect 292942 152504 292948 152516
rect 227772 152476 292948 152504
rect 227772 152464 227778 152476
rect 292942 152464 292948 152476
rect 293000 152464 293006 152516
rect 298646 152464 298652 152516
rect 298704 152504 298710 152516
rect 346854 152504 346860 152516
rect 298704 152476 346860 152504
rect 298704 152464 298710 152476
rect 346854 152464 346860 152476
rect 346912 152464 346918 152516
rect 348142 152464 348148 152516
rect 348200 152504 348206 152516
rect 385034 152504 385040 152516
rect 348200 152476 385040 152504
rect 348200 152464 348206 152476
rect 385034 152464 385040 152476
rect 385092 152464 385098 152516
rect 386414 152464 386420 152516
rect 386472 152504 386478 152516
rect 413646 152504 413652 152516
rect 386472 152476 413652 152504
rect 386472 152464 386478 152476
rect 413646 152464 413652 152476
rect 413704 152464 413710 152516
rect 415394 152464 415400 152516
rect 415452 152504 415458 152516
rect 430850 152504 430856 152516
rect 415452 152476 430856 152504
rect 415452 152464 415458 152476
rect 430850 152464 430856 152476
rect 430908 152464 430914 152516
rect 432570 152504 432598 152680
rect 432874 152668 432880 152720
rect 432932 152708 432938 152720
rect 438026 152708 438032 152720
rect 432932 152680 438032 152708
rect 432932 152668 432938 152680
rect 438026 152668 438032 152680
rect 438084 152668 438090 152720
rect 438118 152668 438124 152720
rect 438176 152708 438182 152720
rect 438176 152680 438992 152708
rect 438176 152668 438182 152680
rect 432690 152600 432696 152652
rect 432748 152640 432754 152652
rect 438762 152640 438768 152652
rect 432748 152612 438768 152640
rect 432748 152600 432754 152612
rect 438762 152600 438768 152612
rect 438820 152600 438826 152652
rect 432966 152532 432972 152584
rect 433024 152572 433030 152584
rect 438854 152572 438860 152584
rect 433024 152544 438860 152572
rect 433024 152532 433030 152544
rect 438854 152532 438860 152544
rect 438912 152532 438918 152584
rect 438964 152572 438992 152680
rect 440326 152668 440332 152720
rect 440384 152708 440390 152720
rect 455414 152708 455420 152720
rect 440384 152680 455420 152708
rect 440384 152668 440390 152680
rect 455414 152668 455420 152680
rect 455472 152668 455478 152720
rect 439038 152600 439044 152652
rect 439096 152640 439102 152652
rect 445754 152640 445760 152652
rect 439096 152612 445760 152640
rect 439096 152600 439102 152612
rect 445754 152600 445760 152612
rect 445812 152600 445818 152652
rect 440602 152572 440608 152584
rect 438964 152544 440608 152572
rect 440602 152532 440608 152544
rect 440660 152532 440666 152584
rect 442810 152532 442816 152584
rect 442868 152572 442874 152584
rect 456794 152572 456800 152584
rect 442868 152544 456800 152572
rect 442868 152532 442874 152544
rect 456794 152532 456800 152544
rect 456852 152532 456858 152584
rect 438118 152504 438124 152516
rect 432570 152476 438124 152504
rect 438118 152464 438124 152476
rect 438176 152464 438182 152516
rect 438578 152464 438584 152516
rect 438636 152504 438642 152516
rect 453482 152504 453488 152516
rect 438636 152476 453488 152504
rect 438636 152464 438642 152476
rect 453482 152464 453488 152476
rect 453540 152464 453546 152516
rect 66622 152396 66628 152448
rect 66680 152436 66686 152448
rect 159358 152436 159364 152448
rect 66680 152408 159364 152436
rect 66680 152396 66686 152408
rect 159358 152396 159364 152408
rect 159416 152396 159422 152448
rect 166994 152396 167000 152448
rect 167052 152436 167058 152448
rect 175918 152436 175924 152448
rect 167052 152408 175924 152436
rect 167052 152396 167058 152408
rect 175918 152396 175924 152408
rect 175976 152396 175982 152448
rect 176102 152396 176108 152448
rect 176160 152436 176166 152448
rect 249242 152436 249248 152448
rect 176160 152408 249248 152436
rect 176160 152396 176166 152408
rect 249242 152396 249248 152408
rect 249300 152396 249306 152448
rect 260834 152396 260840 152448
rect 260892 152436 260898 152448
rect 316034 152436 316040 152448
rect 260892 152408 316040 152436
rect 260892 152396 260898 152408
rect 316034 152396 316040 152408
rect 316092 152396 316098 152448
rect 317506 152396 317512 152448
rect 317564 152436 317570 152448
rect 320818 152436 320824 152448
rect 317564 152408 320824 152436
rect 317564 152396 317570 152408
rect 320818 152396 320824 152408
rect 320876 152396 320882 152448
rect 325878 152396 325884 152448
rect 325936 152436 325942 152448
rect 367370 152436 367376 152448
rect 325936 152408 367376 152436
rect 325936 152396 325942 152408
rect 367370 152396 367376 152408
rect 367428 152396 367434 152448
rect 371326 152396 371332 152448
rect 371384 152436 371390 152448
rect 402054 152436 402060 152448
rect 371384 152408 402060 152436
rect 371384 152396 371390 152408
rect 402054 152396 402060 152408
rect 402112 152396 402118 152448
rect 404170 152396 404176 152448
rect 404228 152436 404234 152448
rect 407942 152436 407948 152448
rect 404228 152408 407948 152436
rect 404228 152396 404234 152408
rect 407942 152396 407948 152408
rect 408000 152396 408006 152448
rect 410886 152396 410892 152448
rect 410944 152436 410950 152448
rect 430942 152436 430948 152448
rect 410944 152408 430948 152436
rect 410944 152396 410950 152408
rect 430942 152396 430948 152408
rect 431000 152396 431006 152448
rect 434714 152396 434720 152448
rect 434772 152436 434778 152448
rect 450906 152436 450912 152448
rect 434772 152408 450912 152436
rect 434772 152396 434778 152408
rect 450906 152396 450912 152408
rect 450964 152396 450970 152448
rect 33594 152328 33600 152380
rect 33652 152368 33658 152380
rect 109678 152368 109684 152380
rect 33652 152340 109684 152368
rect 33652 152328 33658 152340
rect 109678 152328 109684 152340
rect 109736 152328 109742 152380
rect 109770 152328 109776 152380
rect 109828 152368 109834 152380
rect 110506 152368 110512 152380
rect 109828 152340 110512 152368
rect 109828 152328 109834 152340
rect 110506 152328 110512 152340
rect 110564 152328 110570 152380
rect 120074 152328 120080 152380
rect 120132 152368 120138 152380
rect 210786 152368 210792 152380
rect 120132 152340 210792 152368
rect 120132 152328 120138 152340
rect 210786 152328 210792 152340
rect 210844 152328 210850 152380
rect 224034 152328 224040 152380
rect 224092 152368 224098 152380
rect 287790 152368 287796 152380
rect 224092 152340 287796 152368
rect 224092 152328 224098 152340
rect 287790 152328 287796 152340
rect 287848 152328 287854 152380
rect 292206 152328 292212 152380
rect 292264 152368 292270 152380
rect 341702 152368 341708 152380
rect 292264 152340 341708 152368
rect 292264 152328 292270 152340
rect 341702 152328 341708 152340
rect 341760 152328 341766 152380
rect 343818 152328 343824 152380
rect 343876 152368 343882 152380
rect 349798 152368 349804 152380
rect 343876 152340 349804 152368
rect 343876 152328 343882 152340
rect 349798 152328 349804 152340
rect 349856 152328 349862 152380
rect 349890 152328 349896 152380
rect 349948 152368 349954 152380
rect 385402 152368 385408 152380
rect 349948 152340 385408 152368
rect 349948 152328 349954 152340
rect 385402 152328 385408 152340
rect 385460 152328 385466 152380
rect 388346 152328 388352 152380
rect 388404 152368 388410 152380
rect 392026 152368 392032 152380
rect 388404 152340 392032 152368
rect 388404 152328 388410 152340
rect 392026 152328 392032 152340
rect 392084 152328 392090 152380
rect 394602 152328 394608 152380
rect 394660 152368 394666 152380
rect 417510 152368 417516 152380
rect 394660 152340 417516 152368
rect 394660 152328 394666 152340
rect 417510 152328 417516 152340
rect 417568 152328 417574 152380
rect 417602 152328 417608 152380
rect 417660 152368 417666 152380
rect 418890 152368 418896 152380
rect 417660 152340 418896 152368
rect 417660 152328 417666 152340
rect 418890 152328 418896 152340
rect 418948 152328 418954 152380
rect 426894 152328 426900 152380
rect 426952 152368 426958 152380
rect 431586 152368 431592 152380
rect 426952 152340 431592 152368
rect 426952 152328 426958 152340
rect 431586 152328 431592 152340
rect 431644 152328 431650 152380
rect 431862 152328 431868 152380
rect 431920 152368 431926 152380
rect 432506 152368 432512 152380
rect 431920 152340 432512 152368
rect 431920 152328 431926 152340
rect 432506 152328 432512 152340
rect 432564 152328 432570 152380
rect 432598 152328 432604 152380
rect 432656 152368 432662 152380
rect 441890 152368 441896 152380
rect 432656 152340 441896 152368
rect 432656 152328 432662 152340
rect 441890 152328 441896 152340
rect 441948 152328 441954 152380
rect 445294 152328 445300 152380
rect 445352 152368 445358 152380
rect 458542 152368 458548 152380
rect 445352 152340 458548 152368
rect 445352 152328 445358 152340
rect 458542 152328 458548 152340
rect 458600 152328 458606 152380
rect 9490 152260 9496 152312
rect 9548 152300 9554 152312
rect 82814 152300 82820 152312
rect 9548 152272 82820 152300
rect 9548 152260 9554 152272
rect 82814 152260 82820 152272
rect 82872 152260 82878 152312
rect 91094 152260 91100 152312
rect 91152 152300 91158 152312
rect 179966 152300 179972 152312
rect 91152 152272 179972 152300
rect 91152 152260 91158 152272
rect 179966 152260 179972 152272
rect 180024 152260 180030 152312
rect 187878 152260 187884 152312
rect 187936 152300 187942 152312
rect 262214 152300 262220 152312
rect 187936 152272 262220 152300
rect 187936 152260 187942 152272
rect 262214 152260 262220 152272
rect 262272 152260 262278 152312
rect 266354 152260 266360 152312
rect 266412 152300 266418 152312
rect 320542 152300 320548 152312
rect 266412 152272 320548 152300
rect 266412 152260 266418 152272
rect 320542 152260 320548 152272
rect 320600 152260 320606 152312
rect 320818 152260 320824 152312
rect 320876 152300 320882 152312
rect 325694 152300 325700 152312
rect 320876 152272 325700 152300
rect 320876 152260 320882 152272
rect 325694 152260 325700 152272
rect 325752 152260 325758 152312
rect 331214 152260 331220 152312
rect 331272 152300 331278 152312
rect 371878 152300 371884 152312
rect 331272 152272 371884 152300
rect 331272 152260 331278 152272
rect 371878 152260 371884 152272
rect 371936 152260 371942 152312
rect 381078 152260 381084 152312
rect 381136 152300 381142 152312
rect 409874 152300 409880 152312
rect 381136 152272 409880 152300
rect 381136 152260 381142 152272
rect 409874 152260 409880 152272
rect 409932 152260 409938 152312
rect 412606 152272 412864 152300
rect 19794 152192 19800 152244
rect 19852 152232 19858 152244
rect 97902 152232 97908 152244
rect 19852 152204 97908 152232
rect 19852 152192 19858 152204
rect 97902 152192 97908 152204
rect 97960 152192 97966 152244
rect 109034 152192 109040 152244
rect 109092 152232 109098 152244
rect 130562 152232 130568 152244
rect 109092 152204 130568 152232
rect 109092 152192 109098 152204
rect 130562 152192 130568 152204
rect 130620 152192 130626 152244
rect 134058 152192 134064 152244
rect 134116 152232 134122 152244
rect 220998 152232 221004 152244
rect 134116 152204 221004 152232
rect 134116 152192 134122 152204
rect 220998 152192 221004 152204
rect 221056 152192 221062 152244
rect 222102 152192 222108 152244
rect 222160 152232 222166 152244
rect 282914 152232 282920 152244
rect 222160 152204 282920 152232
rect 222160 152192 222166 152204
rect 282914 152192 282920 152204
rect 282972 152192 282978 152244
rect 285766 152192 285772 152244
rect 285824 152232 285830 152244
rect 335906 152232 335912 152244
rect 285824 152204 335912 152232
rect 285824 152192 285830 152204
rect 335906 152192 335912 152204
rect 335964 152192 335970 152244
rect 349154 152192 349160 152244
rect 349212 152232 349218 152244
rect 349890 152232 349896 152244
rect 349212 152204 349896 152232
rect 349212 152192 349218 152204
rect 349890 152192 349896 152204
rect 349948 152192 349954 152244
rect 352006 152192 352012 152244
rect 352064 152232 352070 152244
rect 387978 152232 387984 152244
rect 352064 152204 387984 152232
rect 352064 152192 352070 152204
rect 387978 152192 387984 152204
rect 388036 152192 388042 152244
rect 388438 152192 388444 152244
rect 388496 152232 388502 152244
rect 407206 152232 407212 152244
rect 388496 152204 407212 152232
rect 388496 152192 388502 152204
rect 407206 152192 407212 152204
rect 407264 152192 407270 152244
rect 409230 152192 409236 152244
rect 409288 152232 409294 152244
rect 412606 152232 412634 152272
rect 409288 152204 412634 152232
rect 412836 152232 412864 152272
rect 412910 152260 412916 152312
rect 412968 152300 412974 152312
rect 420914 152300 420920 152312
rect 412968 152272 420920 152300
rect 412968 152260 412974 152272
rect 420914 152260 420920 152272
rect 420972 152260 420978 152312
rect 422294 152260 422300 152312
rect 422352 152300 422358 152312
rect 424042 152300 424048 152312
rect 422352 152272 424048 152300
rect 422352 152260 422358 152272
rect 424042 152260 424048 152272
rect 424100 152260 424106 152312
rect 425146 152260 425152 152312
rect 425204 152300 425210 152312
rect 432414 152300 432420 152312
rect 425204 152272 432420 152300
rect 425204 152260 425210 152272
rect 432414 152260 432420 152272
rect 432472 152260 432478 152312
rect 435542 152300 435548 152312
rect 432892 152272 435548 152300
rect 428366 152232 428372 152244
rect 412836 152204 428372 152232
rect 409288 152192 409294 152204
rect 428366 152192 428372 152204
rect 428424 152192 428430 152244
rect 432892 152232 432920 152272
rect 435542 152260 435548 152272
rect 435600 152260 435606 152312
rect 436094 152260 436100 152312
rect 436152 152300 436158 152312
rect 446490 152300 446496 152312
rect 436152 152272 446496 152300
rect 436152 152260 436158 152272
rect 446490 152260 446496 152272
rect 446548 152260 446554 152312
rect 457346 152300 457352 152312
rect 447796 152272 457352 152300
rect 428476 152204 432920 152232
rect 82906 152124 82912 152176
rect 82964 152164 82970 152176
rect 169754 152164 169760 152176
rect 82964 152136 169760 152164
rect 82964 152124 82970 152136
rect 169754 152124 169760 152136
rect 169812 152124 169818 152176
rect 172698 152124 172704 152176
rect 172756 152164 172762 152176
rect 176102 152164 176108 152176
rect 172756 152136 176108 152164
rect 172756 152124 172762 152136
rect 176102 152124 176108 152136
rect 176160 152124 176166 152176
rect 176194 152124 176200 152176
rect 176252 152164 176258 152176
rect 190178 152164 190184 152176
rect 176252 152136 190184 152164
rect 176252 152124 176258 152136
rect 190178 152124 190184 152136
rect 190236 152124 190242 152176
rect 193398 152124 193404 152176
rect 193456 152164 193462 152176
rect 213270 152164 213276 152176
rect 193456 152136 213276 152164
rect 193456 152124 193462 152136
rect 213270 152124 213276 152136
rect 213328 152124 213334 152176
rect 244366 152124 244372 152176
rect 244424 152164 244430 152176
rect 305730 152164 305736 152176
rect 244424 152136 305736 152164
rect 244424 152124 244430 152136
rect 305730 152124 305736 152136
rect 305788 152124 305794 152176
rect 320726 152124 320732 152176
rect 320784 152164 320790 152176
rect 356514 152164 356520 152176
rect 320784 152136 356520 152164
rect 320784 152124 320790 152136
rect 356514 152124 356520 152136
rect 356572 152124 356578 152176
rect 357526 152124 357532 152176
rect 357584 152164 357590 152176
rect 359090 152164 359096 152176
rect 357584 152136 359096 152164
rect 357584 152124 357590 152136
rect 359090 152124 359096 152136
rect 359148 152124 359154 152176
rect 365714 152124 365720 152176
rect 365772 152164 365778 152176
rect 398190 152164 398196 152176
rect 365772 152136 398196 152164
rect 365772 152124 365778 152136
rect 398190 152124 398196 152136
rect 398248 152124 398254 152176
rect 405458 152124 405464 152176
rect 405516 152164 405522 152176
rect 412726 152164 412732 152176
rect 405516 152136 412732 152164
rect 405516 152124 405522 152136
rect 412726 152124 412732 152136
rect 412784 152124 412790 152176
rect 413002 152164 413008 152176
rect 412836 152136 413008 152164
rect 78766 152056 78772 152108
rect 78824 152096 78830 152108
rect 164510 152096 164516 152108
rect 78824 152068 164516 152096
rect 78824 152056 78830 152068
rect 164510 152056 164516 152068
rect 164568 152056 164574 152108
rect 169846 152056 169852 152108
rect 169904 152096 169910 152108
rect 169904 152068 175872 152096
rect 169904 152056 169910 152068
rect 68922 151988 68928 152040
rect 68980 152028 68986 152040
rect 142798 152028 142804 152040
rect 68980 152000 142804 152028
rect 68980 151988 68986 152000
rect 142798 151988 142804 152000
rect 142856 151988 142862 152040
rect 143350 151988 143356 152040
rect 143408 152028 143414 152040
rect 146662 152028 146668 152040
rect 143408 152000 146668 152028
rect 143408 151988 143414 152000
rect 146662 151988 146668 152000
rect 146720 151988 146726 152040
rect 156414 151988 156420 152040
rect 156472 152028 156478 152040
rect 172514 152028 172520 152040
rect 156472 152000 172520 152028
rect 156472 151988 156478 152000
rect 172514 151988 172520 152000
rect 172572 151988 172578 152040
rect 175844 152028 175872 152068
rect 175918 152056 175924 152108
rect 175976 152096 175982 152108
rect 182450 152096 182456 152108
rect 175976 152068 182456 152096
rect 175976 152056 175982 152068
rect 182450 152056 182456 152068
rect 182508 152056 182514 152108
rect 182542 152056 182548 152108
rect 182600 152096 182606 152108
rect 182600 152068 186314 152096
rect 182600 152056 182606 152068
rect 185026 152028 185032 152040
rect 175844 152000 185032 152028
rect 185026 151988 185032 152000
rect 185084 151988 185090 152040
rect 186286 152028 186314 152068
rect 191650 152056 191656 152108
rect 191708 152096 191714 152108
rect 208394 152096 208400 152108
rect 191708 152068 208400 152096
rect 191708 152056 191714 152068
rect 208394 152056 208400 152068
rect 208452 152056 208458 152108
rect 213638 152056 213644 152108
rect 213696 152096 213702 152108
rect 274266 152096 274272 152108
rect 213696 152068 274272 152096
rect 213696 152056 213702 152068
rect 274266 152056 274272 152068
rect 274324 152056 274330 152108
rect 277394 152056 277400 152108
rect 277452 152096 277458 152108
rect 330846 152096 330852 152108
rect 277452 152068 330852 152096
rect 277452 152056 277458 152068
rect 330846 152056 330852 152068
rect 330904 152056 330910 152108
rect 335354 152056 335360 152108
rect 335412 152096 335418 152108
rect 375374 152096 375380 152108
rect 335412 152068 375380 152096
rect 335412 152056 335418 152068
rect 375374 152056 375380 152068
rect 375432 152056 375438 152108
rect 384942 152056 384948 152108
rect 385000 152096 385006 152108
rect 391934 152096 391940 152108
rect 385000 152068 391940 152096
rect 385000 152056 385006 152068
rect 391934 152056 391940 152068
rect 391992 152056 391998 152108
rect 392026 152056 392032 152108
rect 392084 152096 392090 152108
rect 404630 152096 404636 152108
rect 392084 152068 404636 152096
rect 392084 152056 392090 152068
rect 404630 152056 404636 152068
rect 404688 152056 404694 152108
rect 412836 152096 412864 152136
rect 413002 152124 413008 152136
rect 413060 152124 413066 152176
rect 413922 152124 413928 152176
rect 413980 152164 413986 152176
rect 416222 152164 416228 152176
rect 413980 152136 416228 152164
rect 413980 152124 413986 152136
rect 416222 152124 416228 152136
rect 416280 152124 416286 152176
rect 416590 152124 416596 152176
rect 416648 152164 416654 152176
rect 426526 152164 426532 152176
rect 416648 152136 426532 152164
rect 416648 152124 416654 152136
rect 426526 152124 426532 152136
rect 426584 152124 426590 152176
rect 426636 152136 427400 152164
rect 423306 152096 423312 152108
rect 407776 152068 412864 152096
rect 413664 152068 423312 152096
rect 200482 152028 200488 152040
rect 186286 152000 200488 152028
rect 200482 151988 200488 152000
rect 200540 151988 200546 152040
rect 212626 151988 212632 152040
rect 212684 152028 212690 152040
rect 272426 152028 272432 152040
rect 212684 152000 272432 152028
rect 212684 151988 212690 152000
rect 272426 151988 272432 152000
rect 272484 151988 272490 152040
rect 272518 151988 272524 152040
rect 272576 152028 272582 152040
rect 320818 152028 320824 152040
rect 272576 152000 320824 152028
rect 272576 151988 272582 152000
rect 320818 151988 320824 152000
rect 320876 151988 320882 152040
rect 321554 151988 321560 152040
rect 321612 152028 321618 152040
rect 362310 152028 362316 152040
rect 321612 152000 362316 152028
rect 321612 151988 321618 152000
rect 362310 151988 362316 152000
rect 362368 151988 362374 152040
rect 378594 151988 378600 152040
rect 378652 152028 378658 152040
rect 384114 152028 384120 152040
rect 378652 152000 384120 152028
rect 378652 151988 378658 152000
rect 384114 151988 384120 152000
rect 384172 151988 384178 152040
rect 386322 151988 386328 152040
rect 386380 152028 386386 152040
rect 399478 152028 399484 152040
rect 386380 152000 399484 152028
rect 386380 151988 386386 152000
rect 399478 151988 399484 152000
rect 399536 151988 399542 152040
rect 75086 151920 75092 151972
rect 75144 151960 75150 151972
rect 154206 151960 154212 151972
rect 75144 151932 154212 151960
rect 75144 151920 75150 151932
rect 154206 151920 154212 151932
rect 154264 151920 154270 151972
rect 162578 151920 162584 151972
rect 162636 151960 162642 151972
rect 177390 151960 177396 151972
rect 162636 151932 177396 151960
rect 162636 151920 162642 151932
rect 177390 151920 177396 151932
rect 177448 151920 177454 151972
rect 184658 151920 184664 151972
rect 184716 151960 184722 151972
rect 195330 151960 195336 151972
rect 184716 151932 195336 151960
rect 184716 151920 184722 151932
rect 195330 151920 195336 151932
rect 195388 151920 195394 151972
rect 241606 151920 241612 151972
rect 241664 151960 241670 151972
rect 300854 151960 300860 151972
rect 241664 151932 300860 151960
rect 241664 151920 241670 151932
rect 300854 151920 300860 151932
rect 300912 151920 300918 151972
rect 304074 151920 304080 151972
rect 304132 151960 304138 151972
rect 351362 151960 351368 151972
rect 304132 151932 351368 151960
rect 304132 151920 304138 151932
rect 351362 151920 351368 151932
rect 351420 151920 351426 151972
rect 354674 151920 354680 151972
rect 354732 151960 354738 151972
rect 389910 151960 389916 151972
rect 354732 151932 389916 151960
rect 354732 151920 354738 151932
rect 389910 151920 389916 151932
rect 389968 151920 389974 151972
rect 398926 151920 398932 151972
rect 398984 151960 398990 151972
rect 407776 151960 407804 152068
rect 413554 152028 413560 152040
rect 398984 151932 407804 151960
rect 407868 152000 413560 152028
rect 398984 151920 398990 151932
rect 30190 151852 30196 151904
rect 30248 151892 30254 151904
rect 110322 151892 110328 151904
rect 30248 151864 110328 151892
rect 30248 151852 30254 151864
rect 110322 151852 110328 151864
rect 110380 151852 110386 151904
rect 110506 151852 110512 151904
rect 110564 151892 110570 151904
rect 138290 151892 138296 151904
rect 110564 151864 138296 151892
rect 110564 151852 110570 151864
rect 138290 151852 138296 151864
rect 138348 151852 138354 151904
rect 139302 151852 139308 151904
rect 139360 151892 139366 151904
rect 203058 151892 203064 151904
rect 139360 151864 203064 151892
rect 139360 151852 139366 151864
rect 203058 151852 203064 151864
rect 203116 151852 203122 151904
rect 243354 151852 243360 151904
rect 243412 151892 243418 151904
rect 302602 151892 302608 151904
rect 243412 151864 302608 151892
rect 243412 151852 243418 151864
rect 302602 151852 302608 151864
rect 302660 151852 302666 151904
rect 307386 151852 307392 151904
rect 307444 151892 307450 151904
rect 352006 151892 352012 151904
rect 307444 151864 352012 151892
rect 307444 151852 307450 151864
rect 352006 151852 352012 151864
rect 352064 151852 352070 151904
rect 363230 151852 363236 151904
rect 363288 151892 363294 151904
rect 364334 151892 364340 151904
rect 363288 151864 364340 151892
rect 363288 151852 363294 151864
rect 364334 151852 364340 151864
rect 364392 151852 364398 151904
rect 385126 151852 385132 151904
rect 385184 151892 385190 151904
rect 394694 151892 394700 151904
rect 385184 151864 394700 151892
rect 385184 151852 385190 151864
rect 394694 151852 394700 151864
rect 394752 151852 394758 151904
rect 396258 151852 396264 151904
rect 396316 151892 396322 151904
rect 402974 151892 402980 151904
rect 396316 151864 402980 151892
rect 396316 151852 396322 151864
rect 402974 151852 402980 151864
rect 403032 151852 403038 151904
rect 404262 151852 404268 151904
rect 404320 151892 404326 151904
rect 407868 151892 407896 152000
rect 413554 151988 413560 152000
rect 413612 151988 413618 152040
rect 408586 151920 408592 151972
rect 408644 151960 408650 151972
rect 413664 151960 413692 152068
rect 423306 152056 423312 152068
rect 423364 152056 423370 152108
rect 425974 152056 425980 152108
rect 426032 152096 426038 152108
rect 426636 152096 426664 152136
rect 426032 152068 426664 152096
rect 426032 152056 426038 152068
rect 419718 151988 419724 152040
rect 419776 152028 419782 152040
rect 427078 152028 427084 152040
rect 419776 152000 427084 152028
rect 419776 151988 419782 152000
rect 427078 151988 427084 152000
rect 427136 151988 427142 152040
rect 427372 152028 427400 152136
rect 427998 152124 428004 152176
rect 428056 152164 428062 152176
rect 428476 152164 428504 152204
rect 433058 152192 433064 152244
rect 433116 152232 433122 152244
rect 436186 152232 436192 152244
rect 433116 152204 436192 152232
rect 433116 152192 433122 152204
rect 436186 152192 436192 152204
rect 436244 152192 436250 152244
rect 436278 152192 436284 152244
rect 436336 152232 436342 152244
rect 447686 152232 447692 152244
rect 436336 152204 447692 152232
rect 436336 152192 436342 152204
rect 447686 152192 447692 152204
rect 447744 152192 447750 152244
rect 428056 152136 428504 152164
rect 428056 152124 428062 152136
rect 429286 152124 429292 152176
rect 429344 152164 429350 152176
rect 429344 152136 432828 152164
rect 429344 152124 429350 152136
rect 427446 152056 427452 152108
rect 427504 152096 427510 152108
rect 432414 152096 432420 152108
rect 427504 152068 432420 152096
rect 427504 152056 427510 152068
rect 432414 152056 432420 152068
rect 432472 152056 432478 152108
rect 432800 152096 432828 152136
rect 432966 152124 432972 152176
rect 433024 152164 433030 152176
rect 443822 152164 443828 152176
rect 433024 152136 443828 152164
rect 433024 152124 433030 152136
rect 443822 152124 443828 152136
rect 443880 152124 443886 152176
rect 443914 152124 443920 152176
rect 443972 152164 443978 152176
rect 447796 152164 447824 152272
rect 457346 152260 457352 152272
rect 457404 152260 457410 152312
rect 443972 152136 447824 152164
rect 443972 152124 443978 152136
rect 447870 152124 447876 152176
rect 447928 152164 447934 152176
rect 456058 152164 456064 152176
rect 447928 152136 456064 152164
rect 447928 152124 447934 152136
rect 456058 152124 456064 152136
rect 456116 152124 456122 152176
rect 446306 152096 446312 152108
rect 432800 152068 446312 152096
rect 446306 152056 446312 152068
rect 446364 152056 446370 152108
rect 446398 152056 446404 152108
rect 446456 152096 446462 152108
rect 449894 152096 449900 152108
rect 446456 152068 449900 152096
rect 446456 152056 446462 152068
rect 449894 152056 449900 152068
rect 449952 152056 449958 152108
rect 515766 152056 515772 152108
rect 515824 152096 515830 152108
rect 518986 152096 518992 152108
rect 515824 152068 518992 152096
rect 515824 152056 515830 152068
rect 518986 152056 518992 152068
rect 519044 152056 519050 152108
rect 432322 152028 432328 152040
rect 427372 152000 432328 152028
rect 432322 151988 432328 152000
rect 432380 151988 432386 152040
rect 432874 151988 432880 152040
rect 432932 152028 432938 152040
rect 443178 152028 443184 152040
rect 432932 152000 443184 152028
rect 432932 151988 432938 152000
rect 443178 151988 443184 152000
rect 443236 151988 443242 152040
rect 444466 151988 444472 152040
rect 444524 152028 444530 152040
rect 458174 152028 458180 152040
rect 444524 152000 458180 152028
rect 444524 151988 444530 152000
rect 458174 151988 458180 152000
rect 458232 151988 458238 152040
rect 459554 151988 459560 152040
rect 459612 152028 459618 152040
rect 461762 152028 461768 152040
rect 459612 152000 461768 152028
rect 459612 151988 459618 152000
rect 461762 151988 461768 152000
rect 461820 151988 461826 152040
rect 485774 151988 485780 152040
rect 485832 152028 485838 152040
rect 490006 152028 490012 152040
rect 485832 152000 490012 152028
rect 485832 151988 485838 152000
rect 490006 151988 490012 152000
rect 490064 151988 490070 152040
rect 516042 151988 516048 152040
rect 516100 152028 516106 152040
rect 520182 152028 520188 152040
rect 516100 152000 520188 152028
rect 516100 151988 516106 152000
rect 520182 151988 520188 152000
rect 520240 151988 520246 152040
rect 408644 151932 413692 151960
rect 408644 151920 408650 151932
rect 413830 151920 413836 151972
rect 413888 151960 413894 151972
rect 421374 151960 421380 151972
rect 413888 151932 421380 151960
rect 413888 151920 413894 151932
rect 421374 151920 421380 151932
rect 421432 151920 421438 151972
rect 422754 151920 422760 151972
rect 422812 151960 422818 151972
rect 432598 151960 432604 151972
rect 422812 151932 432604 151960
rect 422812 151920 422818 151932
rect 432598 151920 432604 151932
rect 432656 151920 432662 151972
rect 432690 151920 432696 151972
rect 432748 151960 432754 151972
rect 435450 151960 435456 151972
rect 432748 151932 435456 151960
rect 432748 151920 432754 151932
rect 435450 151920 435456 151932
rect 435508 151920 435514 151972
rect 435542 151920 435548 151972
rect 435600 151960 435606 151972
rect 439314 151960 439320 151972
rect 435600 151932 439320 151960
rect 435600 151920 435606 151932
rect 439314 151920 439320 151932
rect 439372 151920 439378 151972
rect 440234 151920 440240 151972
rect 440292 151960 440298 151972
rect 454770 151960 454776 151972
rect 440292 151932 454776 151960
rect 440292 151920 440298 151932
rect 454770 151920 454776 151932
rect 454828 151920 454834 151972
rect 469214 151920 469220 151972
rect 469272 151960 469278 151972
rect 472066 151960 472072 151972
rect 469272 151932 472072 151960
rect 469272 151920 469278 151932
rect 472066 151920 472072 151932
rect 472124 151920 472130 151972
rect 487338 151920 487344 151972
rect 487396 151960 487402 151972
rect 490650 151960 490656 151972
rect 487396 151932 490656 151960
rect 487396 151920 487402 151932
rect 490650 151920 490656 151932
rect 490708 151920 490714 151972
rect 509142 151920 509148 151972
rect 509200 151960 509206 151972
rect 510890 151960 510896 151972
rect 509200 151932 510896 151960
rect 509200 151920 509206 151932
rect 510890 151920 510896 151932
rect 510948 151920 510954 151972
rect 517422 151920 517428 151972
rect 517480 151960 517486 151972
rect 521562 151960 521568 151972
rect 517480 151932 521568 151960
rect 517480 151920 517486 151932
rect 521562 151920 521568 151932
rect 521620 151920 521626 151972
rect 404320 151864 407896 151892
rect 404320 151852 404326 151864
rect 407942 151852 407948 151904
rect 408000 151892 408006 151904
rect 415670 151892 415676 151904
rect 408000 151864 415676 151892
rect 408000 151852 408006 151864
rect 415670 151852 415676 151864
rect 415728 151852 415734 151904
rect 418154 151892 418160 151904
rect 415780 151864 418160 151892
rect 74810 151784 74816 151836
rect 74868 151824 74874 151836
rect 81342 151824 81348 151836
rect 74868 151796 81348 151824
rect 74868 151784 74874 151796
rect 81342 151784 81348 151796
rect 81400 151784 81406 151836
rect 105814 151784 105820 151836
rect 105872 151824 105878 151836
rect 110230 151824 110236 151836
rect 105872 151796 110236 151824
rect 105872 151784 105878 151796
rect 110230 151784 110236 151796
rect 110288 151784 110294 151836
rect 110414 151784 110420 151836
rect 110472 151824 110478 151836
rect 127894 151824 127900 151836
rect 110472 151796 127900 151824
rect 110472 151784 110478 151796
rect 127894 151784 127900 151796
rect 127952 151784 127958 151836
rect 129734 151784 129740 151836
rect 129792 151824 129798 151836
rect 146570 151824 146576 151836
rect 129792 151796 146576 151824
rect 129792 151784 129798 151796
rect 146570 151784 146576 151796
rect 146628 151784 146634 151836
rect 146662 151784 146668 151836
rect 146720 151824 146726 151836
rect 156782 151824 156788 151836
rect 146720 151796 156788 151824
rect 146720 151784 146726 151796
rect 156782 151784 156788 151796
rect 156840 151784 156846 151836
rect 172422 151784 172428 151836
rect 172480 151824 172486 151836
rect 176194 151824 176200 151836
rect 172480 151796 176200 151824
rect 172480 151784 172486 151796
rect 176194 151784 176200 151796
rect 176252 151784 176258 151836
rect 283190 151784 283196 151836
rect 283248 151824 283254 151836
rect 287146 151824 287152 151836
rect 283248 151796 287152 151824
rect 283248 151784 283254 151796
rect 287146 151784 287152 151796
rect 287204 151784 287210 151836
rect 299658 151784 299664 151836
rect 299716 151824 299722 151836
rect 346394 151824 346400 151836
rect 299716 151796 342944 151824
rect 299716 151784 299722 151796
rect 81710 151716 81716 151768
rect 81768 151756 81774 151768
rect 112806 151756 112812 151768
rect 81768 151728 112812 151756
rect 81768 151716 81774 151728
rect 112806 151716 112812 151728
rect 112864 151716 112870 151768
rect 342916 151756 342944 151796
rect 343744 151796 345060 151824
rect 343744 151756 343772 151796
rect 342916 151728 343772 151756
rect 345032 151756 345060 151796
rect 345676 151796 346400 151824
rect 345676 151756 345704 151796
rect 346394 151784 346400 151796
rect 346452 151784 346458 151836
rect 349798 151784 349804 151836
rect 349856 151824 349862 151836
rect 380250 151824 380256 151836
rect 349856 151796 380256 151824
rect 349856 151784 349862 151796
rect 380250 151784 380256 151796
rect 380308 151784 380314 151836
rect 398098 151784 398104 151836
rect 398156 151824 398162 151836
rect 407850 151824 407856 151836
rect 398156 151796 407856 151824
rect 398156 151784 398162 151796
rect 407850 151784 407856 151796
rect 407908 151784 407914 151836
rect 413554 151784 413560 151836
rect 413612 151824 413618 151836
rect 415780 151824 415808 151864
rect 418154 151852 418160 151864
rect 418212 151852 418218 151904
rect 419626 151852 419632 151904
rect 419684 151892 419690 151904
rect 436738 151892 436744 151904
rect 419684 151864 436744 151892
rect 419684 151852 419690 151864
rect 436738 151852 436744 151864
rect 436796 151852 436802 151904
rect 441246 151892 441252 151904
rect 437446 151864 441252 151892
rect 413612 151796 415808 151824
rect 413612 151784 413618 151796
rect 417418 151784 417424 151836
rect 417476 151824 417482 151836
rect 423950 151824 423956 151836
rect 417476 151796 423956 151824
rect 417476 151784 417482 151796
rect 423950 151784 423956 151796
rect 424008 151784 424014 151836
rect 424042 151784 424048 151836
rect 424100 151824 424106 151836
rect 437446 151824 437474 151864
rect 441246 151852 441252 151864
rect 441304 151852 441310 151904
rect 441798 151852 441804 151904
rect 441856 151892 441862 151904
rect 446214 151892 446220 151904
rect 441856 151864 446220 151892
rect 441856 151852 441862 151864
rect 446214 151852 446220 151864
rect 446272 151852 446278 151904
rect 446490 151852 446496 151904
rect 446548 151892 446554 151904
rect 451550 151892 451556 151904
rect 446548 151864 451556 151892
rect 446548 151852 446554 151864
rect 451550 151852 451556 151864
rect 451608 151852 451614 151904
rect 468018 151852 468024 151904
rect 468076 151892 468082 151904
rect 470778 151892 470784 151904
rect 468076 151864 470784 151892
rect 468076 151852 468082 151864
rect 470778 151852 470784 151864
rect 470836 151852 470842 151904
rect 488166 151852 488172 151904
rect 488224 151852 488230 151904
rect 488534 151852 488540 151904
rect 488592 151892 488598 151904
rect 491938 151892 491944 151904
rect 488592 151864 491944 151892
rect 488592 151852 488598 151864
rect 491938 151852 491944 151864
rect 491996 151852 492002 151904
rect 507762 151852 507768 151904
rect 507820 151892 507826 151904
rect 509510 151892 509516 151904
rect 507820 151864 509516 151892
rect 507820 151852 507826 151864
rect 509510 151852 509516 151864
rect 509568 151852 509574 151904
rect 424100 151796 437474 151824
rect 424100 151784 424106 151796
rect 437750 151784 437756 151836
rect 437808 151824 437814 151836
rect 452838 151824 452844 151836
rect 437808 151796 440188 151824
rect 437808 151784 437814 151796
rect 345032 151728 345704 151756
rect 432414 151716 432420 151768
rect 432472 151756 432478 151768
rect 434162 151756 434168 151768
rect 432472 151728 434168 151756
rect 432472 151716 432478 151728
rect 434162 151716 434168 151728
rect 434220 151716 434226 151768
rect 440160 151756 440188 151796
rect 440712 151796 452844 151824
rect 440712 151756 440740 151796
rect 452838 151784 452844 151796
rect 452896 151784 452902 151836
rect 467926 151784 467932 151836
rect 467984 151824 467990 151836
rect 471422 151824 471428 151836
rect 467984 151796 471428 151824
rect 467984 151784 467990 151796
rect 471422 151784 471428 151796
rect 471480 151784 471486 151836
rect 488184 151824 488212 151852
rect 491294 151824 491300 151836
rect 488184 151796 491300 151824
rect 491294 151784 491300 151796
rect 491352 151784 491358 151836
rect 499114 151784 499120 151836
rect 499172 151824 499178 151836
rect 499758 151824 499764 151836
rect 499172 151796 499764 151824
rect 499172 151784 499178 151796
rect 499758 151784 499764 151796
rect 499816 151784 499822 151836
rect 517054 151784 517060 151836
rect 517112 151824 517118 151836
rect 520274 151824 520280 151836
rect 517112 151796 520280 151824
rect 517112 151784 517118 151796
rect 520274 151784 520280 151796
rect 520332 151784 520338 151836
rect 440160 151728 440740 151756
rect 98914 151648 98920 151700
rect 98972 151688 98978 151700
rect 116026 151688 116032 151700
rect 98972 151660 116032 151688
rect 98972 151648 98978 151660
rect 116026 151648 116032 151660
rect 116084 151648 116090 151700
rect 95510 151580 95516 151632
rect 95568 151620 95574 151632
rect 115290 151620 115296 151632
rect 95568 151592 115296 151620
rect 95568 151580 95574 151592
rect 115290 151580 115296 151592
rect 115348 151580 115354 151632
rect 92014 151512 92020 151564
rect 92072 151552 92078 151564
rect 113082 151552 113088 151564
rect 92072 151524 113088 151552
rect 92072 151512 92078 151524
rect 113082 151512 113088 151524
rect 113140 151512 113146 151564
rect 26694 151444 26700 151496
rect 26752 151484 26758 151496
rect 116946 151484 116952 151496
rect 26752 151456 116952 151484
rect 26752 151444 26758 151456
rect 116946 151444 116952 151456
rect 117004 151444 117010 151496
rect 16390 151376 16396 151428
rect 16448 151416 16454 151428
rect 116762 151416 116768 151428
rect 16448 151388 116768 151416
rect 16448 151376 16454 151388
rect 116762 151376 116768 151388
rect 116820 151376 116826 151428
rect 12986 151308 12992 151360
rect 13044 151348 13050 151360
rect 116670 151348 116676 151360
rect 13044 151320 116676 151348
rect 13044 151308 13050 151320
rect 116670 151308 116676 151320
rect 116728 151308 116734 151360
rect 68002 151240 68008 151292
rect 68060 151280 68066 151292
rect 112714 151280 112720 151292
rect 68060 151252 112720 151280
rect 68060 151240 68066 151252
rect 112714 151240 112720 151252
rect 112772 151240 112778 151292
rect 64506 151172 64512 151224
rect 64564 151212 64570 151224
rect 112622 151212 112628 151224
rect 64564 151184 112628 151212
rect 64564 151172 64570 151184
rect 112622 151172 112628 151184
rect 112680 151172 112686 151224
rect 61102 151104 61108 151156
rect 61160 151144 61166 151156
rect 112530 151144 112536 151156
rect 61160 151116 112536 151144
rect 61160 151104 61166 151116
rect 112530 151104 112536 151116
rect 112588 151104 112594 151156
rect 57698 151036 57704 151088
rect 57756 151076 57762 151088
rect 110966 151076 110972 151088
rect 57756 151048 110972 151076
rect 57756 151036 57762 151048
rect 110966 151036 110972 151048
rect 111024 151036 111030 151088
rect 54202 150968 54208 151020
rect 54260 151008 54266 151020
rect 112438 151008 112444 151020
rect 54260 150980 112444 151008
rect 54260 150968 54266 150980
rect 112438 150968 112444 150980
rect 112496 150968 112502 151020
rect 50798 150900 50804 150952
rect 50856 150940 50862 150952
rect 111702 150940 111708 150952
rect 50856 150912 111708 150940
rect 50856 150900 50862 150912
rect 111702 150900 111708 150912
rect 111760 150900 111766 150952
rect 47302 150832 47308 150884
rect 47360 150872 47366 150884
rect 111610 150872 111616 150884
rect 47360 150844 111616 150872
rect 47360 150832 47366 150844
rect 111610 150832 111616 150844
rect 111668 150832 111674 150884
rect 43898 150764 43904 150816
rect 43956 150804 43962 150816
rect 111518 150804 111524 150816
rect 43956 150776 111524 150804
rect 43956 150764 43962 150776
rect 111518 150764 111524 150776
rect 111576 150764 111582 150816
rect 40494 150696 40500 150748
rect 40552 150736 40558 150748
rect 111426 150736 111432 150748
rect 40552 150708 111432 150736
rect 40552 150696 40558 150708
rect 111426 150696 111432 150708
rect 111484 150696 111490 150748
rect 36998 150628 37004 150680
rect 37056 150668 37062 150680
rect 111242 150668 111248 150680
rect 37056 150640 111248 150668
rect 37056 150628 37062 150640
rect 111242 150628 111248 150640
rect 111300 150628 111306 150680
rect 88610 150560 88616 150612
rect 88668 150600 88674 150612
rect 112990 150600 112996 150612
rect 88668 150572 112996 150600
rect 88668 150560 88674 150572
rect 112990 150560 112996 150572
rect 113048 150560 113054 150612
rect 85206 150492 85212 150544
rect 85264 150532 85270 150544
rect 115198 150532 115204 150544
rect 85264 150504 115204 150532
rect 85264 150492 85270 150504
rect 115198 150492 115204 150504
rect 115256 150492 115262 150544
rect 122834 150492 122840 150544
rect 122892 150532 122898 150544
rect 123386 150532 123392 150544
rect 122892 150504 123392 150532
rect 122892 150492 122898 150504
rect 123386 150492 123392 150504
rect 123444 150492 123450 150544
rect 283098 150492 283104 150544
rect 283156 150532 283162 150544
rect 283926 150532 283932 150544
rect 283156 150504 283932 150532
rect 283156 150492 283162 150504
rect 283926 150492 283932 150504
rect 283984 150492 283990 150544
rect 299474 150492 299480 150544
rect 299532 150532 299538 150544
rect 300026 150532 300032 150544
rect 299532 150504 300032 150532
rect 299532 150492 299538 150504
rect 300026 150492 300032 150504
rect 300084 150492 300090 150544
rect 328454 150492 328460 150544
rect 328512 150532 328518 150544
rect 328914 150532 328920 150544
rect 328512 150504 328920 150532
rect 328512 150492 328518 150504
rect 328914 150492 328920 150504
rect 328972 150492 328978 150544
rect 332686 150492 332692 150544
rect 332744 150532 332750 150544
rect 333422 150532 333428 150544
rect 332744 150504 333428 150532
rect 332744 150492 332750 150504
rect 333422 150492 333428 150504
rect 333480 150492 333486 150544
rect 362954 150492 362960 150544
rect 363012 150532 363018 150544
rect 363598 150532 363604 150544
rect 363012 150504 363604 150532
rect 363012 150492 363018 150504
rect 363598 150492 363604 150504
rect 363656 150492 363662 150544
rect 102318 150424 102324 150476
rect 102376 150464 102382 150476
rect 116118 150464 116124 150476
rect 102376 150436 116124 150464
rect 102376 150424 102382 150436
rect 116118 150424 116124 150436
rect 116176 150424 116182 150476
rect 78306 150288 78312 150340
rect 78364 150328 78370 150340
rect 112898 150328 112904 150340
rect 78364 150300 112904 150328
rect 78364 150288 78370 150300
rect 112898 150288 112904 150300
rect 112956 150288 112962 150340
rect 110322 150220 110328 150272
rect 110380 150260 110386 150272
rect 117130 150260 117136 150272
rect 110380 150232 117136 150260
rect 110380 150220 110386 150232
rect 117130 150220 117136 150232
rect 117188 150220 117194 150272
rect 97902 150152 97908 150204
rect 97960 150192 97966 150204
rect 116854 150192 116860 150204
rect 97960 150164 116860 150192
rect 97960 150152 97966 150164
rect 116854 150152 116860 150164
rect 116912 150152 116918 150204
rect 81342 150084 81348 150136
rect 81400 150124 81406 150136
rect 81400 150096 84194 150124
rect 81400 150084 81406 150096
rect 84166 150056 84194 150096
rect 92474 150084 92480 150136
rect 92532 150124 92538 150136
rect 117222 150124 117228 150136
rect 92532 150096 117228 150124
rect 92532 150084 92538 150096
rect 117222 150084 117228 150096
rect 117280 150084 117286 150136
rect 116486 150056 116492 150068
rect 84166 150028 116492 150056
rect 116486 150016 116492 150028
rect 116544 150016 116550 150068
rect 111150 148316 111156 148368
rect 111208 148356 111214 148368
rect 117038 148356 117044 148368
rect 111208 148328 117044 148356
rect 111208 148316 111214 148328
rect 117038 148316 117044 148328
rect 117096 148316 117102 148368
rect 113082 140700 113088 140752
rect 113140 140740 113146 140752
rect 116118 140740 116124 140752
rect 113140 140712 116124 140740
rect 113140 140700 113146 140712
rect 116118 140700 116124 140712
rect 116176 140700 116182 140752
rect 112990 137912 112996 137964
rect 113048 137952 113054 137964
rect 116118 137952 116124 137964
rect 113048 137924 116124 137952
rect 113048 137912 113054 137924
rect 116118 137912 116124 137924
rect 116176 137912 116182 137964
rect 112806 133832 112812 133884
rect 112864 133872 112870 133884
rect 116026 133872 116032 133884
rect 112864 133844 116032 133872
rect 112864 133832 112870 133844
rect 116026 133832 116032 133844
rect 116084 133832 116090 133884
rect 114186 132608 114192 132660
rect 114244 132648 114250 132660
rect 115198 132648 115204 132660
rect 114244 132620 115204 132648
rect 114244 132608 114250 132620
rect 115198 132608 115204 132620
rect 115256 132608 115262 132660
rect 112898 132404 112904 132456
rect 112956 132444 112962 132456
rect 116118 132444 116124 132456
rect 112956 132416 116124 132444
rect 112956 132404 112962 132416
rect 116118 132404 116124 132416
rect 116176 132404 116182 132456
rect 112714 126896 112720 126948
rect 112772 126936 112778 126948
rect 116118 126936 116124 126948
rect 112772 126908 116124 126936
rect 112772 126896 112778 126908
rect 116118 126896 116124 126908
rect 116176 126896 116182 126948
rect 112622 124108 112628 124160
rect 112680 124148 112686 124160
rect 116118 124148 116124 124160
rect 112680 124120 116124 124148
rect 112680 124108 112686 124120
rect 116118 124108 116124 124120
rect 116176 124108 116182 124160
rect 112530 122748 112536 122800
rect 112588 122788 112594 122800
rect 115934 122788 115940 122800
rect 112588 122760 115940 122788
rect 112588 122748 112594 122760
rect 115934 122748 115940 122760
rect 115992 122748 115998 122800
rect 111702 121388 111708 121440
rect 111760 121428 111766 121440
rect 116118 121428 116124 121440
rect 111760 121400 116124 121428
rect 111760 121388 111766 121400
rect 116118 121388 116124 121400
rect 116176 121388 116182 121440
rect 112438 118600 112444 118652
rect 112496 118640 112502 118652
rect 116118 118640 116124 118652
rect 112496 118612 116124 118640
rect 112496 118600 112502 118612
rect 116118 118600 116124 118612
rect 116176 118600 116182 118652
rect 111610 117240 111616 117292
rect 111668 117280 111674 117292
rect 116118 117280 116124 117292
rect 111668 117252 116124 117280
rect 111668 117240 111674 117252
rect 116118 117240 116124 117252
rect 116176 117240 116182 117292
rect 111518 114452 111524 114504
rect 111576 114492 111582 114504
rect 116118 114492 116124 114504
rect 111576 114464 116124 114492
rect 111576 114452 111582 114464
rect 116118 114452 116124 114464
rect 116176 114452 116182 114504
rect 111426 113092 111432 113144
rect 111484 113132 111490 113144
rect 115934 113132 115940 113144
rect 111484 113104 115940 113132
rect 111484 113092 111490 113104
rect 115934 113092 115940 113104
rect 115992 113092 115998 113144
rect 111334 111732 111340 111784
rect 111392 111772 111398 111784
rect 116118 111772 116124 111784
rect 111392 111744 116124 111772
rect 111392 111732 111398 111744
rect 116118 111732 116124 111744
rect 116176 111732 116182 111784
rect 111150 108944 111156 108996
rect 111208 108984 111214 108996
rect 116118 108984 116124 108996
rect 111208 108956 116124 108984
rect 111208 108944 111214 108956
rect 116118 108944 116124 108956
rect 116176 108944 116182 108996
rect 111242 92420 111248 92472
rect 111300 92460 111306 92472
rect 116118 92460 116124 92472
rect 111300 92432 116124 92460
rect 111300 92420 111306 92432
rect 116118 92420 116124 92432
rect 116176 92420 116182 92472
rect 111058 89632 111064 89684
rect 111116 89672 111122 89684
rect 116118 89672 116124 89684
rect 111116 89644 116124 89672
rect 111116 89632 111122 89644
rect 116118 89632 116124 89644
rect 116176 89632 116182 89684
rect 113818 88272 113824 88324
rect 113876 88312 113882 88324
rect 116026 88312 116032 88324
rect 113876 88284 116032 88312
rect 113876 88272 113882 88284
rect 116026 88272 116032 88284
rect 116084 88272 116090 88324
rect 113910 83920 113916 83972
rect 113968 83960 113974 83972
rect 116578 83960 116584 83972
rect 113968 83932 116584 83960
rect 113968 83920 113974 83932
rect 116578 83920 116584 83932
rect 116636 83920 116642 83972
rect 114002 82764 114008 82816
rect 114060 82804 114066 82816
rect 116210 82804 116216 82816
rect 114060 82776 116216 82804
rect 114060 82764 114066 82776
rect 116210 82764 116216 82776
rect 116268 82764 116274 82816
rect 114094 79976 114100 80028
rect 114152 80016 114158 80028
rect 115934 80016 115940 80028
rect 114152 79988 115940 80016
rect 114152 79976 114158 79988
rect 115934 79976 115940 79988
rect 115992 79976 115998 80028
rect 114186 78616 114192 78668
rect 114244 78656 114250 78668
rect 116118 78656 116124 78668
rect 114244 78628 116124 78656
rect 114244 78616 114250 78628
rect 116118 78616 116124 78628
rect 116176 78616 116182 78668
rect 114186 71748 114192 71800
rect 114244 71788 114250 71800
rect 116578 71788 116584 71800
rect 114244 71760 116584 71788
rect 114244 71748 114250 71760
rect 116578 71748 116584 71760
rect 116636 71748 116642 71800
rect 114094 69028 114100 69080
rect 114152 69068 114158 69080
rect 116302 69068 116308 69080
rect 114152 69040 116308 69068
rect 114152 69028 114158 69040
rect 116302 69028 116308 69040
rect 116360 69028 116366 69080
rect 114002 67600 114008 67652
rect 114060 67640 114066 67652
rect 116118 67640 116124 67652
rect 114060 67612 116124 67640
rect 114060 67600 114066 67612
rect 116118 67600 116124 67612
rect 116176 67600 116182 67652
rect 113910 66240 113916 66292
rect 113968 66280 113974 66292
rect 116578 66280 116584 66292
rect 113968 66252 116584 66280
rect 113968 66240 113974 66252
rect 116578 66240 116584 66252
rect 116636 66240 116642 66292
rect 113358 64676 113364 64728
rect 113416 64716 113422 64728
rect 116578 64716 116584 64728
rect 113416 64688 116584 64716
rect 113416 64676 113422 64688
rect 116578 64676 116584 64688
rect 116636 64676 116642 64728
rect 113818 63520 113824 63572
rect 113876 63560 113882 63572
rect 116210 63560 116216 63572
rect 113876 63532 116216 63560
rect 113876 63520 113882 63532
rect 116210 63520 116216 63532
rect 116268 63520 116274 63572
rect 112438 62092 112444 62144
rect 112496 62132 112502 62144
rect 116118 62132 116124 62144
rect 112496 62104 116124 62132
rect 112496 62092 112502 62104
rect 116118 62092 116124 62104
rect 116176 62092 116182 62144
rect 112530 42780 112536 42832
rect 112588 42820 112594 42832
rect 116118 42820 116124 42832
rect 112588 42792 116124 42820
rect 112588 42780 112594 42792
rect 116118 42780 116124 42792
rect 116176 42780 116182 42832
rect 116394 7624 116400 7676
rect 116452 7624 116458 7676
rect 116302 7420 116308 7472
rect 116360 7460 116366 7472
rect 116412 7460 116440 7624
rect 116360 7432 116440 7460
rect 116360 7420 116366 7432
rect 111058 2796 111064 2848
rect 111116 2836 111122 2848
rect 111116 2808 143672 2836
rect 111116 2796 111122 2808
rect 143644 2508 143672 2808
rect 425808 2808 443684 2836
rect 425808 2508 425836 2808
rect 443656 2508 443684 2808
rect 143626 2456 143632 2508
rect 143684 2456 143690 2508
rect 425790 2456 425796 2508
rect 425848 2456 425854 2508
rect 443638 2456 443644 2508
rect 443696 2456 443702 2508
rect 102612 1924 109816 1952
rect 102612 1896 102640 1924
rect 109788 1896 109816 1924
rect 42058 1844 42064 1896
rect 42116 1884 42122 1896
rect 44726 1884 44732 1896
rect 42116 1856 44732 1884
rect 42116 1844 42122 1856
rect 44726 1844 44732 1856
rect 44784 1844 44790 1896
rect 62390 1844 62396 1896
rect 62448 1884 62454 1896
rect 68278 1884 68284 1896
rect 62448 1856 68284 1884
rect 62448 1844 62454 1856
rect 68278 1844 68284 1856
rect 68336 1844 68342 1896
rect 91922 1844 91928 1896
rect 91980 1884 91986 1896
rect 99190 1884 99196 1896
rect 91980 1856 99196 1884
rect 91980 1844 91986 1856
rect 99190 1844 99196 1856
rect 99248 1844 99254 1896
rect 102594 1844 102600 1896
rect 102652 1844 102658 1896
rect 102686 1844 102692 1896
rect 102744 1884 102750 1896
rect 102744 1856 105860 1884
rect 102744 1844 102750 1856
rect 89346 1776 89352 1828
rect 89404 1816 89410 1828
rect 105832 1816 105860 1856
rect 105906 1844 105912 1896
rect 105964 1884 105970 1896
rect 109126 1884 109132 1896
rect 105964 1856 109132 1884
rect 105964 1844 105970 1856
rect 109126 1844 109132 1856
rect 109184 1844 109190 1896
rect 109678 1884 109684 1896
rect 109236 1856 109684 1884
rect 109236 1816 109264 1856
rect 109678 1844 109684 1856
rect 109736 1844 109742 1896
rect 109770 1844 109776 1896
rect 109828 1844 109834 1896
rect 109862 1844 109868 1896
rect 109920 1884 109926 1896
rect 109920 1856 118694 1884
rect 109920 1844 109926 1856
rect 89404 1788 104204 1816
rect 105832 1788 109264 1816
rect 89404 1776 89410 1788
rect 59354 1708 59360 1760
rect 59412 1748 59418 1760
rect 78766 1748 78772 1760
rect 59412 1720 78772 1748
rect 59412 1708 59418 1720
rect 78766 1708 78772 1720
rect 78824 1708 78830 1760
rect 86034 1708 86040 1760
rect 86092 1748 86098 1760
rect 104176 1748 104204 1788
rect 109310 1776 109316 1828
rect 109368 1816 109374 1828
rect 112438 1816 112444 1828
rect 109368 1788 112444 1816
rect 109368 1776 109374 1788
rect 112438 1776 112444 1788
rect 112496 1776 112502 1828
rect 109954 1748 109960 1760
rect 86092 1720 104112 1748
rect 104176 1720 109960 1748
rect 86092 1708 86098 1720
rect 82630 1640 82636 1692
rect 82688 1680 82694 1692
rect 103974 1680 103980 1692
rect 82688 1652 103980 1680
rect 82688 1640 82694 1652
rect 103974 1640 103980 1652
rect 104032 1640 104038 1692
rect 104084 1680 104112 1720
rect 109954 1708 109960 1720
rect 110012 1708 110018 1760
rect 110046 1708 110052 1760
rect 110104 1748 110110 1760
rect 116578 1748 116584 1760
rect 110104 1720 116584 1748
rect 110104 1708 110110 1720
rect 116578 1708 116584 1720
rect 116636 1708 116642 1760
rect 104084 1652 109172 1680
rect 69290 1572 69296 1624
rect 69348 1612 69354 1624
rect 103790 1612 103796 1624
rect 69348 1584 103796 1612
rect 69348 1572 69354 1584
rect 103790 1572 103796 1584
rect 103848 1572 103854 1624
rect 105906 1612 105912 1624
rect 103900 1584 105912 1612
rect 79318 1504 79324 1556
rect 79376 1544 79382 1556
rect 103900 1544 103928 1584
rect 105906 1572 105912 1584
rect 105964 1572 105970 1624
rect 105998 1572 106004 1624
rect 106056 1612 106062 1624
rect 109034 1612 109040 1624
rect 106056 1584 109040 1612
rect 106056 1572 106062 1584
rect 109034 1572 109040 1584
rect 109092 1572 109098 1624
rect 109144 1612 109172 1652
rect 109218 1640 109224 1692
rect 109276 1680 109282 1692
rect 110598 1680 110604 1692
rect 109276 1652 110604 1680
rect 109276 1640 109282 1652
rect 110598 1640 110604 1652
rect 110656 1640 110662 1692
rect 110138 1612 110144 1624
rect 109144 1584 110144 1612
rect 110138 1572 110144 1584
rect 110196 1572 110202 1624
rect 79376 1516 103928 1544
rect 79376 1504 79382 1516
rect 103974 1504 103980 1556
rect 104032 1544 104038 1556
rect 110230 1544 110236 1556
rect 104032 1516 110236 1544
rect 104032 1504 104038 1516
rect 110230 1504 110236 1516
rect 110288 1504 110294 1556
rect 46014 1436 46020 1488
rect 46072 1476 46078 1488
rect 64046 1476 64052 1488
rect 46072 1448 64052 1476
rect 46072 1436 46078 1448
rect 64046 1436 64052 1448
rect 64104 1436 64110 1488
rect 72694 1436 72700 1488
rect 72752 1476 72758 1488
rect 109586 1476 109592 1488
rect 72752 1448 109592 1476
rect 72752 1436 72758 1448
rect 109586 1436 109592 1448
rect 109644 1436 109650 1488
rect 118666 1476 118694 1856
rect 193582 1476 193588 1488
rect 118666 1448 193588 1476
rect 193582 1436 193588 1448
rect 193640 1436 193646 1488
rect 32674 1368 32680 1420
rect 32732 1408 32738 1420
rect 109126 1408 109132 1420
rect 32732 1380 109132 1408
rect 32732 1368 32738 1380
rect 109126 1368 109132 1380
rect 109184 1368 109190 1420
rect 109218 1368 109224 1420
rect 109276 1408 109282 1420
rect 110046 1408 110052 1420
rect 109276 1380 110052 1408
rect 109276 1368 109282 1380
rect 110046 1368 110052 1380
rect 110104 1368 110110 1420
rect 116394 1408 116400 1420
rect 110156 1380 116400 1408
rect 2682 1300 2688 1352
rect 2740 1340 2746 1352
rect 2740 1312 109356 1340
rect 2740 1300 2746 1312
rect 35986 1232 35992 1284
rect 36044 1272 36050 1284
rect 109328 1272 109356 1312
rect 109402 1300 109408 1352
rect 109460 1340 109466 1352
rect 110156 1340 110184 1380
rect 116394 1368 116400 1380
rect 116452 1368 116458 1420
rect 294782 1368 294788 1420
rect 294840 1408 294846 1420
rect 343634 1408 343640 1420
rect 294840 1380 343640 1408
rect 294840 1368 294846 1380
rect 343634 1368 343640 1380
rect 343692 1368 343698 1420
rect 491294 1368 491300 1420
rect 491352 1408 491358 1420
rect 493594 1408 493600 1420
rect 491352 1380 493600 1408
rect 491352 1368 491358 1380
rect 493594 1368 493600 1380
rect 493652 1368 493658 1420
rect 109460 1312 110184 1340
rect 109460 1300 109466 1312
rect 116302 1272 116308 1284
rect 36044 1244 109264 1272
rect 109328 1244 116308 1272
rect 36044 1232 36050 1244
rect 39298 1164 39304 1216
rect 39356 1204 39362 1216
rect 109034 1204 109040 1216
rect 39356 1176 109040 1204
rect 39356 1164 39362 1176
rect 109034 1164 109040 1176
rect 109092 1164 109098 1216
rect 109236 1204 109264 1244
rect 116302 1232 116308 1244
rect 116360 1232 116366 1284
rect 116486 1204 116492 1216
rect 109236 1176 116492 1204
rect 116486 1164 116492 1176
rect 116544 1164 116550 1216
rect 49326 1096 49332 1148
rect 49384 1136 49390 1148
rect 117038 1136 117044 1148
rect 49384 1108 117044 1136
rect 49384 1096 49390 1108
rect 117038 1096 117044 1108
rect 117096 1096 117102 1148
rect 52638 1028 52644 1080
rect 52696 1068 52702 1080
rect 52696 1040 109172 1068
rect 52696 1028 52702 1040
rect 65978 960 65984 1012
rect 66036 1000 66042 1012
rect 97258 1000 97264 1012
rect 66036 972 97264 1000
rect 66036 960 66042 972
rect 97258 960 97264 972
rect 97316 960 97322 1012
rect 109144 1000 109172 1040
rect 116854 1000 116860 1012
rect 102106 972 106274 1000
rect 109144 972 116860 1000
rect 76006 892 76012 944
rect 76064 932 76070 944
rect 102106 932 102134 972
rect 76064 904 102134 932
rect 106246 932 106274 972
rect 116854 960 116860 972
rect 116912 960 116918 1012
rect 112530 932 112536 944
rect 106246 904 112536 932
rect 76064 892 76070 904
rect 112530 892 112536 904
rect 112588 892 112594 944
rect 91554 824 91560 876
rect 91612 864 91618 876
rect 93854 864 93860 876
rect 91612 836 93860 864
rect 91612 824 91618 836
rect 93854 824 93860 836
rect 93912 824 93918 876
rect 97258 824 97264 876
rect 97316 864 97322 876
rect 116670 864 116676 876
rect 97316 836 116676 864
rect 97316 824 97322 836
rect 116670 824 116676 836
rect 116728 824 116734 876
rect 109034 756 109040 808
rect 109092 796 109098 808
rect 117222 796 117228 808
rect 109092 768 117228 796
rect 109092 756 109098 768
rect 117222 756 117228 768
rect 117280 756 117286 808
rect 103790 688 103796 740
rect 103848 728 103854 740
rect 110782 728 110788 740
rect 103848 700 110788 728
rect 103848 688 103854 700
rect 110782 688 110788 700
rect 110840 688 110846 740
<< via1 >>
rect 63408 160012 63460 160064
rect 146484 160012 146536 160064
rect 146760 160012 146812 160064
rect 154488 160012 154540 160064
rect 156788 160012 156840 160064
rect 191748 160012 191800 160064
rect 197176 160012 197228 160064
rect 207112 160012 207164 160064
rect 211436 160012 211488 160064
rect 280160 160012 280212 160064
rect 281264 160012 281316 160064
rect 332692 160012 332744 160064
rect 335084 160012 335136 160064
rect 338488 160012 338540 160064
rect 339684 160012 339736 160064
rect 374368 160012 374420 160064
rect 378876 160012 378928 160064
rect 398104 160012 398156 160064
rect 409972 160012 410024 160064
rect 417608 160012 417660 160064
rect 454592 160012 454644 160064
rect 465448 160012 465500 160064
rect 25596 159944 25648 159996
rect 109776 159944 109828 159996
rect 117228 159944 117280 159996
rect 191656 159944 191708 159996
rect 198004 159944 198056 159996
rect 269856 159944 269908 159996
rect 271236 159944 271288 159996
rect 272524 159944 272576 159996
rect 275376 159944 275428 159996
rect 328460 159944 328512 159996
rect 329196 159944 329248 159996
rect 369860 159944 369912 159996
rect 374644 159944 374696 159996
rect 388352 159944 388404 159996
rect 389824 159944 389876 159996
rect 413928 159944 413980 159996
rect 452844 159944 452896 159996
rect 464252 159944 464304 159996
rect 468024 159944 468076 159996
rect 476028 159944 476080 159996
rect 76932 159876 76984 159928
rect 162584 159876 162636 159928
rect 166908 159876 166960 159928
rect 186412 159876 186464 159928
rect 191288 159876 191340 159928
rect 264888 159876 264940 159928
rect 268660 159876 268712 159928
rect 323676 159876 323728 159928
rect 328368 159876 328420 159928
rect 369216 159876 369268 159928
rect 372160 159876 372212 159928
rect 396264 159876 396316 159928
rect 403256 159876 403308 159928
rect 416596 159876 416648 159928
rect 455420 159876 455472 159928
rect 466644 159876 466696 159928
rect 467196 159876 467248 159928
rect 473360 159876 473412 159928
rect 70124 159808 70176 159860
rect 156420 159808 156472 159860
rect 156604 159808 156656 159860
rect 160100 159808 160152 159860
rect 56692 159740 56744 159792
rect 137284 159740 137336 159792
rect 137376 159740 137428 159792
rect 139676 159740 139728 159792
rect 139952 159740 140004 159792
rect 147036 159740 147088 159792
rect 153476 159740 153528 159792
rect 180708 159808 180760 159860
rect 184572 159808 184624 159860
rect 259552 159808 259604 159860
rect 261944 159808 261996 159860
rect 312360 159808 312412 159860
rect 312452 159808 312504 159860
rect 313372 159808 313424 159860
rect 322480 159808 322532 159860
rect 364800 159808 364852 159860
rect 376300 159808 376352 159860
rect 405832 159808 405884 159860
rect 449532 159808 449584 159860
rect 459560 159808 459612 159860
rect 472256 159808 472308 159860
rect 479064 159808 479116 159860
rect 177856 159740 177908 159792
rect 254308 159740 254360 159792
rect 255228 159740 255280 159792
rect 313464 159740 313516 159792
rect 314108 159740 314160 159792
rect 357992 159740 358044 159792
rect 365444 159740 365496 159792
rect 395436 159740 395488 159792
rect 396540 159740 396592 159792
rect 413836 159740 413888 159792
rect 420920 159740 420972 159792
rect 440424 159740 440476 159792
rect 453764 159740 453816 159792
rect 464988 159740 465040 159792
rect 18880 159672 18932 159724
rect 109132 159672 109184 159724
rect 113088 159672 113140 159724
rect 126428 159672 126480 159724
rect 126520 159672 126572 159724
rect 156512 159672 156564 159724
rect 49976 159604 50028 159656
rect 143264 159604 143316 159656
rect 143356 159604 143408 159656
rect 156604 159604 156656 159656
rect 43260 159536 43312 159588
rect 136824 159536 136876 159588
rect 137284 159536 137336 159588
rect 144000 159536 144052 159588
rect 144184 159536 144236 159588
rect 36544 159468 36596 159520
rect 32312 159400 32364 159452
rect 126244 159400 126296 159452
rect 126428 159468 126480 159520
rect 127624 159468 127676 159520
rect 129924 159468 129976 159520
rect 146760 159468 146812 159520
rect 147220 159536 147272 159588
rect 164148 159672 164200 159724
rect 167736 159672 167788 159724
rect 246580 159672 246632 159724
rect 248512 159672 248564 159724
rect 308128 159672 308180 159724
rect 308220 159672 308272 159724
rect 161020 159604 161072 159656
rect 241428 159604 241480 159656
rect 244280 159604 244332 159656
rect 305184 159604 305236 159656
rect 309048 159604 309100 159656
rect 342720 159672 342772 159724
rect 343824 159672 343876 159724
rect 347780 159672 347832 159724
rect 378600 159672 378652 159724
rect 379704 159672 379756 159724
rect 405924 159672 405976 159724
rect 414204 159672 414256 159724
rect 434812 159672 434864 159724
rect 446128 159672 446180 159724
rect 456800 159672 456852 159724
rect 458732 159672 458784 159724
rect 465080 159672 465132 159724
rect 470508 159672 470560 159724
rect 476120 159672 476172 159724
rect 478972 159672 479024 159724
rect 484676 159672 484728 159724
rect 157616 159536 157668 159588
rect 239128 159536 239180 159588
rect 250996 159536 251048 159588
rect 310612 159536 310664 159588
rect 315764 159536 315816 159588
rect 342260 159536 342312 159588
rect 147404 159468 147456 159520
rect 129740 159400 129792 159452
rect 130752 159400 130804 159452
rect 137192 159400 137244 159452
rect 6276 159332 6328 159384
rect 122840 159332 122892 159384
rect 123116 159332 123168 159384
rect 144184 159400 144236 159452
rect 144368 159400 144420 159452
rect 225236 159468 225288 159520
rect 231676 159468 231728 159520
rect 295432 159468 295484 159520
rect 295616 159468 295668 159520
rect 335820 159468 335872 159520
rect 147588 159400 147640 159452
rect 149336 159400 149388 159452
rect 150900 159400 150952 159452
rect 233884 159400 233936 159452
rect 234988 159400 235040 159452
rect 298008 159400 298060 159452
rect 301504 159400 301556 159452
rect 336188 159468 336240 159520
rect 353392 159604 353444 159656
rect 357440 159604 357492 159656
rect 363236 159604 363288 159656
rect 369584 159604 369636 159656
rect 400680 159604 400732 159656
rect 407488 159604 407540 159656
rect 429568 159604 429620 159656
rect 450360 159604 450412 159656
rect 462228 159604 462280 159656
rect 468852 159604 468904 159656
rect 474832 159604 474884 159656
rect 477316 159604 477368 159656
rect 483296 159604 483348 159656
rect 342444 159536 342496 159588
rect 359648 159536 359700 159588
rect 362868 159536 362920 159588
rect 395252 159536 395304 159588
rect 399024 159536 399076 159588
rect 408592 159536 408644 159588
rect 410800 159536 410852 159588
rect 432144 159536 432196 159588
rect 451188 159536 451240 159588
rect 461492 159536 461544 159588
rect 463792 159536 463844 159588
rect 471520 159536 471572 159588
rect 479800 159536 479852 159588
rect 484860 159536 484912 159588
rect 341432 159400 341484 159452
rect 354772 159468 354824 159520
rect 358636 159468 358688 159520
rect 392400 159468 392452 159520
rect 424324 159468 424376 159520
rect 442448 159468 442500 159520
rect 452016 159468 452068 159520
rect 463608 159468 463660 159520
rect 465540 159468 465592 159520
rect 472256 159468 472308 159520
rect 343456 159400 343508 159452
rect 137468 159332 137520 159384
rect 223580 159332 223632 159384
rect 224960 159332 225012 159384
rect 290280 159332 290332 159384
rect 294788 159332 294840 159384
rect 336004 159332 336056 159384
rect 336096 159332 336148 159384
rect 342260 159332 342312 159384
rect 342352 159332 342404 159384
rect 348792 159400 348844 159452
rect 356152 159400 356204 159452
rect 390560 159400 390612 159452
rect 404084 159400 404136 159452
rect 426992 159400 427044 159452
rect 427636 159400 427688 159452
rect 445024 159400 445076 159452
rect 447876 159400 447928 159452
rect 460112 159400 460164 159452
rect 518348 159400 518400 159452
rect 523500 159400 523552 159452
rect 346032 159332 346084 159384
rect 382740 159332 382792 159384
rect 383108 159332 383160 159384
rect 411352 159332 411404 159384
rect 417516 159332 417568 159384
rect 437664 159332 437716 159384
rect 448704 159332 448756 159384
rect 461216 159332 461268 159384
rect 461308 159332 461360 159384
rect 468024 159332 468076 159384
rect 469680 159332 469732 159384
rect 477408 159332 477460 159384
rect 478144 159332 478196 159384
rect 483664 159332 483716 159384
rect 517612 159332 517664 159384
rect 522672 159332 522724 159384
rect 73528 159264 73580 159316
rect 80060 159264 80112 159316
rect 83648 159264 83700 159316
rect 167000 159264 167052 159316
rect 170220 159264 170272 159316
rect 198924 159264 198976 159316
rect 201408 159264 201460 159316
rect 212632 159264 212684 159316
rect 214012 159264 214064 159316
rect 282000 159264 282052 159316
rect 282092 159264 282144 159316
rect 333980 159264 334032 159316
rect 334256 159264 334308 159316
rect 374000 159264 374052 159316
rect 388996 159264 389048 159316
rect 404176 159264 404228 159316
rect 457904 159264 457956 159316
rect 468116 159264 468168 159316
rect 80244 159196 80296 159248
rect 91100 159196 91152 159248
rect 100484 159196 100536 159248
rect 184664 159196 184716 159248
rect 187056 159196 187108 159248
rect 214656 159196 214708 159248
rect 218244 159196 218296 159248
rect 285128 159196 285180 159248
rect 287980 159196 288032 159248
rect 338396 159196 338448 159248
rect 339316 159196 339368 159248
rect 377588 159196 377640 159248
rect 385592 159196 385644 159248
rect 398932 159196 398984 159248
rect 400772 159196 400824 159248
rect 424508 159196 424560 159248
rect 457076 159196 457128 159248
rect 467840 159196 467892 159248
rect 86960 159128 87012 159180
rect 93676 159060 93728 159112
rect 162860 159060 162912 159112
rect 163044 159128 163096 159180
rect 172428 159128 172480 159180
rect 193772 159128 193824 159180
rect 218060 159128 218112 159180
rect 220728 159128 220780 159180
rect 283196 159128 283248 159180
rect 284668 159128 284720 159180
rect 285772 159128 285824 159180
rect 169852 159060 169904 159112
rect 171140 159060 171192 159112
rect 172704 159060 172756 159112
rect 173624 159060 173676 159112
rect 197360 159060 197412 159112
rect 224132 159060 224184 159112
rect 288164 159128 288216 159180
rect 288900 159128 288952 159180
rect 339040 159128 339092 159180
rect 341432 159128 341484 159180
rect 348700 159128 348752 159180
rect 348792 159128 348844 159180
rect 374092 159128 374144 159180
rect 302332 159060 302384 159112
rect 349252 159060 349304 159112
rect 107200 158992 107252 159044
rect 182548 158992 182600 159044
rect 183744 158992 183796 159044
rect 200488 158992 200540 159044
rect 200580 158992 200632 159044
rect 224960 158992 225012 159044
rect 230848 158992 230900 159044
rect 294788 158992 294840 159044
rect 298100 158992 298152 159044
rect 299664 158992 299716 159044
rect 307392 158992 307444 159044
rect 351828 159060 351880 159112
rect 351920 159060 351972 159112
rect 385408 159128 385460 159180
rect 392308 159128 392360 159180
rect 404268 159128 404320 159180
rect 456248 159128 456300 159180
rect 466920 159128 466972 159180
rect 378048 159060 378100 159112
rect 388444 159060 388496 159112
rect 395712 159060 395764 159112
rect 405464 159060 405516 159112
rect 460480 159060 460532 159112
rect 466552 159060 466604 159112
rect 471428 159060 471480 159112
rect 478420 159060 478472 159112
rect 351092 158992 351144 159044
rect 382372 158992 382424 159044
rect 459652 158992 459704 159044
rect 466460 158992 466512 159044
rect 473912 158992 473964 159044
rect 480352 158992 480404 159044
rect 480628 158992 480680 159044
rect 485964 158992 486016 159044
rect 96252 158924 96304 158976
rect 121644 158924 121696 158976
rect 124036 158924 124088 158976
rect 193404 158924 193456 158976
rect 194692 158924 194744 158976
rect 203708 158924 203760 158976
rect 207296 158924 207348 158976
rect 230756 158924 230808 158976
rect 237564 158924 237616 158976
rect 299480 158924 299532 158976
rect 314936 158924 314988 158976
rect 357532 158924 357584 158976
rect 357808 158924 357860 158976
rect 384948 158924 385000 158976
rect 409144 158924 409196 158976
rect 410892 158924 410944 158976
rect 413376 158924 413428 158976
rect 419724 158924 419776 158976
rect 462136 158924 462188 158976
rect 467932 158924 467984 158976
rect 475568 158924 475620 158976
rect 481732 158924 481784 158976
rect 506664 158924 506716 158976
rect 508412 158924 508464 158976
rect 102968 158856 103020 158908
rect 125508 158856 125560 158908
rect 109684 158788 109736 158840
rect 137100 158856 137152 158908
rect 137192 158856 137244 158908
rect 195428 158856 195480 158908
rect 208124 158856 208176 158908
rect 212448 158856 212500 158908
rect 217324 158856 217376 158908
rect 220728 158856 220780 158908
rect 241796 158856 241848 158908
rect 303252 158856 303304 158908
rect 305644 158856 305696 158908
rect 307392 158856 307444 158908
rect 310704 158856 310756 158908
rect 311992 158856 312044 158908
rect 312360 158856 312412 158908
rect 318800 158856 318852 158908
rect 320824 158856 320876 158908
rect 133236 158788 133288 158840
rect 158720 158788 158772 158840
rect 163504 158788 163556 158840
rect 197268 158788 197320 158840
rect 203892 158788 203944 158840
rect 213644 158788 213696 158840
rect 214840 158788 214892 158840
rect 222108 158788 222160 158840
rect 238392 158788 238444 158840
rect 241612 158788 241664 158840
rect 261116 158788 261168 158840
rect 316316 158788 316368 158840
rect 319168 158788 319220 158840
rect 90364 158720 90416 158772
rect 92572 158720 92624 158772
rect 92848 158720 92900 158772
rect 114468 158720 114520 158772
rect 119804 158720 119856 158772
rect 146576 158720 146628 158772
rect 146668 158720 146720 158772
rect 176660 158720 176712 158772
rect 180340 158720 180392 158772
rect 204904 158720 204956 158772
rect 210608 158720 210660 158772
rect 215392 158720 215444 158772
rect 221556 158720 221608 158772
rect 224040 158720 224092 158772
rect 240876 158720 240928 158772
rect 243360 158720 243412 158772
rect 254400 158720 254452 158772
rect 255412 158720 255464 158772
rect 258540 158720 258592 158772
rect 260840 158720 260892 158772
rect 264428 158720 264480 158772
rect 266360 158720 266412 158772
rect 267832 158720 267884 158772
rect 320272 158720 320324 158772
rect 321652 158788 321704 158840
rect 357440 158788 357492 158840
rect 361212 158856 361264 158908
rect 385132 158856 385184 158908
rect 391480 158856 391532 158908
rect 394608 158856 394660 158908
rect 412548 158856 412600 158908
rect 413100 158856 413152 158908
rect 420092 158856 420144 158908
rect 423588 158856 423640 158908
rect 462964 158856 463016 158908
rect 469220 158856 469272 158908
rect 474740 158856 474792 158908
rect 481088 158856 481140 158908
rect 482284 158856 482336 158908
rect 487252 158856 487304 158908
rect 507952 158856 508004 158908
rect 510068 158856 510120 158908
rect 362960 158788 363012 158840
rect 367928 158788 367980 158840
rect 327540 158720 327592 158772
rect 368388 158720 368440 158772
rect 386328 158788 386380 158840
rect 374184 158720 374236 158772
rect 379428 158720 379480 158772
rect 384764 158720 384816 158772
rect 389180 158788 389232 158840
rect 405740 158788 405792 158840
rect 409236 158788 409288 158840
rect 416688 158788 416740 158840
rect 419632 158788 419684 158840
rect 466368 158788 466420 158840
rect 472440 158788 472492 158840
rect 476396 158788 476448 158840
rect 482376 158788 482428 158840
rect 506112 158788 506164 158840
rect 507584 158788 507636 158840
rect 388076 158720 388128 158772
rect 390376 158720 390428 158772
rect 464620 158720 464672 158772
rect 471244 158720 471296 158772
rect 473084 158720 473136 158772
rect 479708 158720 479760 158772
rect 481456 158720 481508 158772
rect 486148 158720 486200 158772
rect 505376 158720 505428 158772
rect 506756 158720 506808 158772
rect 509332 158720 509384 158772
rect 511724 158720 511776 158772
rect 514944 158720 514996 158772
rect 518532 158720 518584 158772
rect 81072 158652 81124 158704
rect 180892 158652 180944 158704
rect 181996 158652 182048 158704
rect 257528 158652 257580 158704
rect 321560 158652 321612 158704
rect 67640 158584 67692 158636
rect 170220 158584 170272 158636
rect 171968 158584 172020 158636
rect 249800 158584 249852 158636
rect 74356 158516 74408 158568
rect 175372 158516 175424 158568
rect 178684 158516 178736 158568
rect 255596 158516 255648 158568
rect 71044 158448 71096 158500
rect 172796 158448 172848 158500
rect 175280 158448 175332 158500
rect 252560 158448 252612 158500
rect 60924 158380 60976 158432
rect 165068 158380 165120 158432
rect 165252 158380 165304 158432
rect 244648 158380 244700 158432
rect 64236 158312 64288 158364
rect 167552 158312 167604 158364
rect 168564 158312 168616 158364
rect 247132 158312 247184 158364
rect 54208 158244 54260 158296
rect 160284 158244 160336 158296
rect 161848 158244 161900 158296
rect 242072 158244 242124 158296
rect 50804 158176 50856 158228
rect 157340 158176 157392 158228
rect 158444 158176 158496 158228
rect 239680 158176 239732 158228
rect 256884 158176 256936 158228
rect 314752 158176 314804 158228
rect 47492 158108 47544 158160
rect 154764 158108 154816 158160
rect 155132 158108 155184 158160
rect 237380 158108 237432 158160
rect 246764 158108 246816 158160
rect 306932 158108 306984 158160
rect 37372 158040 37424 158092
rect 146760 158040 146812 158092
rect 148416 158040 148468 158092
rect 231952 158040 232004 158092
rect 243452 158040 243504 158092
rect 304356 158040 304408 158092
rect 388 157972 440 158024
rect 118884 157972 118936 158024
rect 131580 157972 131632 158024
rect 218980 157972 219032 158024
rect 236736 157972 236788 158024
rect 299572 157972 299624 158024
rect 77760 157904 77812 157956
rect 84476 157836 84528 157888
rect 175924 157836 175976 157888
rect 176200 157904 176252 157956
rect 183008 157904 183060 157956
rect 185400 157904 185452 157956
rect 260104 157904 260156 157956
rect 178040 157836 178092 157888
rect 180708 157836 180760 157888
rect 181352 157836 181404 157888
rect 181536 157836 181588 157888
rect 188160 157836 188212 157888
rect 188804 157836 188856 157888
rect 262680 157836 262732 157888
rect 87788 157768 87840 157820
rect 91192 157700 91244 157752
rect 181076 157700 181128 157752
rect 94596 157632 94648 157684
rect 181168 157632 181220 157684
rect 181812 157768 181864 157820
rect 190644 157768 190696 157820
rect 195520 157768 195572 157820
rect 267740 157768 267792 157820
rect 181720 157700 181772 157752
rect 185584 157632 185636 157684
rect 190460 157700 190512 157752
rect 264060 157700 264112 157752
rect 236092 157632 236144 157684
rect 97908 157564 97960 157616
rect 193220 157564 193272 157616
rect 197360 157564 197412 157616
rect 251272 157564 251324 157616
rect 111340 157496 111392 157548
rect 203432 157496 203484 157548
rect 204904 157496 204956 157548
rect 255872 157496 255924 157548
rect 114744 157428 114796 157480
rect 206192 157428 206244 157480
rect 141700 157360 141752 157412
rect 226708 157360 226760 157412
rect 49148 157292 49200 157344
rect 156052 157292 156104 157344
rect 158720 157292 158772 157344
rect 214472 157292 214524 157344
rect 214564 157292 214616 157344
rect 221372 157292 221424 157344
rect 224224 157292 224276 157344
rect 281632 157292 281684 157344
rect 45744 157224 45796 157276
rect 153568 157224 153620 157276
rect 164148 157224 164200 157276
rect 166264 157224 166316 157276
rect 192116 157224 192168 157276
rect 265164 157224 265216 157276
rect 283840 157224 283892 157276
rect 335452 157224 335504 157276
rect 39028 157156 39080 157208
rect 148232 157156 148284 157208
rect 150072 157156 150124 157208
rect 233516 157156 233568 157208
rect 290556 157156 290608 157208
rect 340052 157156 340104 157208
rect 42432 157088 42484 157140
rect 150900 157088 150952 157140
rect 156512 157088 156564 157140
rect 158904 157088 158956 157140
rect 160100 157088 160152 157140
rect 165896 157088 165948 157140
rect 165988 157088 166040 157140
rect 171600 157088 171652 157140
rect 177028 157088 177080 157140
rect 254032 157088 254084 157140
rect 287152 157088 287204 157140
rect 338120 157088 338172 157140
rect 35716 157020 35768 157072
rect 145932 157020 145984 157072
rect 151728 157020 151780 157072
rect 234804 157020 234856 157072
rect 280436 157020 280488 157072
rect 332876 157020 332928 157072
rect 24768 156952 24820 157004
rect 137376 156952 137428 157004
rect 138296 156952 138348 157004
rect 224132 156952 224184 157004
rect 273720 156952 273772 157004
rect 327540 156952 327592 157004
rect 18052 156884 18104 156936
rect 132500 156884 132552 156936
rect 134892 156884 134944 156936
rect 214564 156884 214616 156936
rect 224960 156884 225012 156936
rect 272064 156884 272116 156936
rect 277124 156884 277176 156936
rect 330024 156884 330076 156936
rect 21364 156816 21416 156868
rect 135260 156816 135312 156868
rect 135812 156816 135864 156868
rect 222384 156816 222436 156868
rect 226616 156816 226668 156868
rect 291568 156816 291620 156868
rect 300676 156816 300728 156868
rect 348056 156816 348108 156868
rect 14648 156748 14700 156800
rect 129832 156748 129884 156800
rect 139124 156748 139176 156800
rect 225144 156748 225196 156800
rect 230020 156748 230072 156800
rect 294052 156748 294104 156800
rect 297272 156748 297324 156800
rect 345572 156748 345624 156800
rect 11244 156680 11296 156732
rect 127164 156680 127216 156732
rect 128176 156680 128228 156732
rect 216680 156680 216732 156732
rect 223212 156680 223264 156732
rect 288992 156680 289044 156732
rect 293868 156680 293920 156732
rect 342812 156680 342864 156732
rect 2044 156612 2096 156664
rect 120172 156612 120224 156664
rect 124864 156612 124916 156664
rect 213920 156612 213972 156664
rect 216496 156612 216548 156664
rect 283104 156612 283156 156664
rect 52460 156544 52512 156596
rect 158812 156544 158864 156596
rect 158904 156544 158956 156596
rect 200764 156544 200816 156596
rect 200948 156544 201000 156596
rect 270500 156544 270552 156596
rect 59268 156476 59320 156528
rect 163780 156476 163832 156528
rect 165896 156476 165948 156528
rect 69296 156408 69348 156460
rect 165988 156408 166040 156460
rect 166264 156476 166316 156528
rect 225512 156476 225564 156528
rect 228088 156408 228140 156460
rect 82820 156340 82872 156392
rect 181812 156340 181864 156392
rect 198832 156340 198884 156392
rect 200948 156340 201000 156392
rect 209780 156340 209832 156392
rect 278964 156340 279016 156392
rect 101312 156272 101364 156324
rect 196164 156272 196216 156324
rect 200764 156272 200816 156324
rect 99564 156204 99616 156256
rect 194692 156204 194744 156256
rect 198004 156204 198056 156256
rect 211344 156204 211396 156256
rect 108028 156136 108080 156188
rect 200672 156136 200724 156188
rect 118148 156068 118200 156120
rect 208768 156136 208820 156188
rect 213184 156272 213236 156324
rect 224224 156272 224276 156324
rect 214472 156204 214524 156256
rect 219992 156204 220044 156256
rect 220084 156204 220136 156256
rect 286232 156272 286284 156324
rect 215484 156136 215536 156188
rect 218060 156136 218112 156188
rect 266544 156204 266596 156256
rect 230756 156136 230808 156188
rect 276756 156136 276808 156188
rect 203064 156068 203116 156120
rect 273536 156068 273588 156120
rect 121460 156000 121512 156052
rect 198004 156000 198056 156052
rect 202236 156000 202288 156052
rect 273352 156000 273404 156052
rect 145012 155932 145064 155984
rect 229284 155932 229336 155984
rect 66812 155864 66864 155916
rect 82912 155864 82964 155916
rect 92020 155864 92072 155916
rect 60096 155796 60148 155848
rect 78772 155796 78824 155848
rect 88708 155796 88760 155848
rect 186412 155796 186464 155848
rect 186596 155864 186648 155916
rect 194048 155864 194100 155916
rect 196348 155864 196400 155916
rect 268476 155864 268528 155916
rect 296444 155864 296496 155916
rect 345204 155864 345256 155916
rect 189080 155796 189132 155848
rect 192944 155796 192996 155848
rect 265900 155796 265952 155848
rect 293040 155796 293092 155848
rect 342352 155796 342404 155848
rect 12164 155728 12216 155780
rect 110328 155728 110380 155780
rect 112260 155728 112312 155780
rect 204352 155728 204404 155780
rect 206468 155728 206520 155780
rect 276112 155728 276164 155780
rect 289728 155728 289780 155780
rect 339592 155728 339644 155780
rect 46572 155660 46624 155712
rect 75092 155660 75144 155712
rect 81900 155660 81952 155712
rect 181168 155660 181220 155712
rect 186228 155660 186280 155712
rect 260932 155660 260984 155712
rect 270316 155660 270368 155712
rect 324964 155660 325016 155712
rect 340972 155660 341024 155712
rect 378692 155660 378744 155712
rect 53380 155592 53432 155644
rect 66628 155592 66680 155644
rect 71872 155592 71924 155644
rect 173532 155592 173584 155644
rect 176292 155592 176344 155644
rect 253020 155592 253072 155644
rect 267004 155592 267056 155644
rect 322112 155592 322164 155644
rect 344376 155592 344428 155644
rect 381452 155592 381504 155644
rect 39856 155524 39908 155576
rect 68928 155524 68980 155576
rect 75184 155524 75236 155576
rect 176016 155524 176068 155576
rect 179512 155524 179564 155576
rect 255688 155524 255740 155576
rect 263600 155524 263652 155576
rect 320180 155524 320232 155576
rect 337660 155524 337712 155576
rect 376300 155524 376352 155576
rect 65156 155456 65208 155508
rect 168564 155456 168616 155508
rect 169392 155456 169444 155508
rect 247868 155456 247920 155508
rect 260288 155456 260340 155508
rect 317604 155456 317656 155508
rect 333428 155456 333480 155508
rect 373080 155456 373132 155508
rect 7932 155388 7984 155440
rect 124588 155388 124640 155440
rect 145840 155388 145892 155440
rect 230020 155388 230072 155440
rect 253572 155388 253624 155440
rect 312084 155388 312136 155440
rect 330116 155388 330168 155440
rect 370504 155388 370556 155440
rect 8760 155320 8812 155372
rect 125784 155320 125836 155372
rect 142528 155320 142580 155372
rect 227904 155320 227956 155372
rect 250168 155320 250220 155372
rect 309508 155320 309560 155372
rect 319996 155320 320048 155372
rect 363144 155320 363196 155372
rect 4528 155252 4580 155304
rect 122012 155252 122064 155304
rect 129004 155252 129056 155304
rect 217048 155252 217100 155304
rect 233332 155252 233384 155304
rect 296812 155252 296864 155304
rect 299756 155252 299808 155304
rect 347964 155252 348016 155304
rect 373816 155252 373868 155304
rect 403532 155252 403584 155304
rect 5356 155184 5408 155236
rect 122932 155184 122984 155236
rect 125692 155184 125744 155236
rect 214472 155184 214524 155236
rect 240048 155184 240100 155236
rect 302516 155184 302568 155236
rect 306564 155184 306616 155236
rect 352472 155184 352524 155236
rect 370412 155184 370464 155236
rect 401784 155184 401836 155236
rect 89536 155116 89588 155168
rect 186964 155116 187016 155168
rect 189632 155116 189684 155168
rect 263692 155116 263744 155168
rect 95424 155048 95476 155100
rect 98736 154980 98788 155032
rect 186320 154980 186372 155032
rect 186780 155048 186832 155100
rect 191472 154980 191524 155032
rect 199660 155048 199712 155100
rect 271052 155048 271104 155100
rect 303160 155048 303212 155100
rect 349988 155048 350040 155100
rect 200212 154980 200264 155032
rect 207112 154980 207164 155032
rect 269304 154980 269356 155032
rect 15476 154912 15528 154964
rect 109040 154912 109092 154964
rect 122288 154912 122340 154964
rect 211988 154912 212040 154964
rect 214656 154912 214708 154964
rect 261484 154912 261536 154964
rect 106372 154844 106424 154896
rect 186596 154844 186648 154896
rect 186688 154844 186740 154896
rect 245844 154844 245896 154896
rect 110512 154776 110564 154828
rect 139308 154776 139360 154828
rect 149244 154776 149296 154828
rect 232504 154776 232556 154828
rect 109132 154708 109184 154760
rect 132960 154708 133012 154760
rect 155960 154708 156012 154760
rect 237656 154708 237708 154760
rect 156328 154640 156380 154692
rect 118608 154572 118660 154624
rect 119712 154572 119764 154624
rect 154488 154572 154540 154624
rect 51080 154504 51132 154556
rect 154948 154504 155000 154556
rect 156696 154572 156748 154624
rect 162676 154640 162728 154692
rect 242900 154640 242952 154692
rect 159364 154572 159416 154624
rect 240232 154572 240284 154624
rect 212724 154504 212776 154556
rect 218336 154504 218388 154556
rect 44180 154436 44232 154488
rect 142896 154436 142948 154488
rect 142988 154436 143040 154488
rect 191104 154436 191156 154488
rect 114468 154368 114520 154420
rect 118608 154368 118660 154420
rect 118700 154368 118752 154420
rect 119620 154368 119672 154420
rect 119712 154368 119764 154420
rect 189540 154368 189592 154420
rect 191012 154368 191064 154420
rect 202420 154436 202472 154488
rect 215300 154436 215352 154488
rect 280252 154436 280304 154488
rect 280620 154504 280672 154556
rect 283288 154572 283340 154624
rect 285588 154504 285640 154556
rect 285680 154504 285732 154556
rect 337200 154504 337252 154556
rect 353668 154504 353720 154556
rect 388628 154504 388680 154556
rect 283380 154436 283432 154488
rect 334624 154436 334676 154488
rect 349528 154436 349580 154488
rect 386052 154436 386104 154488
rect 390652 154436 390704 154488
rect 416872 154436 416924 154488
rect 191288 154368 191340 154420
rect 201776 154368 201828 154420
rect 204996 154368 205048 154420
rect 275560 154368 275612 154420
rect 276204 154368 276256 154420
rect 329932 154368 329984 154420
rect 346400 154368 346452 154420
rect 383752 154368 383804 154420
rect 393320 154368 393372 154420
rect 419540 154368 419592 154420
rect 34520 154300 34572 154352
rect 137928 154300 137980 154352
rect 138112 154300 138164 154352
rect 139492 154300 139544 154352
rect 139676 154300 139728 154352
rect 37924 154232 37976 154284
rect 143080 154300 143132 154352
rect 205088 154300 205140 154352
rect 208400 154300 208452 154352
rect 278136 154300 278188 154352
rect 278872 154300 278924 154352
rect 332140 154300 332192 154352
rect 339500 154300 339552 154352
rect 378324 154300 378376 154352
rect 397368 154300 397420 154352
rect 422484 154300 422536 154352
rect 27252 154164 27304 154216
rect 137008 154164 137060 154216
rect 23480 154096 23532 154148
rect 136916 154096 136968 154148
rect 13820 154028 13872 154080
rect 129188 154028 129240 154080
rect 9680 153960 9732 154012
rect 126612 153960 126664 154012
rect 127624 153960 127676 154012
rect 129280 153960 129332 154012
rect 7104 153892 7156 153944
rect 124220 153892 124272 153944
rect 125508 153892 125560 153944
rect 129464 153960 129516 154012
rect 142436 154096 142488 154148
rect 145380 154232 145432 154284
rect 146944 154232 146996 154284
rect 147956 154232 148008 154284
rect 148048 154232 148100 154284
rect 156328 154232 156380 154284
rect 142896 154164 142948 154216
rect 153292 154164 153344 154216
rect 156788 154232 156840 154284
rect 137284 154028 137336 154080
rect 138020 154028 138072 154080
rect 147864 154096 147916 154148
rect 147956 154096 148008 154148
rect 142988 154028 143040 154080
rect 143448 154028 143500 154080
rect 150440 154028 150492 154080
rect 151912 154096 151964 154148
rect 156512 154164 156564 154216
rect 163228 154232 163280 154284
rect 176660 154232 176712 154284
rect 179512 154232 179564 154284
rect 182180 154232 182232 154284
rect 258264 154232 258316 154284
rect 262220 154232 262272 154284
rect 319260 154232 319312 154284
rect 343548 154232 343600 154284
rect 380992 154232 381044 154284
rect 386512 154232 386564 154284
rect 414204 154232 414256 154284
rect 162676 154164 162728 154216
rect 165804 154164 165856 154216
rect 172520 154164 172572 154216
rect 250536 154164 250588 154216
rect 255320 154164 255372 154216
rect 314108 154164 314160 154216
rect 336832 154164 336884 154216
rect 375748 154164 375800 154216
rect 383660 154164 383712 154216
rect 411720 154164 411772 154216
rect 154948 154096 155000 154148
rect 158076 154096 158128 154148
rect 160192 154096 160244 154148
rect 162768 154028 162820 154080
rect 165620 154096 165672 154148
rect 245660 154096 245712 154148
rect 245936 154096 245988 154148
rect 306380 154096 306432 154148
rect 326712 154096 326764 154148
rect 368020 154096 368072 154148
rect 376852 154096 376904 154148
rect 406568 154096 406620 154148
rect 240968 154028 241020 154080
rect 248604 154028 248656 154080
rect 309232 154028 309284 154080
rect 323308 154028 323360 154080
rect 365812 154028 365864 154080
rect 380164 154028 380216 154080
rect 409144 154028 409196 154080
rect 132408 153892 132460 153944
rect 137468 153892 137520 153944
rect 219716 153960 219768 154012
rect 222476 153960 222528 154012
rect 288440 153960 288492 154012
rect 316040 153960 316092 154012
rect 360384 153960 360436 154012
rect 367100 153960 367152 154012
rect 398840 153960 398892 154012
rect 480 153824 532 153876
rect 119528 153824 119580 153876
rect 119620 153824 119672 153876
rect 138204 153824 138256 153876
rect 143540 153892 143592 153944
rect 145288 153892 145340 153944
rect 145380 153892 145432 153944
rect 222936 153892 222988 153944
rect 225052 153892 225104 153944
rect 291292 153892 291344 153944
rect 313280 153892 313332 153944
rect 357808 153892 357860 153944
rect 363052 153892 363104 153944
rect 396356 153892 396408 153944
rect 401600 153892 401652 153944
rect 425336 153892 425388 153944
rect 48320 153756 48372 153808
rect 155500 153756 155552 153808
rect 156788 153824 156840 153876
rect 235172 153824 235224 153876
rect 241888 153824 241940 153876
rect 303804 153824 303856 153876
rect 309140 153824 309192 153876
rect 355232 153824 355284 153876
rect 356244 153824 356296 153876
rect 391204 153824 391256 153876
rect 397460 153824 397512 153876
rect 422668 153824 422720 153876
rect 191012 153756 191064 153808
rect 191104 153756 191156 153808
rect 197360 153756 197412 153808
rect 197452 153756 197504 153808
rect 199292 153756 199344 153808
rect 61108 153688 61160 153740
rect 162676 153688 162728 153740
rect 162768 153688 162820 153740
rect 210148 153756 210200 153808
rect 231860 153756 231912 153808
rect 296168 153756 296220 153808
rect 360476 153756 360528 153808
rect 393780 153756 393832 153808
rect 427820 153756 427872 153808
rect 432696 153756 432748 153808
rect 200488 153688 200540 153740
rect 209780 153688 209832 153740
rect 235080 153688 235132 153740
rect 298744 153688 298796 153740
rect 57980 153620 58032 153672
rect 156512 153620 156564 153672
rect 156696 153620 156748 153672
rect 218060 153620 218112 153672
rect 229100 153620 229152 153672
rect 293592 153620 293644 153672
rect 78680 153552 78732 153604
rect 179420 153552 179472 153604
rect 179512 153552 179564 153604
rect 230664 153552 230716 153604
rect 238852 153552 238904 153604
rect 301320 153552 301372 153604
rect 102140 153484 102192 153536
rect 196624 153484 196676 153536
rect 198924 153484 198976 153536
rect 248604 153484 248656 153536
rect 252652 153484 252704 153536
rect 311532 153484 311584 153536
rect 104900 153416 104952 153468
rect 199200 153416 199252 153468
rect 199292 153416 199344 153468
rect 108304 153348 108356 153400
rect 191288 153348 191340 153400
rect 191748 153348 191800 153400
rect 200120 153348 200172 153400
rect 115940 153280 115992 153332
rect 200580 153416 200632 153468
rect 258908 153416 258960 153468
rect 265440 153416 265492 153468
rect 321836 153416 321888 153468
rect 243452 153348 243504 153400
rect 259460 153348 259512 153400
rect 316776 153348 316828 153400
rect 441620 153348 441672 153400
rect 41604 153212 41656 153264
rect 138112 153212 138164 153264
rect 138204 153212 138256 153264
rect 200304 153212 200356 153264
rect 200856 153280 200908 153332
rect 238392 153280 238444 153332
rect 272892 153280 272944 153332
rect 327080 153280 327132 153332
rect 207572 153212 207624 153264
rect 269212 153212 269264 153264
rect 324412 153212 324464 153264
rect 423588 153212 423640 153264
rect 428004 153212 428056 153264
rect 23296 153144 23348 153196
rect 110972 153144 111024 153196
rect 113180 153144 113232 153196
rect 205640 153144 205692 153196
rect 215392 153144 215444 153196
rect 279424 153144 279476 153196
rect 285496 153144 285548 153196
rect 336740 153144 336792 153196
rect 339684 153144 339736 153196
rect 377036 153144 377088 153196
rect 385408 153144 385460 153196
rect 387340 153144 387392 153196
rect 389180 153144 389232 153196
rect 412640 153144 412692 153196
rect 413100 153144 413152 153196
rect 433432 153144 433484 153196
rect 433524 153144 433576 153196
rect 441804 153144 441856 153196
rect 443000 153144 443052 153196
rect 443920 153144 443972 153196
rect 450268 153144 450320 153196
rect 456800 153144 456852 153196
rect 459192 153144 459244 153196
rect 461492 153144 461544 153196
rect 463056 153144 463108 153196
rect 466460 153144 466512 153196
rect 469496 153144 469548 153196
rect 471244 153144 471296 153196
rect 473544 153144 473596 153196
rect 474832 153144 474884 153196
rect 476580 153144 476632 153196
rect 485688 153144 485740 153196
rect 489368 153144 489420 153196
rect 490748 153144 490800 153196
rect 493232 153144 493284 153196
rect 494152 153144 494204 153196
rect 496452 153144 496504 153196
rect 496636 153144 496688 153196
rect 497740 153144 497792 153196
rect 512552 153144 512604 153196
rect 514852 153144 514904 153196
rect 80060 153076 80112 153128
rect 174820 153076 174872 153128
rect 180800 153076 180852 153128
rect 256976 153076 257028 153128
rect 264980 153076 265032 153128
rect 321192 153076 321244 153128
rect 324320 153076 324372 153128
rect 366732 153076 366784 153128
rect 382188 153076 382240 153128
rect 410432 153076 410484 153128
rect 414296 153076 414348 153128
rect 103520 153008 103572 153060
rect 197912 153008 197964 153060
rect 203708 153008 203760 153060
rect 267280 153008 267332 153060
rect 272156 153008 272208 153060
rect 326344 153008 326396 153060
rect 330944 153008 330996 153060
rect 371240 153008 371292 153060
rect 372620 153008 372672 153060
rect 403348 153008 403400 153060
rect 404360 153008 404412 153060
rect 427912 153008 427964 153060
rect 430672 153076 430724 153128
rect 436284 153076 436336 153128
rect 436928 153076 436980 153128
rect 452200 153076 452252 153128
rect 466552 153076 466604 153128
rect 470140 153076 470192 153128
rect 471520 153076 471572 153128
rect 472716 153076 472768 153128
rect 473360 153076 473412 153128
rect 475292 153076 475344 153128
rect 476120 153076 476172 153128
rect 477868 153076 477920 153128
rect 484032 153076 484084 153128
rect 488080 153076 488132 153128
rect 489920 153076 489972 153128
rect 492772 153076 492824 153128
rect 494060 153076 494112 153128
rect 495808 153076 495860 153128
rect 496820 153076 496872 153128
rect 498384 153076 498436 153128
rect 511264 153076 511316 153128
rect 513472 153076 513524 153128
rect 514484 153076 514536 153128
rect 517428 153076 517480 153128
rect 431868 153008 431920 153060
rect 431960 153008 432012 153060
rect 448980 153008 449032 153060
rect 465080 153008 465132 153060
rect 468852 153008 468904 153060
rect 472440 153008 472492 153060
rect 474740 153008 474792 153060
rect 484492 153008 484544 153060
rect 488724 153008 488776 153060
rect 492680 153008 492732 153060
rect 495440 153008 495492 153060
rect 495532 153008 495584 153060
rect 497096 153008 497148 153060
rect 511724 153008 511776 153060
rect 514300 153008 514352 153060
rect 92572 152940 92624 152992
rect 187700 152940 187752 152992
rect 195428 152940 195480 152992
rect 218428 152940 218480 152992
rect 225236 152940 225288 152992
rect 228732 152940 228784 152992
rect 228824 152940 228876 152992
rect 284576 152940 284628 152992
rect 288164 152940 288216 152992
rect 289912 152940 289964 152992
rect 291384 152940 291436 152992
rect 341064 152940 341116 152992
rect 342260 152940 342312 152992
rect 344284 152940 344336 152992
rect 345296 152940 345348 152992
rect 382280 152940 382332 152992
rect 382372 152940 382424 152992
rect 386696 152940 386748 152992
rect 390376 152940 390428 152992
rect 414940 152940 414992 152992
rect 418160 152940 418212 152992
rect 432880 152940 432932 152992
rect 438860 152940 438912 152992
rect 454224 152940 454276 152992
rect 472256 152940 472308 152992
rect 474004 152940 474056 152992
rect 483204 152940 483256 152992
rect 487528 152940 487580 152992
rect 491300 152940 491352 152992
rect 494060 152940 494112 152992
rect 513196 152940 513248 152992
rect 515956 152940 516008 152992
rect 71412 152872 71464 152924
rect 92480 152872 92532 152924
rect 96620 152872 96672 152924
rect 192760 152872 192812 152924
rect 212448 152872 212500 152924
rect 277492 152872 277544 152924
rect 278780 152872 278832 152924
rect 331496 152872 331548 152924
rect 332600 152872 332652 152924
rect 372620 152872 372672 152924
rect 375472 152872 375524 152924
rect 405280 152872 405332 152924
rect 405924 152872 405976 152924
rect 408500 152872 408552 152924
rect 411260 152872 411312 152924
rect 432604 152872 432656 152924
rect 434352 152872 434404 152924
rect 441620 152872 441672 152924
rect 441712 152872 441764 152924
rect 447876 152872 447928 152924
rect 491668 152872 491720 152924
rect 494520 152872 494572 152924
rect 513840 152872 513892 152924
rect 516140 152872 516192 152924
rect 33140 152804 33192 152856
rect 138296 152804 138348 152856
rect 138572 152804 138624 152856
rect 141424 152804 141476 152856
rect 146484 152804 146536 152856
rect 167092 152804 167144 152856
rect 173900 152804 173952 152856
rect 251824 152804 251876 152856
rect 255412 152804 255464 152856
rect 312820 152804 312872 152856
rect 316316 152804 316368 152856
rect 317972 152804 318024 152856
rect 26424 152736 26476 152788
rect 138848 152736 138900 152788
rect 140872 152736 140924 152788
rect 144000 152736 144052 152788
rect 144092 152736 144144 152788
rect 161940 152736 161992 152788
rect 164332 152736 164384 152788
rect 244280 152736 244332 152788
rect 257712 152736 257764 152788
rect 315396 152736 315448 152788
rect 317420 152736 317472 152788
rect 361028 152804 361080 152856
rect 361580 152804 361632 152856
rect 395068 152804 395120 152856
rect 395436 152804 395488 152856
rect 397552 152804 397604 152856
rect 406660 152804 406712 152856
rect 429200 152804 429252 152856
rect 429384 152804 429436 152856
rect 447140 152804 447192 152856
rect 320272 152736 320324 152788
rect 323124 152736 323176 152788
rect 324228 152736 324280 152788
rect 366088 152736 366140 152788
rect 368480 152736 368532 152788
rect 400220 152736 400272 152788
rect 402428 152736 402480 152788
rect 425888 152736 425940 152788
rect 426440 152736 426492 152788
rect 444564 152736 444616 152788
rect 446312 152736 446364 152788
rect 459836 152736 459888 152788
rect 510528 152736 510580 152788
rect 512000 152736 512052 152788
rect 28172 152668 28224 152720
rect 140780 152668 140832 152720
rect 142804 152668 142856 152720
rect 149152 152668 149204 152720
rect 149336 152668 149388 152720
rect 231308 152668 231360 152720
rect 251180 152668 251232 152720
rect 310888 152668 310940 152720
rect 311992 152668 312044 152720
rect 356060 152668 356112 152720
rect 358820 152668 358872 152720
rect 393320 152668 393372 152720
rect 394884 152668 394936 152720
rect 420092 152668 420144 152720
rect 421012 152668 421064 152720
rect 22192 152600 22244 152652
rect 135628 152600 135680 152652
rect 19340 152532 19392 152584
rect 133880 152532 133932 152584
rect 136824 152532 136876 152584
rect 151820 152600 151872 152652
rect 153660 152600 153712 152652
rect 236460 152600 236512 152652
rect 247040 152600 247092 152652
rect 307760 152600 307812 152652
rect 311624 152600 311676 152652
rect 320732 152600 320784 152652
rect 320824 152600 320876 152652
rect 361672 152600 361724 152652
rect 364524 152600 364576 152652
rect 396908 152600 396960 152652
rect 399116 152600 399168 152652
rect 417424 152600 417476 152652
rect 418620 152600 418672 152652
rect 427728 152600 427780 152652
rect 138296 152532 138348 152584
rect 144000 152532 144052 152584
rect 144092 152532 144144 152584
rect 226340 152532 226392 152584
rect 2872 152464 2924 152516
rect 120816 152464 120868 152516
rect 126980 152464 127032 152516
rect 215852 152464 215904 152516
rect 220728 152464 220780 152516
rect 228824 152532 228876 152584
rect 234160 152532 234212 152584
rect 297456 152532 297508 152584
rect 303620 152532 303672 152584
rect 350724 152532 350776 152584
rect 351920 152532 351972 152584
rect 353300 152532 353352 152584
rect 354496 152532 354548 152584
rect 389272 152532 389324 152584
rect 393136 152532 393188 152584
rect 418804 152532 418856 152584
rect 418896 152532 418948 152584
rect 426900 152532 426952 152584
rect 227720 152464 227772 152516
rect 292948 152464 293000 152516
rect 298652 152464 298704 152516
rect 346860 152464 346912 152516
rect 348148 152464 348200 152516
rect 385040 152464 385092 152516
rect 386420 152464 386472 152516
rect 413652 152464 413704 152516
rect 415400 152464 415452 152516
rect 430856 152464 430908 152516
rect 432880 152668 432932 152720
rect 438032 152668 438084 152720
rect 438124 152668 438176 152720
rect 432696 152600 432748 152652
rect 438768 152600 438820 152652
rect 432972 152532 433024 152584
rect 438860 152532 438912 152584
rect 440332 152668 440384 152720
rect 455420 152668 455472 152720
rect 439044 152600 439096 152652
rect 445760 152600 445812 152652
rect 440608 152532 440660 152584
rect 442816 152532 442868 152584
rect 456800 152532 456852 152584
rect 438124 152464 438176 152516
rect 438584 152464 438636 152516
rect 453488 152464 453540 152516
rect 66628 152396 66680 152448
rect 159364 152396 159416 152448
rect 167000 152396 167052 152448
rect 175924 152396 175976 152448
rect 176108 152396 176160 152448
rect 249248 152396 249300 152448
rect 260840 152396 260892 152448
rect 316040 152396 316092 152448
rect 317512 152396 317564 152448
rect 320824 152396 320876 152448
rect 325884 152396 325936 152448
rect 367376 152396 367428 152448
rect 371332 152396 371384 152448
rect 402060 152396 402112 152448
rect 404176 152396 404228 152448
rect 407948 152396 408000 152448
rect 410892 152396 410944 152448
rect 430948 152396 431000 152448
rect 434720 152396 434772 152448
rect 450912 152396 450964 152448
rect 33600 152328 33652 152380
rect 109684 152328 109736 152380
rect 109776 152328 109828 152380
rect 110512 152328 110564 152380
rect 120080 152328 120132 152380
rect 210792 152328 210844 152380
rect 224040 152328 224092 152380
rect 287796 152328 287848 152380
rect 292212 152328 292264 152380
rect 341708 152328 341760 152380
rect 343824 152328 343876 152380
rect 349804 152328 349856 152380
rect 349896 152328 349948 152380
rect 385408 152328 385460 152380
rect 388352 152328 388404 152380
rect 392032 152328 392084 152380
rect 394608 152328 394660 152380
rect 417516 152328 417568 152380
rect 417608 152328 417660 152380
rect 418896 152328 418948 152380
rect 426900 152328 426952 152380
rect 431592 152328 431644 152380
rect 431868 152328 431920 152380
rect 432512 152328 432564 152380
rect 432604 152328 432656 152380
rect 441896 152328 441948 152380
rect 445300 152328 445352 152380
rect 458548 152328 458600 152380
rect 9496 152260 9548 152312
rect 82820 152260 82872 152312
rect 91100 152260 91152 152312
rect 179972 152260 180024 152312
rect 187884 152260 187936 152312
rect 262220 152260 262272 152312
rect 266360 152260 266412 152312
rect 320548 152260 320600 152312
rect 320824 152260 320876 152312
rect 325700 152260 325752 152312
rect 331220 152260 331272 152312
rect 371884 152260 371936 152312
rect 381084 152260 381136 152312
rect 409880 152260 409932 152312
rect 19800 152192 19852 152244
rect 97908 152192 97960 152244
rect 109040 152192 109092 152244
rect 130568 152192 130620 152244
rect 134064 152192 134116 152244
rect 221004 152192 221056 152244
rect 222108 152192 222160 152244
rect 282920 152192 282972 152244
rect 285772 152192 285824 152244
rect 335912 152192 335964 152244
rect 349160 152192 349212 152244
rect 349896 152192 349948 152244
rect 352012 152192 352064 152244
rect 387984 152192 388036 152244
rect 388444 152192 388496 152244
rect 407212 152192 407264 152244
rect 409236 152192 409288 152244
rect 412916 152260 412968 152312
rect 420920 152260 420972 152312
rect 422300 152260 422352 152312
rect 424048 152260 424100 152312
rect 425152 152260 425204 152312
rect 432420 152260 432472 152312
rect 428372 152192 428424 152244
rect 435548 152260 435600 152312
rect 436100 152260 436152 152312
rect 446496 152260 446548 152312
rect 82912 152124 82964 152176
rect 169760 152124 169812 152176
rect 172704 152124 172756 152176
rect 176108 152124 176160 152176
rect 176200 152124 176252 152176
rect 190184 152124 190236 152176
rect 193404 152124 193456 152176
rect 213276 152124 213328 152176
rect 244372 152124 244424 152176
rect 305736 152124 305788 152176
rect 320732 152124 320784 152176
rect 356520 152124 356572 152176
rect 357532 152124 357584 152176
rect 359096 152124 359148 152176
rect 365720 152124 365772 152176
rect 398196 152124 398248 152176
rect 405464 152124 405516 152176
rect 412732 152124 412784 152176
rect 78772 152056 78824 152108
rect 164516 152056 164568 152108
rect 169852 152056 169904 152108
rect 68928 151988 68980 152040
rect 142804 151988 142856 152040
rect 143356 151988 143408 152040
rect 146668 151988 146720 152040
rect 156420 151988 156472 152040
rect 172520 151988 172572 152040
rect 175924 152056 175976 152108
rect 182456 152056 182508 152108
rect 182548 152056 182600 152108
rect 185032 151988 185084 152040
rect 191656 152056 191708 152108
rect 208400 152056 208452 152108
rect 213644 152056 213696 152108
rect 274272 152056 274324 152108
rect 277400 152056 277452 152108
rect 330852 152056 330904 152108
rect 335360 152056 335412 152108
rect 375380 152056 375432 152108
rect 384948 152056 385000 152108
rect 391940 152056 391992 152108
rect 392032 152056 392084 152108
rect 404636 152056 404688 152108
rect 413008 152124 413060 152176
rect 413928 152124 413980 152176
rect 416228 152124 416280 152176
rect 416596 152124 416648 152176
rect 426532 152124 426584 152176
rect 200488 151988 200540 152040
rect 212632 151988 212684 152040
rect 272432 151988 272484 152040
rect 272524 151988 272576 152040
rect 320824 151988 320876 152040
rect 321560 151988 321612 152040
rect 362316 151988 362368 152040
rect 378600 151988 378652 152040
rect 384120 151988 384172 152040
rect 386328 151988 386380 152040
rect 399484 151988 399536 152040
rect 75092 151920 75144 151972
rect 154212 151920 154264 151972
rect 162584 151920 162636 151972
rect 177396 151920 177448 151972
rect 184664 151920 184716 151972
rect 195336 151920 195388 151972
rect 241612 151920 241664 151972
rect 300860 151920 300912 151972
rect 304080 151920 304132 151972
rect 351368 151920 351420 151972
rect 354680 151920 354732 151972
rect 389916 151920 389968 151972
rect 398932 151920 398984 151972
rect 30196 151852 30248 151904
rect 110328 151852 110380 151904
rect 110512 151852 110564 151904
rect 138296 151852 138348 151904
rect 139308 151852 139360 151904
rect 203064 151852 203116 151904
rect 243360 151852 243412 151904
rect 302608 151852 302660 151904
rect 307392 151852 307444 151904
rect 352012 151852 352064 151904
rect 363236 151852 363288 151904
rect 364340 151852 364392 151904
rect 385132 151852 385184 151904
rect 394700 151852 394752 151904
rect 396264 151852 396316 151904
rect 402980 151852 403032 151904
rect 404268 151852 404320 151904
rect 413560 151988 413612 152040
rect 408592 151920 408644 151972
rect 423312 152056 423364 152108
rect 425980 152056 426032 152108
rect 419724 151988 419776 152040
rect 427084 151988 427136 152040
rect 428004 152124 428056 152176
rect 433064 152192 433116 152244
rect 436192 152192 436244 152244
rect 436284 152192 436336 152244
rect 447692 152192 447744 152244
rect 429292 152124 429344 152176
rect 427452 152056 427504 152108
rect 432420 152056 432472 152108
rect 432972 152124 433024 152176
rect 443828 152124 443880 152176
rect 443920 152124 443972 152176
rect 457352 152260 457404 152312
rect 447876 152124 447928 152176
rect 456064 152124 456116 152176
rect 446312 152056 446364 152108
rect 446404 152056 446456 152108
rect 449900 152056 449952 152108
rect 515772 152056 515824 152108
rect 518992 152056 519044 152108
rect 432328 151988 432380 152040
rect 432880 151988 432932 152040
rect 443184 151988 443236 152040
rect 444472 151988 444524 152040
rect 458180 151988 458232 152040
rect 459560 151988 459612 152040
rect 461768 151988 461820 152040
rect 485780 151988 485832 152040
rect 490012 151988 490064 152040
rect 516048 151988 516100 152040
rect 520188 151988 520240 152040
rect 413836 151920 413888 151972
rect 421380 151920 421432 151972
rect 422760 151920 422812 151972
rect 432604 151920 432656 151972
rect 432696 151920 432748 151972
rect 435456 151920 435508 151972
rect 435548 151920 435600 151972
rect 439320 151920 439372 151972
rect 440240 151920 440292 151972
rect 454776 151920 454828 151972
rect 469220 151920 469272 151972
rect 472072 151920 472124 151972
rect 487344 151920 487396 151972
rect 490656 151920 490708 151972
rect 509148 151920 509200 151972
rect 510896 151920 510948 151972
rect 517428 151920 517480 151972
rect 521568 151920 521620 151972
rect 407948 151852 408000 151904
rect 415676 151852 415728 151904
rect 74816 151784 74868 151836
rect 81348 151784 81400 151836
rect 105820 151784 105872 151836
rect 110236 151784 110288 151836
rect 110420 151784 110472 151836
rect 127900 151784 127952 151836
rect 129740 151784 129792 151836
rect 146576 151784 146628 151836
rect 146668 151784 146720 151836
rect 156788 151784 156840 151836
rect 172428 151784 172480 151836
rect 176200 151784 176252 151836
rect 283196 151784 283248 151836
rect 287152 151784 287204 151836
rect 299664 151784 299716 151836
rect 81716 151716 81768 151768
rect 112812 151716 112864 151768
rect 346400 151784 346452 151836
rect 349804 151784 349856 151836
rect 380256 151784 380308 151836
rect 398104 151784 398156 151836
rect 407856 151784 407908 151836
rect 413560 151784 413612 151836
rect 418160 151852 418212 151904
rect 419632 151852 419684 151904
rect 436744 151852 436796 151904
rect 417424 151784 417476 151836
rect 423956 151784 424008 151836
rect 424048 151784 424100 151836
rect 441252 151852 441304 151904
rect 441804 151852 441856 151904
rect 446220 151852 446272 151904
rect 446496 151852 446548 151904
rect 451556 151852 451608 151904
rect 468024 151852 468076 151904
rect 470784 151852 470836 151904
rect 488172 151852 488224 151904
rect 488540 151852 488592 151904
rect 491944 151852 491996 151904
rect 507768 151852 507820 151904
rect 509516 151852 509568 151904
rect 437756 151784 437808 151836
rect 432420 151716 432472 151768
rect 434168 151716 434220 151768
rect 452844 151784 452896 151836
rect 467932 151784 467984 151836
rect 471428 151784 471480 151836
rect 491300 151784 491352 151836
rect 499120 151784 499172 151836
rect 499764 151784 499816 151836
rect 517060 151784 517112 151836
rect 520280 151784 520332 151836
rect 98920 151648 98972 151700
rect 116032 151648 116084 151700
rect 95516 151580 95568 151632
rect 115296 151580 115348 151632
rect 92020 151512 92072 151564
rect 113088 151512 113140 151564
rect 26700 151444 26752 151496
rect 116952 151444 117004 151496
rect 16396 151376 16448 151428
rect 116768 151376 116820 151428
rect 12992 151308 13044 151360
rect 116676 151308 116728 151360
rect 68008 151240 68060 151292
rect 112720 151240 112772 151292
rect 64512 151172 64564 151224
rect 112628 151172 112680 151224
rect 61108 151104 61160 151156
rect 112536 151104 112588 151156
rect 57704 151036 57756 151088
rect 110972 151036 111024 151088
rect 54208 150968 54260 151020
rect 112444 150968 112496 151020
rect 50804 150900 50856 150952
rect 111708 150900 111760 150952
rect 47308 150832 47360 150884
rect 111616 150832 111668 150884
rect 43904 150764 43956 150816
rect 111524 150764 111576 150816
rect 40500 150696 40552 150748
rect 111432 150696 111484 150748
rect 37004 150628 37056 150680
rect 111248 150628 111300 150680
rect 88616 150560 88668 150612
rect 112996 150560 113048 150612
rect 85212 150492 85264 150544
rect 115204 150492 115256 150544
rect 122840 150492 122892 150544
rect 123392 150492 123444 150544
rect 283104 150492 283156 150544
rect 283932 150492 283984 150544
rect 299480 150492 299532 150544
rect 300032 150492 300084 150544
rect 328460 150492 328512 150544
rect 328920 150492 328972 150544
rect 332692 150492 332744 150544
rect 333428 150492 333480 150544
rect 362960 150492 363012 150544
rect 363604 150492 363656 150544
rect 102324 150424 102376 150476
rect 116124 150424 116176 150476
rect 78312 150288 78364 150340
rect 112904 150288 112956 150340
rect 110328 150220 110380 150272
rect 117136 150220 117188 150272
rect 97908 150152 97960 150204
rect 116860 150152 116912 150204
rect 81348 150084 81400 150136
rect 92480 150084 92532 150136
rect 117228 150084 117280 150136
rect 116492 150016 116544 150068
rect 111156 148316 111208 148368
rect 117044 148316 117096 148368
rect 113088 140700 113140 140752
rect 116124 140700 116176 140752
rect 112996 137912 113048 137964
rect 116124 137912 116176 137964
rect 112812 133832 112864 133884
rect 116032 133832 116084 133884
rect 114192 132608 114244 132660
rect 115204 132608 115256 132660
rect 112904 132404 112956 132456
rect 116124 132404 116176 132456
rect 112720 126896 112772 126948
rect 116124 126896 116176 126948
rect 112628 124108 112680 124160
rect 116124 124108 116176 124160
rect 112536 122748 112588 122800
rect 115940 122748 115992 122800
rect 111708 121388 111760 121440
rect 116124 121388 116176 121440
rect 112444 118600 112496 118652
rect 116124 118600 116176 118652
rect 111616 117240 111668 117292
rect 116124 117240 116176 117292
rect 111524 114452 111576 114504
rect 116124 114452 116176 114504
rect 111432 113092 111484 113144
rect 115940 113092 115992 113144
rect 111340 111732 111392 111784
rect 116124 111732 116176 111784
rect 111156 108944 111208 108996
rect 116124 108944 116176 108996
rect 111248 92420 111300 92472
rect 116124 92420 116176 92472
rect 111064 89632 111116 89684
rect 116124 89632 116176 89684
rect 113824 88272 113876 88324
rect 116032 88272 116084 88324
rect 113916 83920 113968 83972
rect 116584 83920 116636 83972
rect 114008 82764 114060 82816
rect 116216 82764 116268 82816
rect 114100 79976 114152 80028
rect 115940 79976 115992 80028
rect 114192 78616 114244 78668
rect 116124 78616 116176 78668
rect 114192 71748 114244 71800
rect 116584 71748 116636 71800
rect 114100 69028 114152 69080
rect 116308 69028 116360 69080
rect 114008 67600 114060 67652
rect 116124 67600 116176 67652
rect 113916 66240 113968 66292
rect 116584 66240 116636 66292
rect 113364 64676 113416 64728
rect 116584 64676 116636 64728
rect 113824 63520 113876 63572
rect 116216 63520 116268 63572
rect 112444 62092 112496 62144
rect 116124 62092 116176 62144
rect 112536 42780 112588 42832
rect 116124 42780 116176 42832
rect 116400 7624 116452 7676
rect 116308 7420 116360 7472
rect 111064 2796 111116 2848
rect 143632 2456 143684 2508
rect 425796 2456 425848 2508
rect 443644 2456 443696 2508
rect 42064 1844 42116 1896
rect 44732 1844 44784 1896
rect 62396 1844 62448 1896
rect 68284 1844 68336 1896
rect 91928 1844 91980 1896
rect 99196 1844 99248 1896
rect 102600 1844 102652 1896
rect 102692 1844 102744 1896
rect 89352 1776 89404 1828
rect 105912 1844 105964 1896
rect 109132 1844 109184 1896
rect 109684 1844 109736 1896
rect 109776 1844 109828 1896
rect 109868 1844 109920 1896
rect 59360 1708 59412 1760
rect 78772 1708 78824 1760
rect 86040 1708 86092 1760
rect 109316 1776 109368 1828
rect 112444 1776 112496 1828
rect 82636 1640 82688 1692
rect 103980 1640 104032 1692
rect 109960 1708 110012 1760
rect 110052 1708 110104 1760
rect 116584 1708 116636 1760
rect 69296 1572 69348 1624
rect 103796 1572 103848 1624
rect 79324 1504 79376 1556
rect 105912 1572 105964 1624
rect 106004 1572 106056 1624
rect 109040 1572 109092 1624
rect 109224 1640 109276 1692
rect 110604 1640 110656 1692
rect 110144 1572 110196 1624
rect 103980 1504 104032 1556
rect 110236 1504 110288 1556
rect 46020 1436 46072 1488
rect 64052 1436 64104 1488
rect 72700 1436 72752 1488
rect 109592 1436 109644 1488
rect 193588 1436 193640 1488
rect 32680 1368 32732 1420
rect 109132 1368 109184 1420
rect 109224 1368 109276 1420
rect 110052 1368 110104 1420
rect 2688 1300 2740 1352
rect 35992 1232 36044 1284
rect 109408 1300 109460 1352
rect 116400 1368 116452 1420
rect 294788 1368 294840 1420
rect 343640 1368 343692 1420
rect 491300 1368 491352 1420
rect 493600 1368 493652 1420
rect 39304 1164 39356 1216
rect 109040 1164 109092 1216
rect 116308 1232 116360 1284
rect 116492 1164 116544 1216
rect 49332 1096 49384 1148
rect 117044 1096 117096 1148
rect 52644 1028 52696 1080
rect 65984 960 66036 1012
rect 97264 960 97316 1012
rect 76012 892 76064 944
rect 116860 960 116912 1012
rect 112536 892 112588 944
rect 91560 824 91612 876
rect 93860 824 93912 876
rect 97264 824 97316 876
rect 116676 824 116728 876
rect 109040 756 109092 808
rect 117228 756 117280 808
rect 103796 688 103848 740
rect 110788 688 110840 740
<< metal2 >>
rect 386 163200 442 164400
rect 492 163254 1164 163282
rect 400 158030 428 163200
rect 388 158024 440 158030
rect 388 157966 440 157972
rect 492 153882 520 163254
rect 1136 163146 1164 163254
rect 1214 163200 1270 164400
rect 2042 163200 2098 164400
rect 2870 163200 2926 164400
rect 2976 163254 3648 163282
rect 1228 163146 1256 163200
rect 1136 163118 1256 163146
rect 2056 156670 2084 163200
rect 2044 156664 2096 156670
rect 2044 156606 2096 156612
rect 480 153876 532 153882
rect 480 153818 532 153824
rect 2884 152522 2912 163200
rect 2976 153785 3004 163254
rect 3620 163146 3648 163254
rect 3698 163200 3754 164400
rect 4526 163200 4582 164400
rect 5354 163200 5410 164400
rect 6274 163200 6330 164400
rect 7102 163200 7158 164400
rect 7930 163200 7986 164400
rect 8758 163200 8814 164400
rect 8864 163254 9536 163282
rect 3712 163146 3740 163200
rect 3620 163118 3740 163146
rect 4540 155310 4568 163200
rect 4528 155304 4580 155310
rect 4528 155246 4580 155252
rect 5368 155242 5396 163200
rect 6288 159390 6316 163200
rect 6276 159384 6328 159390
rect 6276 159326 6328 159332
rect 5356 155236 5408 155242
rect 5356 155178 5408 155184
rect 7116 153950 7144 163200
rect 7944 155446 7972 163200
rect 7932 155440 7984 155446
rect 7932 155382 7984 155388
rect 8772 155378 8800 163200
rect 8760 155372 8812 155378
rect 8760 155314 8812 155320
rect 7104 153944 7156 153950
rect 7104 153886 7156 153892
rect 2962 153776 3018 153785
rect 2962 153711 3018 153720
rect 2872 152516 2924 152522
rect 2872 152458 2924 152464
rect 8864 152425 8892 163254
rect 9508 163146 9536 163254
rect 9586 163200 9642 164400
rect 9692 163254 10364 163282
rect 9600 163146 9628 163200
rect 9508 163118 9628 163146
rect 9692 154018 9720 163254
rect 10336 163146 10364 163254
rect 10414 163200 10470 164400
rect 11242 163200 11298 164400
rect 12162 163200 12218 164400
rect 12452 163254 12940 163282
rect 10428 163146 10456 163200
rect 10336 163118 10456 163146
rect 11256 156738 11284 163200
rect 11244 156732 11296 156738
rect 11244 156674 11296 156680
rect 12176 155786 12204 163200
rect 12164 155780 12216 155786
rect 12164 155722 12216 155728
rect 9680 154012 9732 154018
rect 9680 153954 9732 153960
rect 12452 152561 12480 163254
rect 12912 163146 12940 163254
rect 12990 163200 13046 164400
rect 13818 163200 13874 164400
rect 14646 163200 14702 164400
rect 15474 163200 15530 164400
rect 16302 163200 16358 164400
rect 16592 163254 17080 163282
rect 13004 163146 13032 163200
rect 12912 163118 13032 163146
rect 13832 154086 13860 163200
rect 14660 156806 14688 163200
rect 14648 156800 14700 156806
rect 14648 156742 14700 156748
rect 15488 154970 15516 163200
rect 16316 159361 16344 163200
rect 16302 159352 16358 159361
rect 16302 159287 16358 159296
rect 15476 154964 15528 154970
rect 15476 154906 15528 154912
rect 13820 154080 13872 154086
rect 13820 154022 13872 154028
rect 16592 153921 16620 163254
rect 17052 163146 17080 163254
rect 17130 163200 17186 164400
rect 18050 163200 18106 164400
rect 18878 163200 18934 164400
rect 19352 163254 19656 163282
rect 17144 163146 17172 163200
rect 17052 163118 17172 163146
rect 18064 156942 18092 163200
rect 18892 159730 18920 163200
rect 18880 159724 18932 159730
rect 18880 159666 18932 159672
rect 18052 156936 18104 156942
rect 18052 156878 18104 156884
rect 16578 153912 16634 153921
rect 16578 153847 16634 153856
rect 19352 152590 19380 163254
rect 19628 163146 19656 163254
rect 19706 163200 19762 164400
rect 19904 163254 20484 163282
rect 19720 163146 19748 163200
rect 19628 163118 19748 163146
rect 19904 154057 19932 163254
rect 20456 163146 20484 163254
rect 20534 163200 20590 164400
rect 21362 163200 21418 164400
rect 22190 163200 22246 164400
rect 23018 163200 23074 164400
rect 23492 163254 23888 163282
rect 20548 163146 20576 163200
rect 20456 163118 20576 163146
rect 21376 156874 21404 163200
rect 21364 156868 21416 156874
rect 21364 156810 21416 156816
rect 19890 154048 19946 154057
rect 19890 153983 19946 153992
rect 22204 152658 22232 163200
rect 23032 159497 23060 163200
rect 23018 159488 23074 159497
rect 23018 159423 23074 159432
rect 23492 154154 23520 163254
rect 23860 163146 23888 163254
rect 23938 163200 23994 164400
rect 24766 163200 24822 164400
rect 25594 163200 25650 164400
rect 26422 163200 26478 164400
rect 27250 163200 27306 164400
rect 28078 163200 28134 164400
rect 28184 163254 28856 163282
rect 23952 163146 23980 163200
rect 23860 163118 23980 163146
rect 24780 157010 24808 163200
rect 25608 160002 25636 163200
rect 25596 159996 25648 160002
rect 25596 159938 25648 159944
rect 24768 157004 24820 157010
rect 24768 156946 24820 156952
rect 23480 154148 23532 154154
rect 23480 154090 23532 154096
rect 23296 153196 23348 153202
rect 23296 153138 23348 153144
rect 22192 152652 22244 152658
rect 22192 152594 22244 152600
rect 19340 152584 19392 152590
rect 12438 152552 12494 152561
rect 19340 152526 19392 152532
rect 12438 152487 12494 152496
rect 8850 152416 8906 152425
rect 8850 152351 8906 152360
rect 9496 152312 9548 152318
rect 9496 152254 9548 152260
rect 6090 150648 6146 150657
rect 6090 150583 6146 150592
rect 2686 150512 2742 150521
rect 2686 150447 2742 150456
rect 2700 149940 2728 150447
rect 6104 149940 6132 150583
rect 9508 149940 9536 152254
rect 19800 152244 19852 152250
rect 19800 152186 19852 152192
rect 16396 151428 16448 151434
rect 16396 151370 16448 151376
rect 12992 151360 13044 151366
rect 12992 151302 13044 151308
rect 13004 149940 13032 151302
rect 16408 149940 16436 151370
rect 19812 149940 19840 152186
rect 23308 149940 23336 153138
rect 26436 152794 26464 163200
rect 27264 154222 27292 163200
rect 28092 156641 28120 163200
rect 28078 156632 28134 156641
rect 28078 156567 28134 156576
rect 27252 154216 27304 154222
rect 27252 154158 27304 154164
rect 26424 152788 26476 152794
rect 26424 152730 26476 152736
rect 28184 152726 28212 163254
rect 28828 163146 28856 163254
rect 28906 163200 28962 164400
rect 29826 163200 29882 164400
rect 30392 163254 30604 163282
rect 28920 163146 28948 163200
rect 28828 163118 28948 163146
rect 29840 159633 29868 163200
rect 29826 159624 29882 159633
rect 29826 159559 29882 159568
rect 30392 154193 30420 163254
rect 30576 163146 30604 163254
rect 30654 163200 30710 164400
rect 31482 163200 31538 164400
rect 32310 163200 32366 164400
rect 33138 163200 33194 164400
rect 33966 163200 34022 164400
rect 34532 163254 34744 163282
rect 30668 163146 30696 163200
rect 30576 163118 30696 163146
rect 31496 156777 31524 163200
rect 32324 159458 32352 163200
rect 32312 159452 32364 159458
rect 32312 159394 32364 159400
rect 31482 156768 31538 156777
rect 31482 156703 31538 156712
rect 30378 154184 30434 154193
rect 30378 154119 30434 154128
rect 33152 152862 33180 163200
rect 33980 158001 34008 163200
rect 33966 157992 34022 158001
rect 33966 157927 34022 157936
rect 34532 154358 34560 163254
rect 34716 163146 34744 163254
rect 34794 163200 34850 164400
rect 35714 163200 35770 164400
rect 36542 163200 36598 164400
rect 37370 163200 37426 164400
rect 37936 163254 38148 163282
rect 34808 163146 34836 163200
rect 34716 163118 34836 163146
rect 35728 157078 35756 163200
rect 36556 159526 36584 163200
rect 36544 159520 36596 159526
rect 36544 159462 36596 159468
rect 37384 158098 37412 163200
rect 37372 158092 37424 158098
rect 37372 158034 37424 158040
rect 35716 157072 35768 157078
rect 35716 157014 35768 157020
rect 34520 154352 34572 154358
rect 34520 154294 34572 154300
rect 37936 154290 37964 163254
rect 38120 163146 38148 163254
rect 38198 163200 38254 164400
rect 39026 163200 39082 164400
rect 39854 163200 39910 164400
rect 40682 163200 40738 164400
rect 41602 163200 41658 164400
rect 42430 163200 42486 164400
rect 43258 163200 43314 164400
rect 44086 163200 44142 164400
rect 44192 163254 44864 163282
rect 38212 163146 38240 163200
rect 38120 163118 38240 163146
rect 39040 157214 39068 163200
rect 39028 157208 39080 157214
rect 39028 157150 39080 157156
rect 39868 155582 39896 163200
rect 40696 158273 40724 163200
rect 40682 158264 40738 158273
rect 40682 158199 40738 158208
rect 39856 155576 39908 155582
rect 39856 155518 39908 155524
rect 37924 154284 37976 154290
rect 37924 154226 37976 154232
rect 41616 153270 41644 163200
rect 42444 157146 42472 163200
rect 43272 159594 43300 163200
rect 43260 159588 43312 159594
rect 43260 159530 43312 159536
rect 44100 158137 44128 163200
rect 44086 158128 44142 158137
rect 44086 158063 44142 158072
rect 42432 157140 42484 157146
rect 42432 157082 42484 157088
rect 44192 154494 44220 163254
rect 44836 163146 44864 163254
rect 44914 163200 44970 164400
rect 45742 163200 45798 164400
rect 46570 163200 46626 164400
rect 47490 163200 47546 164400
rect 48318 163200 48374 164400
rect 49146 163200 49202 164400
rect 49974 163200 50030 164400
rect 50802 163200 50858 164400
rect 51092 163254 51580 163282
rect 44928 163146 44956 163200
rect 44836 163118 44956 163146
rect 45756 157282 45784 163200
rect 45744 157276 45796 157282
rect 45744 157218 45796 157224
rect 46584 155718 46612 163200
rect 47504 158166 47532 163200
rect 47492 158160 47544 158166
rect 47492 158102 47544 158108
rect 46572 155712 46624 155718
rect 46572 155654 46624 155660
rect 44180 154488 44232 154494
rect 44180 154430 44232 154436
rect 48332 153814 48360 163200
rect 49160 157350 49188 163200
rect 49988 159662 50016 163200
rect 49976 159656 50028 159662
rect 49976 159598 50028 159604
rect 50816 158234 50844 163200
rect 50804 158228 50856 158234
rect 50804 158170 50856 158176
rect 49148 157344 49200 157350
rect 49148 157286 49200 157292
rect 51092 154562 51120 163254
rect 51552 163146 51580 163254
rect 51630 163200 51686 164400
rect 52458 163200 52514 164400
rect 53378 163200 53434 164400
rect 54206 163200 54262 164400
rect 54312 163254 54984 163282
rect 51644 163146 51672 163200
rect 51552 163118 51672 163146
rect 52472 156602 52500 163200
rect 52460 156596 52512 156602
rect 52460 156538 52512 156544
rect 53392 155650 53420 163200
rect 54220 158302 54248 163200
rect 54208 158296 54260 158302
rect 54208 158238 54260 158244
rect 53380 155644 53432 155650
rect 53380 155586 53432 155592
rect 51080 154556 51132 154562
rect 51080 154498 51132 154504
rect 54312 154329 54340 163254
rect 54956 163146 54984 163254
rect 55034 163200 55090 164400
rect 55862 163200 55918 164400
rect 56690 163200 56746 164400
rect 57518 163200 57574 164400
rect 57992 163254 58296 163282
rect 55048 163146 55076 163200
rect 54956 163118 55076 163146
rect 55876 156913 55904 163200
rect 56704 159798 56732 163200
rect 56692 159792 56744 159798
rect 56692 159734 56744 159740
rect 57532 158409 57560 163200
rect 57518 158400 57574 158409
rect 57518 158335 57574 158344
rect 55862 156904 55918 156913
rect 55862 156839 55918 156848
rect 54298 154320 54354 154329
rect 54298 154255 54354 154264
rect 48320 153808 48372 153814
rect 48320 153750 48372 153756
rect 57992 153678 58020 163254
rect 58268 163146 58296 163254
rect 58346 163200 58402 164400
rect 59266 163200 59322 164400
rect 60094 163200 60150 164400
rect 60922 163200 60978 164400
rect 61120 163254 61700 163282
rect 58360 163146 58388 163200
rect 58268 163118 58388 163146
rect 59280 156534 59308 163200
rect 59268 156528 59320 156534
rect 59268 156470 59320 156476
rect 60108 155854 60136 163200
rect 60936 158438 60964 163200
rect 60924 158432 60976 158438
rect 60924 158374 60976 158380
rect 60096 155848 60148 155854
rect 60096 155790 60148 155796
rect 61120 153746 61148 163254
rect 61672 163146 61700 163254
rect 61750 163200 61806 164400
rect 62578 163200 62634 164400
rect 63406 163200 63462 164400
rect 64234 163200 64290 164400
rect 65154 163200 65210 164400
rect 65982 163200 66038 164400
rect 66810 163200 66866 164400
rect 67638 163200 67694 164400
rect 68466 163200 68522 164400
rect 69294 163200 69350 164400
rect 70122 163200 70178 164400
rect 71042 163200 71098 164400
rect 71870 163200 71926 164400
rect 72698 163200 72754 164400
rect 73526 163200 73582 164400
rect 74354 163200 74410 164400
rect 75182 163200 75238 164400
rect 76010 163200 76066 164400
rect 76930 163200 76986 164400
rect 77758 163200 77814 164400
rect 78586 163200 78642 164400
rect 78692 163254 79364 163282
rect 61764 163146 61792 163200
rect 61672 163118 61792 163146
rect 62592 155417 62620 163200
rect 63420 160070 63448 163200
rect 63408 160064 63460 160070
rect 63408 160006 63460 160012
rect 64248 158370 64276 163200
rect 64236 158364 64288 158370
rect 64236 158306 64288 158312
rect 65168 155514 65196 163200
rect 65996 155553 66024 163200
rect 66824 155922 66852 163200
rect 67652 158642 67680 163200
rect 67640 158636 67692 158642
rect 67640 158578 67692 158584
rect 66812 155916 66864 155922
rect 66812 155858 66864 155864
rect 66628 155644 66680 155650
rect 66628 155586 66680 155592
rect 65982 155544 66038 155553
rect 65156 155508 65208 155514
rect 65982 155479 66038 155488
rect 65156 155450 65208 155456
rect 62578 155408 62634 155417
rect 62578 155343 62634 155352
rect 61108 153740 61160 153746
rect 61108 153682 61160 153688
rect 57980 153672 58032 153678
rect 57980 153614 58032 153620
rect 41604 153264 41656 153270
rect 41604 153206 41656 153212
rect 33140 152856 33192 152862
rect 33140 152798 33192 152804
rect 28172 152720 28224 152726
rect 28172 152662 28224 152668
rect 66640 152454 66668 155586
rect 68480 155281 68508 163200
rect 69308 156466 69336 163200
rect 70136 159866 70164 163200
rect 70124 159860 70176 159866
rect 70124 159802 70176 159808
rect 71056 158506 71084 163200
rect 71044 158500 71096 158506
rect 71044 158442 71096 158448
rect 69296 156460 69348 156466
rect 69296 156402 69348 156408
rect 71884 155650 71912 163200
rect 72712 157049 72740 163200
rect 73540 159322 73568 163200
rect 73528 159316 73580 159322
rect 73528 159258 73580 159264
rect 74368 158574 74396 163200
rect 74356 158568 74408 158574
rect 74356 158510 74408 158516
rect 72698 157040 72754 157049
rect 72698 156975 72754 156984
rect 75092 155712 75144 155718
rect 75092 155654 75144 155660
rect 71872 155644 71924 155650
rect 71872 155586 71924 155592
rect 68928 155576 68980 155582
rect 68928 155518 68980 155524
rect 68466 155272 68522 155281
rect 68466 155207 68522 155216
rect 66628 152448 66680 152454
rect 66628 152390 66680 152396
rect 33600 152380 33652 152386
rect 33600 152322 33652 152328
rect 30196 151904 30248 151910
rect 30196 151846 30248 151852
rect 26700 151496 26752 151502
rect 26700 151438 26752 151444
rect 26712 149940 26740 151438
rect 30208 149940 30236 151846
rect 33612 149940 33640 152322
rect 68940 152046 68968 155518
rect 71412 152924 71464 152930
rect 71412 152866 71464 152872
rect 68928 152040 68980 152046
rect 68928 151982 68980 151988
rect 68008 151292 68060 151298
rect 68008 151234 68060 151240
rect 64512 151224 64564 151230
rect 64512 151166 64564 151172
rect 61108 151156 61160 151162
rect 61108 151098 61160 151104
rect 57704 151088 57756 151094
rect 57704 151030 57756 151036
rect 54208 151020 54260 151026
rect 54208 150962 54260 150968
rect 50804 150952 50856 150958
rect 50804 150894 50856 150900
rect 47308 150884 47360 150890
rect 47308 150826 47360 150832
rect 43904 150816 43956 150822
rect 43904 150758 43956 150764
rect 40500 150748 40552 150754
rect 40500 150690 40552 150696
rect 37004 150680 37056 150686
rect 37004 150622 37056 150628
rect 37016 149940 37044 150622
rect 40512 149940 40540 150690
rect 43916 149940 43944 150758
rect 47320 149940 47348 150826
rect 50816 149940 50844 150894
rect 54220 149940 54248 150962
rect 57716 149940 57744 151030
rect 61120 149940 61148 151098
rect 64524 149940 64552 151166
rect 68020 149940 68048 151234
rect 71424 149940 71452 152866
rect 75104 151978 75132 155654
rect 75196 155582 75224 163200
rect 76024 155825 76052 163200
rect 76944 159934 76972 163200
rect 76932 159928 76984 159934
rect 76932 159870 76984 159876
rect 77772 157962 77800 163200
rect 77760 157956 77812 157962
rect 77760 157898 77812 157904
rect 76010 155816 76066 155825
rect 76010 155751 76066 155760
rect 78600 155689 78628 163200
rect 78586 155680 78642 155689
rect 78586 155615 78642 155624
rect 75184 155576 75236 155582
rect 75184 155518 75236 155524
rect 78692 153610 78720 163254
rect 79336 163146 79364 163254
rect 79414 163200 79470 164400
rect 80242 163200 80298 164400
rect 81070 163200 81126 164400
rect 81898 163200 81954 164400
rect 82818 163200 82874 164400
rect 83646 163200 83702 164400
rect 84474 163200 84530 164400
rect 85302 163200 85358 164400
rect 85592 163254 86080 163282
rect 79428 163146 79456 163200
rect 79336 163118 79456 163146
rect 80060 159316 80112 159322
rect 80060 159258 80112 159264
rect 78772 155848 78824 155854
rect 78772 155790 78824 155796
rect 78680 153604 78732 153610
rect 78680 153546 78732 153552
rect 78784 152114 78812 155790
rect 80072 153134 80100 159258
rect 80256 159254 80284 163200
rect 80244 159248 80296 159254
rect 80244 159190 80296 159196
rect 81084 158710 81112 163200
rect 81072 158704 81124 158710
rect 81072 158646 81124 158652
rect 81912 155718 81940 163200
rect 82832 156398 82860 163200
rect 83660 159322 83688 163200
rect 83648 159316 83700 159322
rect 83648 159258 83700 159264
rect 84488 157894 84516 163200
rect 84476 157888 84528 157894
rect 84476 157830 84528 157836
rect 82820 156392 82872 156398
rect 82820 156334 82872 156340
rect 85316 155961 85344 163200
rect 85302 155952 85358 155961
rect 82912 155916 82964 155922
rect 85302 155887 85358 155896
rect 82912 155858 82964 155864
rect 81900 155712 81952 155718
rect 81900 155654 81952 155660
rect 80060 153128 80112 153134
rect 80060 153070 80112 153076
rect 82820 152312 82872 152318
rect 82820 152254 82872 152260
rect 78772 152108 78824 152114
rect 78772 152050 78824 152056
rect 75092 151972 75144 151978
rect 75092 151914 75144 151920
rect 74816 151836 74868 151842
rect 81348 151836 81400 151842
rect 74868 151786 74948 151814
rect 74816 151778 74868 151784
rect 74920 149954 74948 151786
rect 81348 151778 81400 151784
rect 78312 150340 78364 150346
rect 78312 150282 78364 150288
rect 74842 149926 74948 149954
rect 78324 149940 78352 150282
rect 81360 150142 81388 151778
rect 81716 151768 81768 151774
rect 81716 151710 81768 151716
rect 81348 150136 81400 150142
rect 81348 150078 81400 150084
rect 81728 149940 81756 151710
rect 82832 149705 82860 152254
rect 82924 152182 82952 155858
rect 85592 154465 85620 163254
rect 86052 163146 86080 163254
rect 86130 163200 86186 164400
rect 86958 163200 87014 164400
rect 87786 163200 87842 164400
rect 88706 163200 88762 164400
rect 89534 163200 89590 164400
rect 90362 163200 90418 164400
rect 91190 163200 91246 164400
rect 92018 163200 92074 164400
rect 92846 163200 92902 164400
rect 93674 163200 93730 164400
rect 94594 163200 94650 164400
rect 95422 163200 95478 164400
rect 96250 163200 96306 164400
rect 96632 163254 97028 163282
rect 86144 163146 86172 163200
rect 86052 163118 86172 163146
rect 86972 159186 87000 163200
rect 86960 159180 87012 159186
rect 86960 159122 87012 159128
rect 87800 157826 87828 163200
rect 87788 157820 87840 157826
rect 87788 157762 87840 157768
rect 88720 155854 88748 163200
rect 88708 155848 88760 155854
rect 88708 155790 88760 155796
rect 89548 155174 89576 163200
rect 90376 158778 90404 163200
rect 91100 159248 91152 159254
rect 91100 159190 91152 159196
rect 90364 158772 90416 158778
rect 90364 158714 90416 158720
rect 89536 155168 89588 155174
rect 89536 155110 89588 155116
rect 85578 154456 85634 154465
rect 85578 154391 85634 154400
rect 91112 152318 91140 159190
rect 91204 157758 91232 163200
rect 91192 157752 91244 157758
rect 91192 157694 91244 157700
rect 92032 155922 92060 163200
rect 92860 158778 92888 163200
rect 93688 159118 93716 163200
rect 93676 159112 93728 159118
rect 93676 159054 93728 159060
rect 92572 158772 92624 158778
rect 92572 158714 92624 158720
rect 92848 158772 92900 158778
rect 92848 158714 92900 158720
rect 92020 155916 92072 155922
rect 92020 155858 92072 155864
rect 92584 152998 92612 158714
rect 94608 157690 94636 163200
rect 94596 157684 94648 157690
rect 94596 157626 94648 157632
rect 95436 155106 95464 163200
rect 96264 158982 96292 163200
rect 96252 158976 96304 158982
rect 96252 158918 96304 158924
rect 95424 155100 95476 155106
rect 95424 155042 95476 155048
rect 92572 152992 92624 152998
rect 92572 152934 92624 152940
rect 96632 152930 96660 163254
rect 97000 163146 97028 163254
rect 97078 163200 97134 164400
rect 97906 163200 97962 164400
rect 98734 163200 98790 164400
rect 99562 163200 99618 164400
rect 100482 163200 100538 164400
rect 101310 163200 101366 164400
rect 102138 163200 102194 164400
rect 102966 163200 103022 164400
rect 103532 163254 103744 163282
rect 97092 163146 97120 163200
rect 97000 163118 97120 163146
rect 97920 157622 97948 163200
rect 97908 157616 97960 157622
rect 97908 157558 97960 157564
rect 98748 155038 98776 163200
rect 99576 156262 99604 163200
rect 100496 159254 100524 163200
rect 100484 159248 100536 159254
rect 100484 159190 100536 159196
rect 101324 156330 101352 163200
rect 101312 156324 101364 156330
rect 101312 156266 101364 156272
rect 99564 156256 99616 156262
rect 99564 156198 99616 156204
rect 98736 155032 98788 155038
rect 98736 154974 98788 154980
rect 102152 153542 102180 163200
rect 102980 158914 103008 163200
rect 102968 158908 103020 158914
rect 102968 158850 103020 158856
rect 102140 153536 102192 153542
rect 102140 153478 102192 153484
rect 103532 153066 103560 163254
rect 103716 163146 103744 163254
rect 103794 163200 103850 164400
rect 104622 163200 104678 164400
rect 104912 163254 105400 163282
rect 103808 163146 103836 163200
rect 103716 163118 103836 163146
rect 104636 158545 104664 163200
rect 104622 158536 104678 158545
rect 104622 158471 104678 158480
rect 104912 153474 104940 163254
rect 105372 163146 105400 163254
rect 105450 163200 105506 164400
rect 106370 163200 106426 164400
rect 107198 163200 107254 164400
rect 108026 163200 108082 164400
rect 108316 163254 108804 163282
rect 105464 163146 105492 163200
rect 105372 163118 105492 163146
rect 106384 154902 106412 163200
rect 107212 159050 107240 163200
rect 107200 159044 107252 159050
rect 107200 158986 107252 158992
rect 108040 156194 108068 163200
rect 108028 156188 108080 156194
rect 108028 156130 108080 156136
rect 106372 154896 106424 154902
rect 106372 154838 106424 154844
rect 104900 153468 104952 153474
rect 104900 153410 104952 153416
rect 108316 153406 108344 163254
rect 108776 163146 108804 163254
rect 108854 163200 108910 164400
rect 109682 163200 109738 164400
rect 110510 163200 110566 164400
rect 111338 163200 111394 164400
rect 112258 163200 112314 164400
rect 113086 163200 113142 164400
rect 113192 163254 113864 163282
rect 108868 163146 108896 163200
rect 108776 163118 108896 163146
rect 109132 159724 109184 159730
rect 109132 159666 109184 159672
rect 109040 154964 109092 154970
rect 109040 154906 109092 154912
rect 108304 153400 108356 153406
rect 108304 153342 108356 153348
rect 103520 153060 103572 153066
rect 103520 153002 103572 153008
rect 92480 152924 92532 152930
rect 92480 152866 92532 152872
rect 96620 152924 96672 152930
rect 96620 152866 96672 152872
rect 91100 152312 91152 152318
rect 91100 152254 91152 152260
rect 82912 152176 82964 152182
rect 82912 152118 82964 152124
rect 92020 151564 92072 151570
rect 92020 151506 92072 151512
rect 88616 150612 88668 150618
rect 88616 150554 88668 150560
rect 85212 150544 85264 150550
rect 85212 150486 85264 150492
rect 85224 149940 85252 150486
rect 88628 149940 88656 150554
rect 92032 149940 92060 151506
rect 92492 150142 92520 152866
rect 109052 152250 109080 154906
rect 109144 154766 109172 159666
rect 109696 158846 109724 163200
rect 109776 159996 109828 160002
rect 109776 159938 109828 159944
rect 109684 158840 109736 158846
rect 109684 158782 109736 158788
rect 109132 154760 109184 154766
rect 109132 154702 109184 154708
rect 109788 152386 109816 159938
rect 110328 155780 110380 155786
rect 110328 155722 110380 155728
rect 109684 152380 109736 152386
rect 109684 152322 109736 152328
rect 109776 152380 109828 152386
rect 109776 152322 109828 152328
rect 97908 152244 97960 152250
rect 97908 152186 97960 152192
rect 109040 152244 109092 152250
rect 109040 152186 109092 152192
rect 95516 151632 95568 151638
rect 95516 151574 95568 151580
rect 92480 150136 92532 150142
rect 92480 150078 92532 150084
rect 95528 149940 95556 151574
rect 97920 150210 97948 152186
rect 105820 151836 105872 151842
rect 105740 151786 105820 151814
rect 98920 151700 98972 151706
rect 98920 151642 98972 151648
rect 97908 150204 97960 150210
rect 97908 150146 97960 150152
rect 98932 149940 98960 151642
rect 102324 150476 102376 150482
rect 102324 150418 102376 150424
rect 102336 149940 102364 150418
rect 105740 149954 105768 151786
rect 105820 151778 105872 151784
rect 105740 149926 105846 149954
rect 82818 149696 82874 149705
rect 82818 149631 82874 149640
rect 109250 149382 109632 149410
rect 109604 148073 109632 149382
rect 109590 148064 109646 148073
rect 109590 147999 109646 148008
rect 109696 132494 109724 152322
rect 110340 151994 110368 155722
rect 110524 154834 110552 163200
rect 111352 157554 111380 163200
rect 111340 157548 111392 157554
rect 111340 157490 111392 157496
rect 112272 155786 112300 163200
rect 113100 159730 113128 163200
rect 113088 159724 113140 159730
rect 113088 159666 113140 159672
rect 112260 155780 112312 155786
rect 112260 155722 112312 155728
rect 110512 154828 110564 154834
rect 110512 154770 110564 154776
rect 113192 153202 113220 163254
rect 113836 163146 113864 163254
rect 113914 163200 113970 164400
rect 114742 163200 114798 164400
rect 115570 163200 115626 164400
rect 115952 163254 116348 163282
rect 113928 163146 113956 163200
rect 113836 163118 113956 163146
rect 114468 158772 114520 158778
rect 114468 158714 114520 158720
rect 114480 154426 114508 158714
rect 114756 157486 114784 163200
rect 114744 157480 114796 157486
rect 114744 157422 114796 157428
rect 115584 157185 115612 163200
rect 115570 157176 115626 157185
rect 115570 157111 115626 157120
rect 114468 154420 114520 154426
rect 114468 154362 114520 154368
rect 115952 153338 115980 163254
rect 116320 163146 116348 163254
rect 116398 163200 116454 164400
rect 117226 163200 117282 164400
rect 118146 163200 118202 164400
rect 118712 163254 118924 163282
rect 116412 163146 116440 163200
rect 116320 163118 116440 163146
rect 117240 160002 117268 163200
rect 117228 159996 117280 160002
rect 117228 159938 117280 159944
rect 118160 156126 118188 163200
rect 118148 156120 118200 156126
rect 118148 156062 118200 156068
rect 118608 154624 118660 154630
rect 118608 154566 118660 154572
rect 118620 154426 118648 154566
rect 118712 154426 118740 163254
rect 118896 163146 118924 163254
rect 118974 163200 119030 164400
rect 119802 163200 119858 164400
rect 120092 163254 120580 163282
rect 118988 163146 119016 163200
rect 118896 163118 119016 163146
rect 119816 158778 119844 163200
rect 119804 158772 119856 158778
rect 119804 158714 119856 158720
rect 118884 158024 118936 158030
rect 118884 157966 118936 157972
rect 118608 154420 118660 154426
rect 118608 154362 118660 154368
rect 118700 154420 118752 154426
rect 118700 154362 118752 154368
rect 115940 153332 115992 153338
rect 115940 153274 115992 153280
rect 110972 153196 111024 153202
rect 110972 153138 111024 153144
rect 113180 153196 113232 153202
rect 113180 153138 113232 153144
rect 110512 152380 110564 152386
rect 110512 152322 110564 152328
rect 110340 151966 110460 151994
rect 110328 151904 110380 151910
rect 110328 151846 110380 151852
rect 110236 151836 110288 151842
rect 110236 151778 110288 151784
rect 110248 146418 110276 151778
rect 110340 150278 110368 151846
rect 110432 151842 110460 151966
rect 110524 151910 110552 152322
rect 110512 151904 110564 151910
rect 110512 151846 110564 151852
rect 110420 151836 110472 151842
rect 110984 151814 111012 153138
rect 110984 151786 111196 151814
rect 110420 151778 110472 151784
rect 110972 151088 111024 151094
rect 110972 151030 111024 151036
rect 110328 150272 110380 150278
rect 110328 150214 110380 150220
rect 110984 147393 111012 151030
rect 111062 150512 111118 150521
rect 111062 150447 111118 150456
rect 110970 147384 111026 147393
rect 110970 147319 111026 147328
rect 110326 146432 110382 146441
rect 110248 146390 110326 146418
rect 110326 146367 110382 146376
rect 109696 132466 110368 132494
rect 110340 106321 110368 132466
rect 110326 106312 110382 106321
rect 110326 106247 110382 106256
rect 111076 89690 111104 150447
rect 111168 148374 111196 151786
rect 112812 151768 112864 151774
rect 112812 151710 112864 151716
rect 112720 151292 112772 151298
rect 112720 151234 112772 151240
rect 112628 151224 112680 151230
rect 112628 151166 112680 151172
rect 112536 151156 112588 151162
rect 112536 151098 112588 151104
rect 112444 151020 112496 151026
rect 112444 150962 112496 150968
rect 111708 150952 111760 150958
rect 111708 150894 111760 150900
rect 111616 150884 111668 150890
rect 111616 150826 111668 150832
rect 111524 150816 111576 150822
rect 111524 150758 111576 150764
rect 111432 150748 111484 150754
rect 111432 150690 111484 150696
rect 111248 150680 111300 150686
rect 111248 150622 111300 150628
rect 111338 150648 111394 150657
rect 111156 148368 111208 148374
rect 111156 148310 111208 148316
rect 111260 148186 111288 150622
rect 111338 150583 111394 150592
rect 111168 148158 111288 148186
rect 111168 109002 111196 148158
rect 111352 148050 111380 150583
rect 111260 148022 111380 148050
rect 111156 108996 111208 109002
rect 111156 108938 111208 108944
rect 111260 92478 111288 148022
rect 111444 147914 111472 150690
rect 111352 147886 111472 147914
rect 111352 111790 111380 147886
rect 111536 147778 111564 150758
rect 111444 147750 111564 147778
rect 111444 113150 111472 147750
rect 111628 147642 111656 150826
rect 111536 147614 111656 147642
rect 111536 114510 111564 147614
rect 111720 147506 111748 150894
rect 111628 147478 111748 147506
rect 111628 117298 111656 147478
rect 111706 147384 111762 147393
rect 111706 147319 111762 147328
rect 111720 121446 111748 147319
rect 111708 121440 111760 121446
rect 111708 121382 111760 121388
rect 112456 118658 112484 150962
rect 112548 122806 112576 151098
rect 112640 124166 112668 151166
rect 112732 126954 112760 151234
rect 112824 133890 112852 151710
rect 116032 151700 116084 151706
rect 116032 151642 116084 151648
rect 115296 151632 115348 151638
rect 115296 151574 115348 151580
rect 113088 151564 113140 151570
rect 113088 151506 113140 151512
rect 112996 150612 113048 150618
rect 112996 150554 113048 150560
rect 112904 150340 112956 150346
rect 112904 150282 112956 150288
rect 112812 133884 112864 133890
rect 112812 133826 112864 133832
rect 112916 132462 112944 150282
rect 113008 137970 113036 150554
rect 113100 140758 113128 151506
rect 115204 150544 115256 150550
rect 115204 150486 115256 150492
rect 113822 144256 113878 144265
rect 113822 144191 113878 144200
rect 113088 140752 113140 140758
rect 113088 140694 113140 140700
rect 112996 137964 113048 137970
rect 112996 137906 113048 137912
rect 112904 132456 112956 132462
rect 112904 132398 112956 132404
rect 112720 126948 112772 126954
rect 112720 126890 112772 126896
rect 112628 124160 112680 124166
rect 112628 124102 112680 124108
rect 112536 122800 112588 122806
rect 112536 122742 112588 122748
rect 112444 118652 112496 118658
rect 112444 118594 112496 118600
rect 111616 117292 111668 117298
rect 111616 117234 111668 117240
rect 111524 114504 111576 114510
rect 111524 114446 111576 114452
rect 111432 113144 111484 113150
rect 111432 113086 111484 113092
rect 111340 111784 111392 111790
rect 111340 111726 111392 111732
rect 111248 92472 111300 92478
rect 111248 92414 111300 92420
rect 111064 89684 111116 89690
rect 111064 89626 111116 89632
rect 113836 88330 113864 144191
rect 115216 135561 115244 150486
rect 115308 141409 115336 151574
rect 116044 143313 116072 151642
rect 116952 151496 117004 151502
rect 116952 151438 117004 151444
rect 116768 151428 116820 151434
rect 116768 151370 116820 151376
rect 116676 151360 116728 151366
rect 116676 151302 116728 151308
rect 116124 150476 116176 150482
rect 116124 150418 116176 150424
rect 116136 145217 116164 150418
rect 116492 150068 116544 150074
rect 116492 150010 116544 150016
rect 116122 145208 116178 145217
rect 116122 145143 116178 145152
rect 116030 143304 116086 143313
rect 116030 143239 116086 143248
rect 115294 141400 115350 141409
rect 115294 141335 115350 141344
rect 116124 140752 116176 140758
rect 116124 140694 116176 140700
rect 116136 139505 116164 140694
rect 116122 139496 116178 139505
rect 116122 139431 116178 139440
rect 116124 137964 116176 137970
rect 116124 137906 116176 137912
rect 116136 137601 116164 137906
rect 116122 137592 116178 137601
rect 116122 137527 116178 137536
rect 115202 135552 115258 135561
rect 115202 135487 115258 135496
rect 116032 133884 116084 133890
rect 116032 133826 116084 133832
rect 116044 133657 116072 133826
rect 116030 133648 116086 133657
rect 116030 133583 116086 133592
rect 114190 132832 114246 132841
rect 114190 132767 114246 132776
rect 114204 132666 114232 132767
rect 114192 132660 114244 132666
rect 114192 132602 114244 132608
rect 115204 132660 115256 132666
rect 115204 132602 115256 132608
rect 113914 121408 113970 121417
rect 113914 121343 113970 121352
rect 113824 88324 113876 88330
rect 113824 88266 113876 88272
rect 113928 83978 113956 121343
rect 114006 110120 114062 110129
rect 114006 110055 114062 110064
rect 113916 83972 113968 83978
rect 113916 83914 113968 83920
rect 114020 82822 114048 110055
rect 114098 98696 114154 98705
rect 114098 98631 114154 98640
rect 114008 82816 114060 82822
rect 114008 82758 114060 82764
rect 114112 80034 114140 98631
rect 114190 87272 114246 87281
rect 114190 87207 114246 87216
rect 114100 80028 114152 80034
rect 114100 79970 114152 79976
rect 114204 78674 114232 87207
rect 115216 85649 115244 132602
rect 116124 132456 116176 132462
rect 116124 132398 116176 132404
rect 116136 131753 116164 132398
rect 116122 131744 116178 131753
rect 116122 131679 116178 131688
rect 116504 129849 116532 150010
rect 116582 149696 116638 149705
rect 116582 149631 116638 149640
rect 116490 129840 116546 129849
rect 116490 129775 116546 129784
rect 116124 126948 116176 126954
rect 116124 126890 116176 126896
rect 116136 126041 116164 126890
rect 116122 126032 116178 126041
rect 116122 125967 116178 125976
rect 116124 124160 116176 124166
rect 116122 124128 116124 124137
rect 116176 124128 116178 124137
rect 116122 124063 116178 124072
rect 115940 122800 115992 122806
rect 115940 122742 115992 122748
rect 115952 122233 115980 122742
rect 115938 122224 115994 122233
rect 115938 122159 115994 122168
rect 116124 121440 116176 121446
rect 116124 121382 116176 121388
rect 116136 120193 116164 121382
rect 116122 120184 116178 120193
rect 116122 120119 116178 120128
rect 116124 118652 116176 118658
rect 116124 118594 116176 118600
rect 116136 118289 116164 118594
rect 116122 118280 116178 118289
rect 116122 118215 116178 118224
rect 116124 117292 116176 117298
rect 116124 117234 116176 117240
rect 116136 116385 116164 117234
rect 116122 116376 116178 116385
rect 116122 116311 116178 116320
rect 116124 114504 116176 114510
rect 116122 114472 116124 114481
rect 116176 114472 116178 114481
rect 116122 114407 116178 114416
rect 115940 113144 115992 113150
rect 115940 113086 115992 113092
rect 115952 112577 115980 113086
rect 115938 112568 115994 112577
rect 115938 112503 115994 112512
rect 116124 111784 116176 111790
rect 116124 111726 116176 111732
rect 116136 110673 116164 111726
rect 116122 110664 116178 110673
rect 116122 110599 116178 110608
rect 116124 108996 116176 109002
rect 116124 108938 116176 108944
rect 116136 108769 116164 108938
rect 116122 108760 116178 108769
rect 116122 108695 116178 108704
rect 116596 93401 116624 149631
rect 116688 95305 116716 151302
rect 116780 97209 116808 151370
rect 116860 150204 116912 150210
rect 116860 150146 116912 150152
rect 116872 99113 116900 150146
rect 116964 102921 116992 151438
rect 117136 150272 117188 150278
rect 117136 150214 117188 150220
rect 117044 148368 117096 148374
rect 117044 148310 117096 148316
rect 116950 102912 117006 102921
rect 116950 102847 117006 102856
rect 117056 101017 117084 148310
rect 117148 104825 117176 150214
rect 117228 150136 117280 150142
rect 117228 150078 117280 150084
rect 117240 132546 117268 150078
rect 118896 149954 118924 157966
rect 119712 154624 119764 154630
rect 119712 154566 119764 154572
rect 119724 154426 119752 154566
rect 119620 154420 119672 154426
rect 119620 154362 119672 154368
rect 119712 154420 119764 154426
rect 119712 154362 119764 154368
rect 119632 153882 119660 154362
rect 119528 153876 119580 153882
rect 119528 153818 119580 153824
rect 119620 153876 119672 153882
rect 119620 153818 119672 153824
rect 119540 149954 119568 153818
rect 120092 152386 120120 163254
rect 120552 163146 120580 163254
rect 120630 163200 120686 164400
rect 121458 163200 121514 164400
rect 122286 163200 122342 164400
rect 123114 163200 123170 164400
rect 124034 163200 124090 164400
rect 124862 163200 124918 164400
rect 125690 163200 125746 164400
rect 126518 163200 126574 164400
rect 126992 163254 127296 163282
rect 120644 163146 120672 163200
rect 120552 163118 120672 163146
rect 120172 156664 120224 156670
rect 120172 156606 120224 156612
rect 120080 152380 120132 152386
rect 120080 152322 120132 152328
rect 120184 149954 120212 156606
rect 121472 156058 121500 163200
rect 121644 158976 121696 158982
rect 121644 158918 121696 158924
rect 121460 156052 121512 156058
rect 121460 155994 121512 156000
rect 121656 153785 121684 158918
rect 122012 155304 122064 155310
rect 122012 155246 122064 155252
rect 121458 153776 121514 153785
rect 121458 153711 121514 153720
rect 121642 153776 121698 153785
rect 121642 153711 121698 153720
rect 120816 152516 120868 152522
rect 120816 152458 120868 152464
rect 120828 149954 120856 152458
rect 121472 149954 121500 153711
rect 122024 149954 122052 155246
rect 122300 154970 122328 163200
rect 123128 159390 123156 163200
rect 122840 159384 122892 159390
rect 122840 159326 122892 159332
rect 123116 159384 123168 159390
rect 123116 159326 123168 159332
rect 122288 154964 122340 154970
rect 122288 154906 122340 154912
rect 122852 150550 122880 159326
rect 124048 158982 124076 163200
rect 124036 158976 124088 158982
rect 124036 158918 124088 158924
rect 124876 156670 124904 163200
rect 125508 158908 125560 158914
rect 125508 158850 125560 158856
rect 124864 156664 124916 156670
rect 124864 156606 124916 156612
rect 124588 155440 124640 155446
rect 124588 155382 124640 155388
rect 122932 155236 122984 155242
rect 122932 155178 122984 155184
rect 122840 150544 122892 150550
rect 122840 150486 122892 150492
rect 122944 149954 122972 155178
rect 124220 153944 124272 153950
rect 124220 153886 124272 153892
rect 123392 150544 123444 150550
rect 123392 150486 123444 150492
rect 123404 149954 123432 150486
rect 124232 149954 124260 153886
rect 124600 149954 124628 155382
rect 125520 153950 125548 158850
rect 125704 155242 125732 163200
rect 126532 159730 126560 163200
rect 126428 159724 126480 159730
rect 126428 159666 126480 159672
rect 126520 159724 126572 159730
rect 126520 159666 126572 159672
rect 126440 159526 126468 159666
rect 126428 159520 126480 159526
rect 126428 159462 126480 159468
rect 126244 159452 126296 159458
rect 126244 159394 126296 159400
rect 125784 155372 125836 155378
rect 125784 155314 125836 155320
rect 125692 155236 125744 155242
rect 125692 155178 125744 155184
rect 125508 153944 125560 153950
rect 125508 153886 125560 153892
rect 125796 149954 125824 155314
rect 126256 152425 126284 159394
rect 126612 154012 126664 154018
rect 126612 153954 126664 153960
rect 125966 152416 126022 152425
rect 125966 152351 126022 152360
rect 126242 152416 126298 152425
rect 126242 152351 126298 152360
rect 118896 149926 119324 149954
rect 119540 149926 119876 149954
rect 120184 149926 120520 149954
rect 120828 149926 121164 149954
rect 121472 149926 121808 149954
rect 122024 149926 122452 149954
rect 122944 149926 123096 149954
rect 123404 149926 123740 149954
rect 124232 149926 124384 149954
rect 124600 149926 125028 149954
rect 125672 149926 125824 149954
rect 125980 149954 126008 152351
rect 126624 149954 126652 153954
rect 126992 152522 127020 163254
rect 127268 163146 127296 163254
rect 127346 163200 127402 164400
rect 128174 163200 128230 164400
rect 129002 163200 129058 164400
rect 129922 163200 129978 164400
rect 130750 163200 130806 164400
rect 131578 163200 131634 164400
rect 132406 163200 132462 164400
rect 133234 163200 133290 164400
rect 134062 163200 134118 164400
rect 134890 163200 134946 164400
rect 135810 163200 135866 164400
rect 136638 163200 136694 164400
rect 136744 163254 137416 163282
rect 127360 163146 127388 163200
rect 127268 163118 127388 163146
rect 127624 159520 127676 159526
rect 127624 159462 127676 159468
rect 127164 156732 127216 156738
rect 127164 156674 127216 156680
rect 126980 152516 127032 152522
rect 126980 152458 127032 152464
rect 127176 149954 127204 156674
rect 127636 154018 127664 159462
rect 128188 156738 128216 163200
rect 128176 156732 128228 156738
rect 128176 156674 128228 156680
rect 129016 155310 129044 163200
rect 129936 159526 129964 163200
rect 129924 159520 129976 159526
rect 129924 159462 129976 159468
rect 130764 159458 130792 163200
rect 129740 159452 129792 159458
rect 129740 159394 129792 159400
rect 130752 159452 130804 159458
rect 130752 159394 130804 159400
rect 129004 155304 129056 155310
rect 129004 155246 129056 155252
rect 129188 154080 129240 154086
rect 129188 154022 129240 154028
rect 127624 154012 127676 154018
rect 127624 153954 127676 153960
rect 128542 152552 128598 152561
rect 128542 152487 128598 152496
rect 127900 151836 127952 151842
rect 127900 151778 127952 151784
rect 127912 149954 127940 151778
rect 128556 149954 128584 152487
rect 129200 149954 129228 154022
rect 129292 154018 129504 154034
rect 129280 154012 129516 154018
rect 129332 154006 129464 154012
rect 129280 153954 129332 153960
rect 129464 153954 129516 153960
rect 129752 151842 129780 159394
rect 131026 159352 131082 159361
rect 131026 159287 131082 159296
rect 129832 156800 129884 156806
rect 129832 156742 129884 156748
rect 129740 151836 129792 151842
rect 129740 151778 129792 151784
rect 129844 149954 129872 156742
rect 130568 152244 130620 152250
rect 130568 152186 130620 152192
rect 130580 149954 130608 152186
rect 131040 151814 131068 159287
rect 131592 158030 131620 163200
rect 131580 158024 131632 158030
rect 131580 157966 131632 157972
rect 132420 153950 132448 163200
rect 133248 158846 133276 163200
rect 133602 159488 133658 159497
rect 133602 159423 133658 159432
rect 133236 158840 133288 158846
rect 133236 158782 133288 158788
rect 132500 156936 132552 156942
rect 132500 156878 132552 156884
rect 132408 153944 132460 153950
rect 131762 153912 131818 153921
rect 132408 153886 132460 153892
rect 131762 153847 131818 153856
rect 131040 151786 131160 151814
rect 131132 149954 131160 151786
rect 131776 149954 131804 153847
rect 132512 149954 132540 156878
rect 132960 154760 133012 154766
rect 132960 154702 133012 154708
rect 132972 149954 133000 154702
rect 133616 153105 133644 159423
rect 133602 153096 133658 153105
rect 133602 153031 133658 153040
rect 133880 152584 133932 152590
rect 133880 152526 133932 152532
rect 133892 149954 133920 152526
rect 134076 152250 134104 163200
rect 134904 156942 134932 163200
rect 134892 156936 134944 156942
rect 134892 156878 134944 156884
rect 135824 156874 135852 163200
rect 136652 163146 136680 163200
rect 136744 163146 136772 163254
rect 136652 163118 136772 163146
rect 137388 159798 137416 163254
rect 137466 163200 137522 164400
rect 138294 163200 138350 164400
rect 139122 163200 139178 164400
rect 139950 163200 140006 164400
rect 140778 163200 140834 164400
rect 141698 163200 141754 164400
rect 142526 163200 142582 164400
rect 143354 163200 143410 164400
rect 144182 163200 144238 164400
rect 145010 163200 145066 164400
rect 145838 163200 145894 164400
rect 146666 163200 146722 164400
rect 147586 163200 147642 164400
rect 148414 163200 148470 164400
rect 149242 163200 149298 164400
rect 150070 163200 150126 164400
rect 150898 163200 150954 164400
rect 151726 163200 151782 164400
rect 151924 163254 152504 163282
rect 137284 159792 137336 159798
rect 137284 159734 137336 159740
rect 137376 159792 137428 159798
rect 137376 159734 137428 159740
rect 137296 159594 137324 159734
rect 136824 159588 136876 159594
rect 136824 159530 136876 159536
rect 137284 159588 137336 159594
rect 137284 159530 137336 159536
rect 135260 156868 135312 156874
rect 135260 156810 135312 156816
rect 135812 156868 135864 156874
rect 135812 156810 135864 156816
rect 134338 154048 134394 154057
rect 134338 153983 134394 153992
rect 134064 152244 134116 152250
rect 134064 152186 134116 152192
rect 134352 149954 134380 153983
rect 135272 150226 135300 156810
rect 136270 153096 136326 153105
rect 136270 153031 136326 153040
rect 135628 152652 135680 152658
rect 135628 152594 135680 152600
rect 135272 150198 135346 150226
rect 125980 149926 126316 149954
rect 126624 149926 126960 149954
rect 127176 149926 127604 149954
rect 127912 149926 128248 149954
rect 128556 149926 128892 149954
rect 129200 149926 129536 149954
rect 129844 149926 130180 149954
rect 130580 149926 130824 149954
rect 131132 149926 131468 149954
rect 131776 149926 132112 149954
rect 132512 149926 132756 149954
rect 132972 149926 133400 149954
rect 133892 149926 134044 149954
rect 134352 149926 134688 149954
rect 135318 149940 135346 150198
rect 135640 149954 135668 152594
rect 136284 149954 136312 153031
rect 136836 152590 136864 159530
rect 137192 159452 137244 159458
rect 137192 159394 137244 159400
rect 137204 158914 137232 159394
rect 137480 159390 137508 163200
rect 137468 159384 137520 159390
rect 137468 159326 137520 159332
rect 137100 158908 137152 158914
rect 137100 158850 137152 158856
rect 137192 158908 137244 158914
rect 137192 158850 137244 158856
rect 137112 158794 137140 158850
rect 137112 158766 137508 158794
rect 137376 157004 137428 157010
rect 137376 156946 137428 156952
rect 137008 154216 137060 154222
rect 137060 154164 137324 154170
rect 137008 154158 137324 154164
rect 136916 154148 136968 154154
rect 137020 154142 137324 154158
rect 136916 154090 136968 154096
rect 136824 152584 136876 152590
rect 136824 152526 136876 152532
rect 136928 149954 136956 154090
rect 137296 154086 137324 154142
rect 137284 154080 137336 154086
rect 137284 154022 137336 154028
rect 137388 151814 137416 156946
rect 137480 153950 137508 158766
rect 138308 157010 138336 163200
rect 138386 159624 138442 159633
rect 138386 159559 138442 159568
rect 138400 157334 138428 159559
rect 138400 157306 138612 157334
rect 138296 157004 138348 157010
rect 138296 156946 138348 156952
rect 137928 154352 137980 154358
rect 137928 154294 137980 154300
rect 138112 154352 138164 154358
rect 138112 154294 138164 154300
rect 137940 154057 137968 154294
rect 138124 154170 138152 154294
rect 138032 154142 138152 154170
rect 138032 154086 138060 154142
rect 138020 154080 138072 154086
rect 137926 154048 137982 154057
rect 138020 154022 138072 154028
rect 137926 153983 137982 153992
rect 137468 153944 137520 153950
rect 137468 153886 137520 153892
rect 138204 153876 138256 153882
rect 138204 153818 138256 153824
rect 138110 153640 138166 153649
rect 138110 153575 138166 153584
rect 138124 153270 138152 153575
rect 138216 153270 138244 153818
rect 138112 153264 138164 153270
rect 138112 153206 138164 153212
rect 138204 153264 138256 153270
rect 138204 153206 138256 153212
rect 138584 152862 138612 157306
rect 139136 156806 139164 163200
rect 139964 159798 139992 163200
rect 140792 161474 140820 163200
rect 140792 161446 140912 161474
rect 139676 159792 139728 159798
rect 139676 159734 139728 159740
rect 139952 159792 140004 159798
rect 139952 159734 140004 159740
rect 139124 156800 139176 156806
rect 139124 156742 139176 156748
rect 139308 154828 139360 154834
rect 139308 154770 139360 154776
rect 138296 152856 138348 152862
rect 138296 152798 138348 152804
rect 138572 152856 138624 152862
rect 138572 152798 138624 152804
rect 138308 152590 138336 152798
rect 138848 152788 138900 152794
rect 138848 152730 138900 152736
rect 138296 152584 138348 152590
rect 138296 152526 138348 152532
rect 138296 151904 138348 151910
rect 138296 151846 138348 151852
rect 137388 151786 137508 151814
rect 137480 149954 137508 151786
rect 138308 149954 138336 151846
rect 138860 149954 138888 152730
rect 139320 151910 139348 154770
rect 139688 154358 139716 159734
rect 140134 156632 140190 156641
rect 140134 156567 140190 156576
rect 139492 154352 139544 154358
rect 139492 154294 139544 154300
rect 139676 154352 139728 154358
rect 139676 154294 139728 154300
rect 139308 151904 139360 151910
rect 139308 151846 139360 151852
rect 139504 149954 139532 154294
rect 140148 149954 140176 156567
rect 140884 152794 140912 161446
rect 141712 157418 141740 163200
rect 141700 157412 141752 157418
rect 141700 157354 141752 157360
rect 142540 155378 142568 163200
rect 143368 159662 143396 163200
rect 144196 161474 144224 163200
rect 144196 161446 144408 161474
rect 143264 159656 143316 159662
rect 143264 159598 143316 159604
rect 143356 159656 143408 159662
rect 143356 159598 143408 159604
rect 143276 157334 143304 159598
rect 144000 159588 144052 159594
rect 144000 159530 144052 159536
rect 144184 159588 144236 159594
rect 144184 159530 144236 159536
rect 144012 159474 144040 159530
rect 144012 159446 144132 159474
rect 144196 159458 144224 159530
rect 144380 159458 144408 161446
rect 143276 157306 143396 157334
rect 143262 156768 143318 156777
rect 143262 156703 143318 156712
rect 142528 155372 142580 155378
rect 142528 155314 142580 155320
rect 142896 154488 142948 154494
rect 142896 154430 142948 154436
rect 142988 154488 143040 154494
rect 142988 154430 143040 154436
rect 142908 154222 142936 154430
rect 142896 154216 142948 154222
rect 142158 154184 142214 154193
rect 142158 154119 142214 154128
rect 142434 154184 142490 154193
rect 142896 154158 142948 154164
rect 142434 154119 142436 154128
rect 141424 152856 141476 152862
rect 141424 152798 141476 152804
rect 140872 152788 140924 152794
rect 140872 152730 140924 152736
rect 140780 152720 140832 152726
rect 140780 152662 140832 152668
rect 140792 149954 140820 152662
rect 141436 149954 141464 152798
rect 142172 149954 142200 154119
rect 142488 154119 142490 154128
rect 142436 154090 142488 154096
rect 143000 154086 143028 154430
rect 143080 154352 143132 154358
rect 143080 154294 143132 154300
rect 143092 154193 143120 154294
rect 143078 154184 143134 154193
rect 143078 154119 143134 154128
rect 142988 154080 143040 154086
rect 142988 154022 143040 154028
rect 142804 152720 142856 152726
rect 142804 152662 142856 152668
rect 142816 152046 142844 152662
rect 142804 152040 142856 152046
rect 142804 151982 142856 151988
rect 143276 149954 143304 156703
rect 143368 152046 143396 157306
rect 143448 154080 143500 154086
rect 143448 154022 143500 154028
rect 143538 154048 143594 154057
rect 143460 153649 143488 154022
rect 143538 153983 143594 153992
rect 143552 153950 143580 153983
rect 143540 153944 143592 153950
rect 143540 153886 143592 153892
rect 143446 153640 143502 153649
rect 143446 153575 143502 153584
rect 144104 152794 144132 159446
rect 144184 159452 144236 159458
rect 144184 159394 144236 159400
rect 144368 159452 144420 159458
rect 144368 159394 144420 159400
rect 145024 155990 145052 163200
rect 145102 157992 145158 158001
rect 145102 157927 145158 157936
rect 145012 155984 145064 155990
rect 145012 155926 145064 155932
rect 144000 152788 144052 152794
rect 144000 152730 144052 152736
rect 144092 152788 144144 152794
rect 144092 152730 144144 152736
rect 144012 152674 144040 152730
rect 144012 152646 144132 152674
rect 144104 152590 144132 152646
rect 144000 152584 144052 152590
rect 144000 152526 144052 152532
rect 144092 152584 144144 152590
rect 144092 152526 144144 152532
rect 143538 152416 143594 152425
rect 143538 152351 143594 152360
rect 143356 152040 143408 152046
rect 143356 151982 143408 151988
rect 135640 149926 135976 149954
rect 136284 149926 136620 149954
rect 136928 149926 137264 149954
rect 137480 149926 137908 149954
rect 138308 149926 138552 149954
rect 138860 149926 139196 149954
rect 139504 149926 139840 149954
rect 140148 149926 140484 149954
rect 140792 149926 141128 149954
rect 141436 149926 141772 149954
rect 142172 149926 142416 149954
rect 143060 149926 143304 149954
rect 143552 149954 143580 152351
rect 144012 149954 144040 152526
rect 145116 149954 145144 157927
rect 145852 155446 145880 163200
rect 146484 160064 146536 160070
rect 146484 160006 146536 160012
rect 145932 157072 145984 157078
rect 145932 157014 145984 157020
rect 145840 155440 145892 155446
rect 145840 155382 145892 155388
rect 145380 154284 145432 154290
rect 145380 154226 145432 154232
rect 145392 153950 145420 154226
rect 145288 153944 145340 153950
rect 145288 153886 145340 153892
rect 145380 153944 145432 153950
rect 145380 153886 145432 153892
rect 143552 149926 143704 149954
rect 144012 149926 144348 149954
rect 144992 149926 145144 149954
rect 145300 149954 145328 153886
rect 145944 149954 145972 157014
rect 146496 152862 146524 160006
rect 146680 158778 146708 163200
rect 146760 160064 146812 160070
rect 146760 160006 146812 160012
rect 146772 159526 146800 160006
rect 147036 159792 147088 159798
rect 147088 159740 147260 159746
rect 147036 159734 147260 159740
rect 147048 159718 147260 159734
rect 147232 159594 147260 159718
rect 147220 159588 147272 159594
rect 147220 159530 147272 159536
rect 146760 159520 146812 159526
rect 146760 159462 146812 159468
rect 147404 159520 147456 159526
rect 147404 159462 147456 159468
rect 147416 159338 147444 159462
rect 147600 159458 147628 163200
rect 147588 159452 147640 159458
rect 147588 159394 147640 159400
rect 147416 159310 148088 159338
rect 146576 158772 146628 158778
rect 146576 158714 146628 158720
rect 146668 158772 146720 158778
rect 146668 158714 146720 158720
rect 146588 158658 146616 158714
rect 146588 158630 146984 158658
rect 146760 158092 146812 158098
rect 146760 158034 146812 158040
rect 146772 157334 146800 158034
rect 146772 157306 146892 157334
rect 146484 152856 146536 152862
rect 146484 152798 146536 152804
rect 146668 152040 146720 152046
rect 146668 151982 146720 151988
rect 146680 151842 146708 151982
rect 146576 151836 146628 151842
rect 146576 151778 146628 151784
rect 146668 151836 146720 151842
rect 146668 151778 146720 151784
rect 146588 149954 146616 151778
rect 146864 150090 146892 157306
rect 146956 154290 146984 158630
rect 148060 154290 148088 159310
rect 148428 158098 148456 163200
rect 148416 158092 148468 158098
rect 148416 158034 148468 158040
rect 148232 157208 148284 157214
rect 148232 157150 148284 157156
rect 146944 154284 146996 154290
rect 146944 154226 146996 154232
rect 147956 154284 148008 154290
rect 147956 154226 148008 154232
rect 148048 154284 148100 154290
rect 148048 154226 148100 154232
rect 147968 154154 147996 154226
rect 147864 154148 147916 154154
rect 147864 154090 147916 154096
rect 147956 154148 148008 154154
rect 147956 154090 148008 154096
rect 146864 150062 147168 150090
rect 147140 149954 147168 150062
rect 147876 149954 147904 154090
rect 148244 151814 148272 157150
rect 149256 154834 149284 163200
rect 149336 159452 149388 159458
rect 149336 159394 149388 159400
rect 149244 154828 149296 154834
rect 149244 154770 149296 154776
rect 149348 152726 149376 159394
rect 149610 158264 149666 158273
rect 149610 158199 149666 158208
rect 149152 152720 149204 152726
rect 149152 152662 149204 152668
rect 149336 152720 149388 152726
rect 149336 152662 149388 152668
rect 148244 151786 148456 151814
rect 148428 149954 148456 151786
rect 149164 149954 149192 152662
rect 149624 149954 149652 158199
rect 150084 157214 150112 163200
rect 150912 159458 150940 163200
rect 150900 159452 150952 159458
rect 150900 159394 150952 159400
rect 150072 157208 150124 157214
rect 150072 157150 150124 157156
rect 150900 157140 150952 157146
rect 150900 157082 150952 157088
rect 150440 154080 150492 154086
rect 150440 154022 150492 154028
rect 150452 149954 150480 154022
rect 150912 149954 150940 157082
rect 151740 157078 151768 163200
rect 151728 157072 151780 157078
rect 151728 157014 151780 157020
rect 151924 154154 151952 163254
rect 152476 163146 152504 163254
rect 152554 163200 152610 164400
rect 153474 163200 153530 164400
rect 153672 163254 154252 163282
rect 152568 163146 152596 163200
rect 152476 163118 152596 163146
rect 153488 159798 153516 163200
rect 153476 159792 153528 159798
rect 153476 159734 153528 159740
rect 152186 158128 152242 158137
rect 152186 158063 152242 158072
rect 151912 154148 151964 154154
rect 151912 154090 151964 154096
rect 151820 152652 151872 152658
rect 151820 152594 151872 152600
rect 151832 149954 151860 152594
rect 152200 149954 152228 158063
rect 153568 157276 153620 157282
rect 153568 157218 153620 157224
rect 153292 154216 153344 154222
rect 153292 154158 153344 154164
rect 153304 150226 153332 154158
rect 153258 150198 153332 150226
rect 145300 149926 145636 149954
rect 145944 149926 146280 149954
rect 146588 149926 146924 149954
rect 147140 149926 147568 149954
rect 147876 149926 148212 149954
rect 148428 149926 148856 149954
rect 149164 149926 149500 149954
rect 149624 149926 150052 149954
rect 150452 149926 150696 149954
rect 150912 149926 151340 149954
rect 151832 149926 151984 149954
rect 152200 149926 152628 149954
rect 153258 149940 153286 150198
rect 153580 149954 153608 157218
rect 153672 152658 153700 163254
rect 154224 163146 154252 163254
rect 154302 163200 154358 164400
rect 155130 163200 155186 164400
rect 155958 163200 156014 164400
rect 156786 163200 156842 164400
rect 157614 163200 157670 164400
rect 158442 163200 158498 164400
rect 159362 163200 159418 164400
rect 160190 163200 160246 164400
rect 161018 163200 161074 164400
rect 161846 163200 161902 164400
rect 162674 163200 162730 164400
rect 163502 163200 163558 164400
rect 164330 163200 164386 164400
rect 165250 163200 165306 164400
rect 165632 163254 166028 163282
rect 154316 163146 154344 163200
rect 154224 163118 154344 163146
rect 154488 160064 154540 160070
rect 154488 160006 154540 160012
rect 154500 154630 154528 160006
rect 155144 158166 155172 163200
rect 154764 158160 154816 158166
rect 154764 158102 154816 158108
rect 155132 158160 155184 158166
rect 155132 158102 155184 158108
rect 154488 154624 154540 154630
rect 154488 154566 154540 154572
rect 153660 152652 153712 152658
rect 153660 152594 153712 152600
rect 154212 151972 154264 151978
rect 154212 151914 154264 151920
rect 154224 149954 154252 151914
rect 154776 149954 154804 158102
rect 155972 154766 156000 163200
rect 156800 160070 156828 163200
rect 156788 160064 156840 160070
rect 156788 160006 156840 160012
rect 156420 159860 156472 159866
rect 156420 159802 156472 159808
rect 156604 159860 156656 159866
rect 156604 159802 156656 159808
rect 156052 157344 156104 157350
rect 156052 157286 156104 157292
rect 155960 154760 156012 154766
rect 155960 154702 156012 154708
rect 154948 154556 155000 154562
rect 154948 154498 155000 154504
rect 154960 154154 154988 154498
rect 154948 154148 155000 154154
rect 154948 154090 155000 154096
rect 155500 153808 155552 153814
rect 155500 153750 155552 153756
rect 155512 149954 155540 153750
rect 156064 149954 156092 157286
rect 156328 154692 156380 154698
rect 156328 154634 156380 154640
rect 156340 154290 156368 154634
rect 156328 154284 156380 154290
rect 156328 154226 156380 154232
rect 156432 152046 156460 159802
rect 156512 159724 156564 159730
rect 156512 159666 156564 159672
rect 156524 157146 156552 159666
rect 156616 159662 156644 159802
rect 156604 159656 156656 159662
rect 156604 159598 156656 159604
rect 157628 159594 157656 163200
rect 157616 159588 157668 159594
rect 157616 159530 157668 159536
rect 158456 158234 158484 163200
rect 158720 158840 158772 158846
rect 158720 158782 158772 158788
rect 157340 158228 157392 158234
rect 157340 158170 157392 158176
rect 158444 158228 158496 158234
rect 158444 158170 158496 158176
rect 156512 157140 156564 157146
rect 156512 157082 156564 157088
rect 156696 154624 156748 154630
rect 156696 154566 156748 154572
rect 156512 154216 156564 154222
rect 156512 154158 156564 154164
rect 156524 153678 156552 154158
rect 156708 153678 156736 154566
rect 156788 154284 156840 154290
rect 156788 154226 156840 154232
rect 156800 153882 156828 154226
rect 156788 153876 156840 153882
rect 156788 153818 156840 153824
rect 156512 153672 156564 153678
rect 156512 153614 156564 153620
rect 156696 153672 156748 153678
rect 156696 153614 156748 153620
rect 156420 152040 156472 152046
rect 156420 151982 156472 151988
rect 156788 151836 156840 151842
rect 156788 151778 156840 151784
rect 156800 149954 156828 151778
rect 157352 149954 157380 158170
rect 158732 157350 158760 158782
rect 158720 157344 158772 157350
rect 158720 157286 158772 157292
rect 158904 157140 158956 157146
rect 158904 157082 158956 157088
rect 158916 156602 158944 157082
rect 158812 156596 158864 156602
rect 158812 156538 158864 156544
rect 158904 156596 158956 156602
rect 158904 156538 158956 156544
rect 158076 154148 158128 154154
rect 158076 154090 158128 154096
rect 158088 149954 158116 154090
rect 158824 149954 158852 156538
rect 159376 154630 159404 163200
rect 160100 159860 160152 159866
rect 160100 159802 160152 159808
rect 160112 157146 160140 159802
rect 160100 157140 160152 157146
rect 160100 157082 160152 157088
rect 159364 154624 159416 154630
rect 159364 154566 159416 154572
rect 160204 154154 160232 163200
rect 161032 159662 161060 163200
rect 161020 159656 161072 159662
rect 161020 159598 161072 159604
rect 161860 158302 161888 163200
rect 162584 159928 162636 159934
rect 162584 159870 162636 159876
rect 160284 158296 160336 158302
rect 160284 158238 160336 158244
rect 161848 158296 161900 158302
rect 161848 158238 161900 158244
rect 160192 154148 160244 154154
rect 160192 154090 160244 154096
rect 159364 152448 159416 152454
rect 159364 152390 159416 152396
rect 159376 149954 159404 152390
rect 160296 150226 160324 158238
rect 161570 156904 161626 156913
rect 161570 156839 161626 156848
rect 160650 154320 160706 154329
rect 160650 154255 160706 154264
rect 160296 150198 160370 150226
rect 153580 149926 153916 149954
rect 154224 149926 154560 149954
rect 154776 149926 155204 149954
rect 155512 149926 155848 149954
rect 156064 149926 156492 149954
rect 156800 149926 157136 149954
rect 157352 149926 157780 149954
rect 158088 149926 158424 149954
rect 158824 149926 159068 149954
rect 159376 149926 159712 149954
rect 160342 149940 160370 150198
rect 160664 149954 160692 154255
rect 161584 150226 161612 156839
rect 161940 152788 161992 152794
rect 161940 152730 161992 152736
rect 161584 150198 161658 150226
rect 160664 149926 161000 149954
rect 161630 149940 161658 150198
rect 161952 149954 161980 152730
rect 162596 151978 162624 159870
rect 162688 154698 162716 163200
rect 162872 159186 163084 159202
rect 162872 159180 163096 159186
rect 162872 159174 163044 159180
rect 162872 159118 162900 159174
rect 163044 159122 163096 159128
rect 162860 159112 162912 159118
rect 162860 159054 162912 159060
rect 163516 158846 163544 163200
rect 164148 159724 164200 159730
rect 164148 159666 164200 159672
rect 163504 158840 163556 158846
rect 163504 158782 163556 158788
rect 162858 158400 162914 158409
rect 162858 158335 162914 158344
rect 162676 154692 162728 154698
rect 162676 154634 162728 154640
rect 162676 154216 162728 154222
rect 162676 154158 162728 154164
rect 162688 153746 162716 154158
rect 162768 154080 162820 154086
rect 162768 154022 162820 154028
rect 162780 153746 162808 154022
rect 162676 153740 162728 153746
rect 162676 153682 162728 153688
rect 162768 153740 162820 153746
rect 162768 153682 162820 153688
rect 162584 151972 162636 151978
rect 162584 151914 162636 151920
rect 162872 150226 162900 158335
rect 164160 157282 164188 159666
rect 164148 157276 164200 157282
rect 164148 157218 164200 157224
rect 163780 156528 163832 156534
rect 163780 156470 163832 156476
rect 163228 154284 163280 154290
rect 163228 154226 163280 154232
rect 162872 150198 162946 150226
rect 161952 149926 162288 149954
rect 162918 149940 162946 150198
rect 163240 149954 163268 154226
rect 163792 149954 163820 156470
rect 164344 152794 164372 163200
rect 165264 158438 165292 163200
rect 165068 158432 165120 158438
rect 165068 158374 165120 158380
rect 165252 158432 165304 158438
rect 165252 158374 165304 158380
rect 164332 152788 164384 152794
rect 164332 152730 164384 152736
rect 164516 152108 164568 152114
rect 164516 152050 164568 152056
rect 164528 149954 164556 152050
rect 165080 149954 165108 158374
rect 165632 154154 165660 163254
rect 166000 163146 166028 163254
rect 166078 163200 166134 164400
rect 166906 163200 166962 164400
rect 167734 163200 167790 164400
rect 168562 163200 168618 164400
rect 169390 163200 169446 164400
rect 170218 163200 170274 164400
rect 171138 163200 171194 164400
rect 171966 163200 172022 164400
rect 172532 163254 172744 163282
rect 166092 163146 166120 163200
rect 166000 163118 166120 163146
rect 166920 159934 166948 163200
rect 166908 159928 166960 159934
rect 166908 159870 166960 159876
rect 167748 159730 167776 163200
rect 167736 159724 167788 159730
rect 167736 159666 167788 159672
rect 167000 159316 167052 159322
rect 167000 159258 167052 159264
rect 166264 157276 166316 157282
rect 166264 157218 166316 157224
rect 165896 157140 165948 157146
rect 165896 157082 165948 157088
rect 165988 157140 166040 157146
rect 165988 157082 166040 157088
rect 165908 156534 165936 157082
rect 165896 156528 165948 156534
rect 165896 156470 165948 156476
rect 166000 156466 166028 157082
rect 166276 156534 166304 157218
rect 166264 156528 166316 156534
rect 166264 156470 166316 156476
rect 165988 156460 166040 156466
rect 165988 156402 166040 156408
rect 166354 155408 166410 155417
rect 166354 155343 166410 155352
rect 165804 154216 165856 154222
rect 165804 154158 165856 154164
rect 165620 154148 165672 154154
rect 165620 154090 165672 154096
rect 165816 149954 165844 154158
rect 166368 149954 166396 155343
rect 167012 152454 167040 159258
rect 168576 158370 168604 163200
rect 167552 158364 167604 158370
rect 167552 158306 167604 158312
rect 168564 158364 168616 158370
rect 168564 158306 168616 158312
rect 167092 152856 167144 152862
rect 167092 152798 167144 152804
rect 167000 152448 167052 152454
rect 167000 152390 167052 152396
rect 167104 149954 167132 152798
rect 167564 151814 167592 158306
rect 169022 155544 169078 155553
rect 168564 155508 168616 155514
rect 169404 155514 169432 163200
rect 170232 159322 170260 163200
rect 170220 159316 170272 159322
rect 170220 159258 170272 159264
rect 171152 159118 171180 163200
rect 169852 159112 169904 159118
rect 169852 159054 169904 159060
rect 171140 159112 171192 159118
rect 171140 159054 171192 159060
rect 169022 155479 169078 155488
rect 169392 155508 169444 155514
rect 168564 155450 168616 155456
rect 167564 151786 167684 151814
rect 167656 149954 167684 151786
rect 168576 149954 168604 155450
rect 169036 149954 169064 155479
rect 169392 155450 169444 155456
rect 169760 152176 169812 152182
rect 169760 152118 169812 152124
rect 169772 149954 169800 152118
rect 169864 152114 169892 159054
rect 171980 158642 172008 163200
rect 172428 159180 172480 159186
rect 172428 159122 172480 159128
rect 170220 158636 170272 158642
rect 170220 158578 170272 158584
rect 171968 158636 172020 158642
rect 171968 158578 172020 158584
rect 169852 152108 169904 152114
rect 169852 152050 169904 152056
rect 170232 149954 170260 158578
rect 171600 157140 171652 157146
rect 171600 157082 171652 157088
rect 171230 155272 171286 155281
rect 171230 155207 171286 155216
rect 171244 150226 171272 155207
rect 171244 150198 171318 150226
rect 163240 149926 163576 149954
rect 163792 149926 164220 149954
rect 164528 149926 164864 149954
rect 165080 149926 165508 149954
rect 165816 149926 166152 149954
rect 166368 149926 166796 149954
rect 167104 149926 167440 149954
rect 167656 149926 168084 149954
rect 168576 149926 168728 149954
rect 169036 149926 169372 149954
rect 169772 149926 170016 149954
rect 170232 149926 170660 149954
rect 171290 149940 171318 150198
rect 171612 149954 171640 157082
rect 172440 151842 172468 159122
rect 172532 154222 172560 163254
rect 172716 163146 172744 163254
rect 172794 163200 172850 164400
rect 173622 163200 173678 164400
rect 173912 163254 174400 163282
rect 172808 163146 172836 163200
rect 172716 163118 172836 163146
rect 173636 159118 173664 163200
rect 172704 159112 172756 159118
rect 172704 159054 172756 159060
rect 173624 159112 173676 159118
rect 173624 159054 173676 159060
rect 172520 154216 172572 154222
rect 172520 154158 172572 154164
rect 172716 152182 172744 159054
rect 172796 158500 172848 158506
rect 172796 158442 172848 158448
rect 172704 152176 172756 152182
rect 172704 152118 172756 152124
rect 172520 152040 172572 152046
rect 172520 151982 172572 151988
rect 172428 151836 172480 151842
rect 172428 151778 172480 151784
rect 172532 150226 172560 151982
rect 172532 150198 172606 150226
rect 171612 149926 171948 149954
rect 172578 149940 172606 150198
rect 172808 149954 172836 158442
rect 173532 155644 173584 155650
rect 173532 155586 173584 155592
rect 173544 149954 173572 155586
rect 173912 152862 173940 163254
rect 174372 163146 174400 163254
rect 174450 163200 174506 164400
rect 175278 163200 175334 164400
rect 176106 163200 176162 164400
rect 177026 163200 177082 164400
rect 177854 163200 177910 164400
rect 178682 163200 178738 164400
rect 179510 163200 179566 164400
rect 180338 163200 180394 164400
rect 180812 163254 181116 163282
rect 174464 163146 174492 163200
rect 174372 163118 174492 163146
rect 175292 158506 175320 163200
rect 176120 161474 176148 163200
rect 176120 161446 176332 161474
rect 175372 158568 175424 158574
rect 175372 158510 175424 158516
rect 175280 158500 175332 158506
rect 175280 158442 175332 158448
rect 174082 157040 174138 157049
rect 174082 156975 174138 156984
rect 173900 152856 173952 152862
rect 173900 152798 173952 152804
rect 174096 149954 174124 156975
rect 174820 153128 174872 153134
rect 174820 153070 174872 153076
rect 174832 149954 174860 153070
rect 175384 149954 175412 158510
rect 176200 157956 176252 157962
rect 176200 157898 176252 157904
rect 175924 157888 175976 157894
rect 176212 157842 176240 157898
rect 175976 157836 176240 157842
rect 175924 157830 176240 157836
rect 175936 157814 176240 157830
rect 176304 155650 176332 161446
rect 176660 158772 176712 158778
rect 176660 158714 176712 158720
rect 176292 155644 176344 155650
rect 176292 155586 176344 155592
rect 176016 155576 176068 155582
rect 176016 155518 176068 155524
rect 175924 152448 175976 152454
rect 175924 152390 175976 152396
rect 175936 152114 175964 152390
rect 175924 152108 175976 152114
rect 175924 152050 175976 152056
rect 176028 149954 176056 155518
rect 176672 154290 176700 158714
rect 177040 157146 177068 163200
rect 177868 159798 177896 163200
rect 177856 159792 177908 159798
rect 177856 159734 177908 159740
rect 178696 158574 178724 163200
rect 178684 158568 178736 158574
rect 178684 158510 178736 158516
rect 178040 157888 178092 157894
rect 178040 157830 178092 157836
rect 177028 157140 177080 157146
rect 177028 157082 177080 157088
rect 176842 155816 176898 155825
rect 176842 155751 176898 155760
rect 176660 154284 176712 154290
rect 176660 154226 176712 154232
rect 176108 152448 176160 152454
rect 176108 152390 176160 152396
rect 176120 152182 176148 152390
rect 176108 152176 176160 152182
rect 176108 152118 176160 152124
rect 176200 152176 176252 152182
rect 176200 152118 176252 152124
rect 176212 151842 176240 152118
rect 176200 151836 176252 151842
rect 176200 151778 176252 151784
rect 176856 149954 176884 155751
rect 177396 151972 177448 151978
rect 177396 151914 177448 151920
rect 177408 149954 177436 151914
rect 178052 149954 178080 157830
rect 178682 155680 178738 155689
rect 178682 155615 178738 155624
rect 178696 149954 178724 155615
rect 179524 155582 179552 163200
rect 180352 158778 180380 163200
rect 180708 159860 180760 159866
rect 180708 159802 180760 159808
rect 180340 158772 180392 158778
rect 180340 158714 180392 158720
rect 180720 157894 180748 159802
rect 180708 157888 180760 157894
rect 180708 157830 180760 157836
rect 179512 155576 179564 155582
rect 179512 155518 179564 155524
rect 179512 154284 179564 154290
rect 179512 154226 179564 154232
rect 179524 153610 179552 154226
rect 179420 153604 179472 153610
rect 179420 153546 179472 153552
rect 179512 153604 179564 153610
rect 179512 153546 179564 153552
rect 179432 149954 179460 153546
rect 180812 153134 180840 163254
rect 181088 163146 181116 163254
rect 181166 163200 181222 164400
rect 181994 163200 182050 164400
rect 182192 163254 182864 163282
rect 181180 163146 181208 163200
rect 181088 163118 181208 163146
rect 182008 158710 182036 163200
rect 180892 158704 180944 158710
rect 180892 158646 180944 158652
rect 181996 158704 182048 158710
rect 181996 158646 182048 158652
rect 180800 153128 180852 153134
rect 180800 153070 180852 153076
rect 179972 152312 180024 152318
rect 179972 152254 180024 152260
rect 179984 149954 180012 152254
rect 180904 150226 180932 158646
rect 181088 157950 181576 157978
rect 181088 157758 181116 157950
rect 181548 157894 181576 157950
rect 181352 157888 181404 157894
rect 181352 157830 181404 157836
rect 181536 157888 181588 157894
rect 181536 157830 181588 157836
rect 181076 157752 181128 157758
rect 181076 157694 181128 157700
rect 181364 157706 181392 157830
rect 181812 157820 181864 157826
rect 181812 157762 181864 157768
rect 181720 157752 181772 157758
rect 181364 157700 181720 157706
rect 181364 157694 181772 157700
rect 181168 157684 181220 157690
rect 181364 157678 181760 157694
rect 181168 157626 181220 157632
rect 181180 157570 181208 157626
rect 181824 157570 181852 157762
rect 181180 157542 181852 157570
rect 181812 156392 181864 156398
rect 181812 156334 181864 156340
rect 181168 155712 181220 155718
rect 181168 155654 181220 155660
rect 180858 150198 180932 150226
rect 172808 149926 173236 149954
rect 173544 149926 173880 149954
rect 174096 149926 174524 149954
rect 174832 149926 175168 149954
rect 175384 149926 175812 149954
rect 176028 149926 176456 149954
rect 176856 149926 177100 149954
rect 177408 149926 177744 149954
rect 178052 149926 178388 149954
rect 178696 149926 179032 149954
rect 179432 149926 179676 149954
rect 179984 149926 180320 149954
rect 180858 149940 180886 150198
rect 181180 149954 181208 155654
rect 181824 149954 181852 156334
rect 182192 154290 182220 163254
rect 182836 163146 182864 163254
rect 182914 163200 182970 164400
rect 183742 163200 183798 164400
rect 184570 163200 184626 164400
rect 185398 163200 185454 164400
rect 186226 163200 186282 164400
rect 187054 163200 187110 164400
rect 187882 163200 187938 164400
rect 188802 163200 188858 164400
rect 189630 163200 189686 164400
rect 190458 163200 190514 164400
rect 191286 163200 191342 164400
rect 192114 163200 192170 164400
rect 192942 163200 192998 164400
rect 193770 163200 193826 164400
rect 194690 163200 194746 164400
rect 195518 163200 195574 164400
rect 196346 163200 196402 164400
rect 197174 163200 197230 164400
rect 198002 163200 198058 164400
rect 198830 163200 198886 164400
rect 199658 163200 199714 164400
rect 200578 163200 200634 164400
rect 201406 163200 201462 164400
rect 202234 163200 202290 164400
rect 203062 163200 203118 164400
rect 203890 163200 203946 164400
rect 204718 163200 204774 164400
rect 205008 163254 205496 163282
rect 182928 163146 182956 163200
rect 182836 163118 182956 163146
rect 183756 159050 183784 163200
rect 184584 159866 184612 163200
rect 184572 159860 184624 159866
rect 184572 159802 184624 159808
rect 184664 159248 184716 159254
rect 184664 159190 184716 159196
rect 182548 159044 182600 159050
rect 182548 158986 182600 158992
rect 183744 159044 183796 159050
rect 183744 158986 183796 158992
rect 182180 154284 182232 154290
rect 182180 154226 182232 154232
rect 182560 152114 182588 158986
rect 183008 157956 183060 157962
rect 183008 157898 183060 157904
rect 182456 152108 182508 152114
rect 182456 152050 182508 152056
rect 182548 152108 182600 152114
rect 182548 152050 182600 152056
rect 182468 149954 182496 152050
rect 183020 149954 183048 157898
rect 183742 155952 183798 155961
rect 183742 155887 183798 155896
rect 183756 149954 183784 155887
rect 184386 154456 184442 154465
rect 184386 154391 184442 154400
rect 184400 149954 184428 154391
rect 184676 151978 184704 159190
rect 185412 157962 185440 163200
rect 185400 157956 185452 157962
rect 185400 157898 185452 157904
rect 185584 157684 185636 157690
rect 185584 157626 185636 157632
rect 185032 152040 185084 152046
rect 185032 151982 185084 151988
rect 184664 151972 184716 151978
rect 184664 151914 184716 151920
rect 185044 149954 185072 151982
rect 185596 149954 185624 157626
rect 186240 155718 186268 163200
rect 186412 159928 186464 159934
rect 186412 159870 186464 159876
rect 186424 157334 186452 159870
rect 187068 159254 187096 163200
rect 187056 159248 187108 159254
rect 187056 159190 187108 159196
rect 186424 157306 186728 157334
rect 186332 155922 186636 155938
rect 186332 155916 186648 155922
rect 186332 155910 186596 155916
rect 186228 155712 186280 155718
rect 186228 155654 186280 155660
rect 186332 155038 186360 155910
rect 186596 155858 186648 155864
rect 186412 155848 186464 155854
rect 186412 155790 186464 155796
rect 186320 155032 186372 155038
rect 186320 154974 186372 154980
rect 186424 149954 186452 155790
rect 186700 154902 186728 157306
rect 186964 155168 187016 155174
rect 186964 155110 187016 155116
rect 186780 155100 186832 155106
rect 186780 155042 186832 155048
rect 186596 154896 186648 154902
rect 186596 154838 186648 154844
rect 186688 154896 186740 154902
rect 186688 154838 186740 154844
rect 186608 154714 186636 154838
rect 186792 154714 186820 155042
rect 186608 154686 186820 154714
rect 186976 149954 187004 155110
rect 187700 152992 187752 152998
rect 187700 152934 187752 152940
rect 187712 149954 187740 152934
rect 187896 152318 187924 163200
rect 188816 157894 188844 163200
rect 188160 157888 188212 157894
rect 188160 157830 188212 157836
rect 188804 157888 188856 157894
rect 188804 157830 188856 157836
rect 187884 152312 187936 152318
rect 187884 152254 187936 152260
rect 188172 149954 188200 157830
rect 189080 155848 189132 155854
rect 189080 155790 189132 155796
rect 189092 149954 189120 155790
rect 189644 155174 189672 163200
rect 190472 157758 190500 163200
rect 191300 159934 191328 163200
rect 191748 160064 191800 160070
rect 191748 160006 191800 160012
rect 191656 159996 191708 160002
rect 191656 159938 191708 159944
rect 191288 159928 191340 159934
rect 191288 159870 191340 159876
rect 190644 157820 190696 157826
rect 190644 157762 190696 157768
rect 190460 157752 190512 157758
rect 190460 157694 190512 157700
rect 190656 157334 190684 157762
rect 190656 157306 190776 157334
rect 189632 155168 189684 155174
rect 189632 155110 189684 155116
rect 189540 154420 189592 154426
rect 189540 154362 189592 154368
rect 189552 149954 189580 154362
rect 190184 152176 190236 152182
rect 190184 152118 190236 152124
rect 190196 149954 190224 152118
rect 190748 149954 190776 157306
rect 191472 155032 191524 155038
rect 191472 154974 191524 154980
rect 191104 154488 191156 154494
rect 191104 154430 191156 154436
rect 191012 154420 191064 154426
rect 191012 154362 191064 154368
rect 191024 153814 191052 154362
rect 191116 153814 191144 154430
rect 191288 154420 191340 154426
rect 191288 154362 191340 154368
rect 191012 153808 191064 153814
rect 191012 153750 191064 153756
rect 191104 153808 191156 153814
rect 191104 153750 191156 153756
rect 191300 153406 191328 154362
rect 191288 153400 191340 153406
rect 191288 153342 191340 153348
rect 191484 149954 191512 154974
rect 191668 152114 191696 159938
rect 191760 153406 191788 160006
rect 192128 157282 192156 163200
rect 192116 157276 192168 157282
rect 192116 157218 192168 157224
rect 192956 155854 192984 163200
rect 193784 159186 193812 163200
rect 193772 159180 193824 159186
rect 193772 159122 193824 159128
rect 194704 158982 194732 163200
rect 193404 158976 193456 158982
rect 193404 158918 193456 158924
rect 194692 158976 194744 158982
rect 194692 158918 194744 158924
rect 193220 157616 193272 157622
rect 193220 157558 193272 157564
rect 193232 157334 193260 157558
rect 193232 157306 193352 157334
rect 192944 155848 192996 155854
rect 192944 155790 192996 155796
rect 192114 153776 192170 153785
rect 192114 153711 192170 153720
rect 191748 153400 191800 153406
rect 191748 153342 191800 153348
rect 191656 152108 191708 152114
rect 191656 152050 191708 152056
rect 192128 149954 192156 153711
rect 192760 152924 192812 152930
rect 192760 152866 192812 152872
rect 192772 149954 192800 152866
rect 193324 149954 193352 157306
rect 193416 152182 193444 158918
rect 195428 158908 195480 158914
rect 195428 158850 195480 158856
rect 194692 156256 194744 156262
rect 194692 156198 194744 156204
rect 194048 155916 194100 155922
rect 194048 155858 194100 155864
rect 193404 152176 193456 152182
rect 193404 152118 193456 152124
rect 194060 149954 194088 155858
rect 194704 149954 194732 156198
rect 195440 152998 195468 158850
rect 195532 157826 195560 163200
rect 195520 157820 195572 157826
rect 195520 157762 195572 157768
rect 196164 156324 196216 156330
rect 196164 156266 196216 156272
rect 195428 152992 195480 152998
rect 195428 152934 195480 152940
rect 195336 151972 195388 151978
rect 195336 151914 195388 151920
rect 195348 149954 195376 151914
rect 196176 149954 196204 156266
rect 196360 155922 196388 163200
rect 197188 160070 197216 163200
rect 197176 160064 197228 160070
rect 197176 160006 197228 160012
rect 198016 160002 198044 163200
rect 198004 159996 198056 160002
rect 198004 159938 198056 159944
rect 197360 159112 197412 159118
rect 197360 159054 197412 159060
rect 197268 158840 197320 158846
rect 197268 158782 197320 158788
rect 196348 155916 196400 155922
rect 196348 155858 196400 155864
rect 197280 153898 197308 158782
rect 197372 157622 197400 159054
rect 198738 158536 198794 158545
rect 198738 158471 198794 158480
rect 197360 157616 197412 157622
rect 197360 157558 197412 157564
rect 198004 156256 198056 156262
rect 198004 156198 198056 156204
rect 198016 156058 198044 156198
rect 198004 156052 198056 156058
rect 198004 155994 198056 156000
rect 197280 153870 197492 153898
rect 197464 153814 197492 153870
rect 197360 153808 197412 153814
rect 197360 153750 197412 153756
rect 197452 153808 197504 153814
rect 197452 153750 197504 153756
rect 196624 153536 196676 153542
rect 196624 153478 196676 153484
rect 196636 149954 196664 153478
rect 197372 149954 197400 153750
rect 197912 153060 197964 153066
rect 197912 153002 197964 153008
rect 197924 149954 197952 153002
rect 198752 149954 198780 158471
rect 198844 156398 198872 163200
rect 198924 159316 198976 159322
rect 198924 159258 198976 159264
rect 198832 156392 198884 156398
rect 198832 156334 198884 156340
rect 198936 153542 198964 159258
rect 199672 155106 199700 163200
rect 200592 159050 200620 163200
rect 201420 159322 201448 163200
rect 201408 159316 201460 159322
rect 201408 159258 201460 159264
rect 200488 159044 200540 159050
rect 200488 158986 200540 158992
rect 200580 159044 200632 159050
rect 200580 158986 200632 158992
rect 200500 157334 200528 158986
rect 200500 157306 200620 157334
rect 199660 155100 199712 155106
rect 199660 155042 199712 155048
rect 200212 155032 200264 155038
rect 200212 154974 200264 154980
rect 199292 153808 199344 153814
rect 199292 153750 199344 153756
rect 198924 153536 198976 153542
rect 198924 153478 198976 153484
rect 199304 153474 199332 153750
rect 199200 153468 199252 153474
rect 199200 153410 199252 153416
rect 199292 153468 199344 153474
rect 199292 153410 199344 153416
rect 199212 149954 199240 153410
rect 200120 153400 200172 153406
rect 200118 153368 200120 153377
rect 200172 153368 200174 153377
rect 200118 153303 200174 153312
rect 200224 150090 200252 154974
rect 200488 153740 200540 153746
rect 200488 153682 200540 153688
rect 200500 153354 200528 153682
rect 200592 153474 200620 157306
rect 200764 156596 200816 156602
rect 200764 156538 200816 156544
rect 200948 156596 201000 156602
rect 200948 156538 201000 156544
rect 200776 156330 200804 156538
rect 200960 156398 200988 156538
rect 200948 156392 201000 156398
rect 200948 156334 201000 156340
rect 200764 156324 200816 156330
rect 200764 156266 200816 156272
rect 200672 156188 200724 156194
rect 200672 156130 200724 156136
rect 200580 153468 200632 153474
rect 200580 153410 200632 153416
rect 200316 153326 200528 153354
rect 200316 153270 200344 153326
rect 200304 153264 200356 153270
rect 200304 153206 200356 153212
rect 200488 152040 200540 152046
rect 200488 151982 200540 151988
rect 200224 150062 200344 150090
rect 181180 149926 181516 149954
rect 181824 149926 182160 149954
rect 182468 149926 182804 149954
rect 183020 149926 183448 149954
rect 183756 149926 184092 149954
rect 184400 149926 184736 149954
rect 185044 149926 185380 149954
rect 185596 149926 186024 149954
rect 186424 149926 186668 149954
rect 186976 149926 187312 149954
rect 187712 149926 187956 149954
rect 188172 149926 188600 149954
rect 189092 149926 189244 149954
rect 189552 149926 189888 149954
rect 190196 149926 190532 149954
rect 190748 149926 191176 149954
rect 191484 149926 191820 149954
rect 192128 149926 192464 149954
rect 192772 149926 193108 149954
rect 193324 149926 193752 149954
rect 194060 149926 194396 149954
rect 194704 149926 195040 149954
rect 195348 149926 195684 149954
rect 196176 149926 196328 149954
rect 196636 149926 196972 149954
rect 197372 149926 197616 149954
rect 197924 149926 198260 149954
rect 198752 149926 198904 149954
rect 199212 149926 199548 149954
rect 200316 149818 200344 150062
rect 200500 149954 200528 151982
rect 200684 150090 200712 156130
rect 202248 156058 202276 163200
rect 203076 156126 203104 163200
rect 203708 158976 203760 158982
rect 203708 158918 203760 158924
rect 203432 157548 203484 157554
rect 203432 157490 203484 157496
rect 203444 157334 203472 157490
rect 203444 157306 203656 157334
rect 203064 156120 203116 156126
rect 203064 156062 203116 156068
rect 202236 156052 202288 156058
rect 202236 155994 202288 156000
rect 202420 154488 202472 154494
rect 202420 154430 202472 154436
rect 201776 154420 201828 154426
rect 201776 154362 201828 154368
rect 200854 153368 200910 153377
rect 200854 153303 200856 153312
rect 200908 153303 200910 153312
rect 200856 153274 200908 153280
rect 200684 150062 201080 150090
rect 201052 149954 201080 150062
rect 201788 149954 201816 154362
rect 202432 149954 202460 154430
rect 203064 151904 203116 151910
rect 203064 151846 203116 151852
rect 203076 149954 203104 151846
rect 203628 149954 203656 157306
rect 203720 153066 203748 158918
rect 203904 158846 203932 163200
rect 204732 159361 204760 163200
rect 204718 159352 204774 159361
rect 204718 159287 204774 159296
rect 203892 158840 203944 158846
rect 203892 158782 203944 158788
rect 204904 158772 204956 158778
rect 204904 158714 204956 158720
rect 204916 157554 204944 158714
rect 204904 157548 204956 157554
rect 204904 157490 204956 157496
rect 204352 155780 204404 155786
rect 204352 155722 204404 155728
rect 203708 153060 203760 153066
rect 203708 153002 203760 153008
rect 204364 149954 204392 155722
rect 205008 154426 205036 163254
rect 205468 163146 205496 163254
rect 205546 163200 205602 164400
rect 206466 163200 206522 164400
rect 207294 163200 207350 164400
rect 208122 163200 208178 164400
rect 208412 163254 208900 163282
rect 205560 163146 205588 163200
rect 205468 163118 205588 163146
rect 206192 157480 206244 157486
rect 206192 157422 206244 157428
rect 204996 154420 205048 154426
rect 204996 154362 205048 154368
rect 205088 154352 205140 154358
rect 205088 154294 205140 154300
rect 205100 149954 205128 154294
rect 205640 153196 205692 153202
rect 205640 153138 205692 153144
rect 205652 149954 205680 153138
rect 206204 149954 206232 157422
rect 206480 155786 206508 163200
rect 207112 160064 207164 160070
rect 207112 160006 207164 160012
rect 207018 157176 207074 157185
rect 207018 157111 207074 157120
rect 206468 155780 206520 155786
rect 206468 155722 206520 155728
rect 207032 149954 207060 157111
rect 207124 155038 207152 160006
rect 207308 158982 207336 163200
rect 207296 158976 207348 158982
rect 207296 158918 207348 158924
rect 208136 158914 208164 163200
rect 208124 158908 208176 158914
rect 208124 158850 208176 158856
rect 207112 155032 207164 155038
rect 207112 154974 207164 154980
rect 208412 154358 208440 163254
rect 208872 163146 208900 163254
rect 208950 163200 209006 164400
rect 209778 163200 209834 164400
rect 210606 163200 210662 164400
rect 211434 163200 211490 164400
rect 211540 163254 212304 163282
rect 208964 163146 208992 163200
rect 208872 163118 208992 163146
rect 209792 156398 209820 163200
rect 210620 158778 210648 163200
rect 211448 160070 211476 163200
rect 211436 160064 211488 160070
rect 211436 160006 211488 160012
rect 210608 158772 210660 158778
rect 210608 158714 210660 158720
rect 209780 156392 209832 156398
rect 209780 156334 209832 156340
rect 211344 156256 211396 156262
rect 211344 156198 211396 156204
rect 208768 156188 208820 156194
rect 208768 156130 208820 156136
rect 208400 154352 208452 154358
rect 208400 154294 208452 154300
rect 207572 153264 207624 153270
rect 207572 153206 207624 153212
rect 207584 149954 207612 153206
rect 208400 152108 208452 152114
rect 208400 152050 208452 152056
rect 208412 149954 208440 152050
rect 208780 149954 208808 156130
rect 210148 153808 210200 153814
rect 210148 153750 210200 153756
rect 209780 153740 209832 153746
rect 209780 153682 209832 153688
rect 209792 150226 209820 153682
rect 209792 150198 209866 150226
rect 200500 149926 200836 149954
rect 201052 149926 201480 149954
rect 201788 149926 202124 149954
rect 202432 149926 202768 149954
rect 203076 149926 203412 149954
rect 203628 149926 204056 149954
rect 204364 149926 204700 149954
rect 205100 149926 205344 149954
rect 205652 149926 205988 149954
rect 206204 149926 206632 149954
rect 207032 149926 207276 149954
rect 207584 149926 207920 149954
rect 208412 149926 208564 149954
rect 208780 149926 209208 149954
rect 209838 149940 209866 150198
rect 210160 149954 210188 153750
rect 210792 152380 210844 152386
rect 210792 152322 210844 152328
rect 210804 149954 210832 152322
rect 211356 149954 211384 156198
rect 211540 153785 211568 163254
rect 212276 163146 212304 163254
rect 212354 163200 212410 164400
rect 213182 163200 213238 164400
rect 214010 163200 214066 164400
rect 214838 163200 214894 164400
rect 215312 163254 215616 163282
rect 212368 163146 212396 163200
rect 212276 163118 212396 163146
rect 212632 159316 212684 159322
rect 212632 159258 212684 159264
rect 212448 158908 212500 158914
rect 212448 158850 212500 158856
rect 211988 154964 212040 154970
rect 211988 154906 212040 154912
rect 211526 153776 211582 153785
rect 211526 153711 211582 153720
rect 212000 149954 212028 154906
rect 212460 152930 212488 158850
rect 212448 152924 212500 152930
rect 212448 152866 212500 152872
rect 212644 152046 212672 159258
rect 213196 156330 213224 163200
rect 214024 159322 214052 163200
rect 214012 159316 214064 159322
rect 214012 159258 214064 159264
rect 214656 159248 214708 159254
rect 214656 159190 214708 159196
rect 213644 158840 213696 158846
rect 213644 158782 213696 158788
rect 213184 156324 213236 156330
rect 213184 156266 213236 156272
rect 212724 154556 212776 154562
rect 212724 154498 212776 154504
rect 212632 152040 212684 152046
rect 212632 151982 212684 151988
rect 212736 149954 212764 154498
rect 213276 152176 213328 152182
rect 213276 152118 213328 152124
rect 213288 149954 213316 152118
rect 213656 152114 213684 158782
rect 214472 157344 214524 157350
rect 214472 157286 214524 157292
rect 214564 157344 214616 157350
rect 214564 157286 214616 157292
rect 213920 156664 213972 156670
rect 213920 156606 213972 156612
rect 213644 152108 213696 152114
rect 213644 152050 213696 152056
rect 213932 149954 213960 156606
rect 214484 156262 214512 157286
rect 214576 156942 214604 157286
rect 214564 156936 214616 156942
rect 214564 156878 214616 156884
rect 214472 156256 214524 156262
rect 214472 156198 214524 156204
rect 214472 155236 214524 155242
rect 214472 155178 214524 155184
rect 214484 149954 214512 155178
rect 214668 154970 214696 159190
rect 214852 158846 214880 163200
rect 214840 158840 214892 158846
rect 214840 158782 214892 158788
rect 214656 154964 214708 154970
rect 214656 154906 214708 154912
rect 215312 154494 215340 163254
rect 215588 163146 215616 163254
rect 215666 163200 215722 164400
rect 216494 163200 216550 164400
rect 217322 163200 217378 164400
rect 218242 163200 218298 164400
rect 218348 163254 219020 163282
rect 215680 163146 215708 163200
rect 215588 163118 215708 163146
rect 215392 158772 215444 158778
rect 215392 158714 215444 158720
rect 215300 154488 215352 154494
rect 215300 154430 215352 154436
rect 215404 153202 215432 158714
rect 216508 156670 216536 163200
rect 217336 158914 217364 163200
rect 218256 159254 218284 163200
rect 218244 159248 218296 159254
rect 218244 159190 218296 159196
rect 218060 159180 218112 159186
rect 218060 159122 218112 159128
rect 217324 158908 217376 158914
rect 217324 158850 217376 158856
rect 216680 156732 216732 156738
rect 216680 156674 216732 156680
rect 216496 156664 216548 156670
rect 216496 156606 216548 156612
rect 215484 156188 215536 156194
rect 215484 156130 215536 156136
rect 215392 153196 215444 153202
rect 215392 153138 215444 153144
rect 215496 150226 215524 156130
rect 215852 152516 215904 152522
rect 215852 152458 215904 152464
rect 215496 150198 215570 150226
rect 210160 149926 210496 149954
rect 210804 149926 211140 149954
rect 211356 149926 211692 149954
rect 212000 149926 212336 149954
rect 212736 149926 212980 149954
rect 213288 149926 213624 149954
rect 213932 149926 214268 149954
rect 214484 149926 214912 149954
rect 215542 149940 215570 150198
rect 215864 149954 215892 152458
rect 216692 149954 216720 156674
rect 218072 156194 218100 159122
rect 218060 156188 218112 156194
rect 218060 156130 218112 156136
rect 217048 155304 217100 155310
rect 217048 155246 217100 155252
rect 217060 149954 217088 155246
rect 218348 154562 218376 163254
rect 218992 163146 219020 163254
rect 219070 163200 219126 164400
rect 219898 163200 219954 164400
rect 220726 163200 220782 164400
rect 221554 163200 221610 164400
rect 222382 163200 222438 164400
rect 223210 163200 223266 164400
rect 224130 163200 224186 164400
rect 224958 163200 225014 164400
rect 225064 163254 225736 163282
rect 219084 163146 219112 163200
rect 218992 163118 219112 163146
rect 219912 161474 219940 163200
rect 219912 161446 220124 161474
rect 218980 158024 219032 158030
rect 218980 157966 219032 157972
rect 218336 154556 218388 154562
rect 218336 154498 218388 154504
rect 218060 153672 218112 153678
rect 218060 153614 218112 153620
rect 218072 150226 218100 153614
rect 218428 152992 218480 152998
rect 218428 152934 218480 152940
rect 218072 150198 218146 150226
rect 215864 149926 216200 149954
rect 216692 149926 216844 149954
rect 217060 149926 217488 149954
rect 218118 149940 218146 150198
rect 218440 149954 218468 152934
rect 218992 149954 219020 157966
rect 220096 156262 220124 161446
rect 220740 159186 220768 163200
rect 220728 159180 220780 159186
rect 220728 159122 220780 159128
rect 220728 158908 220780 158914
rect 220728 158850 220780 158856
rect 219992 156256 220044 156262
rect 219992 156198 220044 156204
rect 220084 156256 220136 156262
rect 220084 156198 220136 156204
rect 219716 154012 219768 154018
rect 219716 153954 219768 153960
rect 219728 149954 219756 153954
rect 220004 151814 220032 156198
rect 220740 152522 220768 158850
rect 221568 158778 221596 163200
rect 222396 161474 222424 163200
rect 222396 161446 222516 161474
rect 222108 158840 222160 158846
rect 222108 158782 222160 158788
rect 221556 158772 221608 158778
rect 221556 158714 221608 158720
rect 221372 157344 221424 157350
rect 221372 157286 221424 157292
rect 220728 152516 220780 152522
rect 220728 152458 220780 152464
rect 221004 152244 221056 152250
rect 221004 152186 221056 152192
rect 220004 151786 220308 151814
rect 220280 149954 220308 151786
rect 221016 149954 221044 152186
rect 221384 151814 221412 157286
rect 222120 152250 222148 158782
rect 222384 156868 222436 156874
rect 222384 156810 222436 156816
rect 222108 152244 222160 152250
rect 222108 152186 222160 152192
rect 221384 151786 221596 151814
rect 221568 149954 221596 151786
rect 222396 149954 222424 156810
rect 222488 154018 222516 161446
rect 223224 156738 223252 163200
rect 223580 159384 223632 159390
rect 223580 159326 223632 159332
rect 223212 156732 223264 156738
rect 223212 156674 223264 156680
rect 222476 154012 222528 154018
rect 222476 153954 222528 153960
rect 222936 153944 222988 153950
rect 222936 153886 222988 153892
rect 222948 149954 222976 153886
rect 223592 149954 223620 159326
rect 224144 159118 224172 163200
rect 224972 159390 225000 163200
rect 224960 159384 225012 159390
rect 224960 159326 225012 159332
rect 224132 159112 224184 159118
rect 224132 159054 224184 159060
rect 224960 159044 225012 159050
rect 224960 158986 225012 158992
rect 224040 158772 224092 158778
rect 224040 158714 224092 158720
rect 224052 152386 224080 158714
rect 224224 157344 224276 157350
rect 224224 157286 224276 157292
rect 224132 157004 224184 157010
rect 224132 156946 224184 156952
rect 224040 152380 224092 152386
rect 224040 152322 224092 152328
rect 224144 149954 224172 156946
rect 224236 156330 224264 157286
rect 224972 156942 225000 158986
rect 224960 156936 225012 156942
rect 224960 156878 225012 156884
rect 224224 156324 224276 156330
rect 224224 156266 224276 156272
rect 225064 153950 225092 163254
rect 225708 163146 225736 163254
rect 225786 163200 225842 164400
rect 226614 163200 226670 164400
rect 226812 163254 227392 163282
rect 225800 163146 225828 163200
rect 225708 163118 225828 163146
rect 225236 159520 225288 159526
rect 225236 159462 225288 159468
rect 225144 156800 225196 156806
rect 225144 156742 225196 156748
rect 225052 153944 225104 153950
rect 225052 153886 225104 153892
rect 225156 150226 225184 156742
rect 225248 152998 225276 159462
rect 226628 156874 226656 163200
rect 226708 157412 226760 157418
rect 226708 157354 226760 157360
rect 226616 156868 226668 156874
rect 226616 156810 226668 156816
rect 225512 156528 225564 156534
rect 225512 156470 225564 156476
rect 225236 152992 225288 152998
rect 225236 152934 225288 152940
rect 225156 150198 225230 150226
rect 218440 149926 218776 149954
rect 218992 149926 219420 149954
rect 219728 149926 220064 149954
rect 220280 149926 220708 149954
rect 221016 149926 221352 149954
rect 221568 149926 221996 149954
rect 222396 149926 222640 149954
rect 222948 149926 223284 149954
rect 223592 149926 223928 149954
rect 224144 149926 224572 149954
rect 225202 149940 225230 150198
rect 225524 149954 225552 156470
rect 226340 152584 226392 152590
rect 226340 152526 226392 152532
rect 226352 149954 226380 152526
rect 226720 149954 226748 157354
rect 226812 152425 226840 163254
rect 227364 163146 227392 163254
rect 227442 163200 227498 164400
rect 227732 163254 228220 163282
rect 227456 163146 227484 163200
rect 227364 163118 227484 163146
rect 227732 152522 227760 163254
rect 228192 163146 228220 163254
rect 228270 163200 228326 164400
rect 229098 163200 229154 164400
rect 230018 163200 230074 164400
rect 230846 163200 230902 164400
rect 231674 163200 231730 164400
rect 231872 163254 232452 163282
rect 228284 163146 228312 163200
rect 228192 163118 228312 163146
rect 228088 156460 228140 156466
rect 228088 156402 228140 156408
rect 227904 155372 227956 155378
rect 227904 155314 227956 155320
rect 227720 152516 227772 152522
rect 227720 152458 227772 152464
rect 226798 152416 226854 152425
rect 226798 152351 226854 152360
rect 227916 149954 227944 155314
rect 225524 149926 225860 149954
rect 226352 149926 226504 149954
rect 226720 149926 227148 149954
rect 227792 149926 227944 149954
rect 228100 149954 228128 156402
rect 229112 153678 229140 163200
rect 230032 156806 230060 163200
rect 230860 159050 230888 163200
rect 231688 159526 231716 163200
rect 231676 159520 231728 159526
rect 231676 159462 231728 159468
rect 230848 159044 230900 159050
rect 230848 158986 230900 158992
rect 230756 158976 230808 158982
rect 230756 158918 230808 158924
rect 230020 156800 230072 156806
rect 230020 156742 230072 156748
rect 230768 156194 230796 158918
rect 230756 156188 230808 156194
rect 230756 156130 230808 156136
rect 229284 155984 229336 155990
rect 229284 155926 229336 155932
rect 229100 153672 229152 153678
rect 229100 153614 229152 153620
rect 228732 152992 228784 152998
rect 228732 152934 228784 152940
rect 228824 152992 228876 152998
rect 228824 152934 228876 152940
rect 228744 149954 228772 152934
rect 228836 152590 228864 152934
rect 228824 152584 228876 152590
rect 228824 152526 228876 152532
rect 229296 149954 229324 155926
rect 230020 155440 230072 155446
rect 230020 155382 230072 155388
rect 230032 149954 230060 155382
rect 231872 153814 231900 163254
rect 232424 163146 232452 163254
rect 232502 163200 232558 164400
rect 233330 163200 233386 164400
rect 234158 163200 234214 164400
rect 234986 163200 235042 164400
rect 235092 163254 235856 163282
rect 232516 163146 232544 163200
rect 232424 163118 232544 163146
rect 231952 158092 232004 158098
rect 231952 158034 232004 158040
rect 231860 153808 231912 153814
rect 231860 153750 231912 153756
rect 230664 153604 230716 153610
rect 230664 153546 230716 153552
rect 230676 149954 230704 153546
rect 231308 152720 231360 152726
rect 231308 152662 231360 152668
rect 231320 149954 231348 152662
rect 231964 149954 231992 158034
rect 233344 155310 233372 163200
rect 233884 159452 233936 159458
rect 233884 159394 233936 159400
rect 233516 157208 233568 157214
rect 233516 157150 233568 157156
rect 233332 155304 233384 155310
rect 233332 155246 233384 155252
rect 232504 154828 232556 154834
rect 232504 154770 232556 154776
rect 232516 149954 232544 154770
rect 233528 150226 233556 157150
rect 233528 150198 233602 150226
rect 228100 149926 228436 149954
rect 228744 149926 229080 149954
rect 229296 149926 229724 149954
rect 230032 149926 230368 149954
rect 230676 149926 231012 149954
rect 231320 149926 231656 149954
rect 231964 149926 232300 149954
rect 232516 149926 232944 149954
rect 233574 149940 233602 150198
rect 233896 149954 233924 159394
rect 234172 152590 234200 163200
rect 235000 159458 235028 163200
rect 234988 159452 235040 159458
rect 234988 159394 235040 159400
rect 234804 157072 234856 157078
rect 234804 157014 234856 157020
rect 234160 152584 234212 152590
rect 234160 152526 234212 152532
rect 234816 150226 234844 157014
rect 235092 153746 235120 163254
rect 235828 163146 235856 163254
rect 235906 163200 235962 164400
rect 236734 163200 236790 164400
rect 237562 163200 237618 164400
rect 238390 163200 238446 164400
rect 238864 163254 239168 163282
rect 235920 163146 235948 163200
rect 235828 163118 235948 163146
rect 236748 158030 236776 163200
rect 237576 158982 237604 163200
rect 237564 158976 237616 158982
rect 237564 158918 237616 158924
rect 238404 158846 238432 163200
rect 238392 158840 238444 158846
rect 238392 158782 238444 158788
rect 237380 158160 237432 158166
rect 237380 158102 237432 158108
rect 236736 158024 236788 158030
rect 236736 157966 236788 157972
rect 236092 157684 236144 157690
rect 236092 157626 236144 157632
rect 235172 153876 235224 153882
rect 235172 153818 235224 153824
rect 235080 153740 235132 153746
rect 235080 153682 235132 153688
rect 234816 150198 234890 150226
rect 233896 149926 234232 149954
rect 234862 149940 234890 150198
rect 235184 149954 235212 153818
rect 236104 150226 236132 157626
rect 236460 152652 236512 152658
rect 236460 152594 236512 152600
rect 236104 150198 236178 150226
rect 235184 149926 235520 149954
rect 236150 149940 236178 150198
rect 236472 149954 236500 152594
rect 237392 150226 237420 158102
rect 237656 154760 237708 154766
rect 237656 154702 237708 154708
rect 237392 150198 237466 150226
rect 236472 149926 236808 149954
rect 237438 149940 237466 150198
rect 237668 149954 237696 154702
rect 238864 153610 238892 163254
rect 239140 163146 239168 163254
rect 239218 163200 239274 164400
rect 240046 163200 240102 164400
rect 240874 163200 240930 164400
rect 241794 163200 241850 164400
rect 241900 163254 242572 163282
rect 239232 163146 239260 163200
rect 239140 163118 239260 163146
rect 239128 159588 239180 159594
rect 239128 159530 239180 159536
rect 238852 153604 238904 153610
rect 238852 153546 238904 153552
rect 238392 153332 238444 153338
rect 238392 153274 238444 153280
rect 238404 149954 238432 153274
rect 239140 149954 239168 159530
rect 239680 158228 239732 158234
rect 239680 158170 239732 158176
rect 239692 149954 239720 158170
rect 240060 155242 240088 163200
rect 240888 158778 240916 163200
rect 241428 159656 241480 159662
rect 241428 159598 241480 159604
rect 240876 158772 240928 158778
rect 240876 158714 240928 158720
rect 240048 155236 240100 155242
rect 240048 155178 240100 155184
rect 240232 154624 240284 154630
rect 240232 154566 240284 154572
rect 240244 149954 240272 154566
rect 240968 154080 241020 154086
rect 240968 154022 241020 154028
rect 240980 149954 241008 154022
rect 241440 151814 241468 159598
rect 241808 158914 241836 163200
rect 241796 158908 241848 158914
rect 241796 158850 241848 158856
rect 241612 158840 241664 158846
rect 241612 158782 241664 158788
rect 241624 151978 241652 158782
rect 241900 153882 241928 163254
rect 242544 163146 242572 163254
rect 242622 163200 242678 164400
rect 243450 163200 243506 164400
rect 244278 163200 244334 164400
rect 244384 163254 245056 163282
rect 242636 163146 242664 163200
rect 242544 163118 242664 163146
rect 243360 158772 243412 158778
rect 243360 158714 243412 158720
rect 242072 158296 242124 158302
rect 242072 158238 242124 158244
rect 241888 153876 241940 153882
rect 241888 153818 241940 153824
rect 241612 151972 241664 151978
rect 241612 151914 241664 151920
rect 241440 151786 241560 151814
rect 241532 149954 241560 151786
rect 242084 149954 242112 158238
rect 242900 154692 242952 154698
rect 242900 154634 242952 154640
rect 242912 149954 242940 154634
rect 243372 151910 243400 158714
rect 243464 158098 243492 163200
rect 244292 159662 244320 163200
rect 244280 159656 244332 159662
rect 244280 159598 244332 159604
rect 243452 158092 243504 158098
rect 243452 158034 243504 158040
rect 243452 153400 243504 153406
rect 243452 153342 243504 153348
rect 243360 151904 243412 151910
rect 243360 151846 243412 151852
rect 243464 149954 243492 153342
rect 244280 152788 244332 152794
rect 244280 152730 244332 152736
rect 244292 149954 244320 152730
rect 244384 152182 244412 163254
rect 245028 163146 245056 163254
rect 245106 163200 245162 164400
rect 245934 163200 245990 164400
rect 246762 163200 246818 164400
rect 247052 163254 247632 163282
rect 245120 163146 245148 163200
rect 245028 163118 245148 163146
rect 244648 158432 244700 158438
rect 244648 158374 244700 158380
rect 244372 152176 244424 152182
rect 244372 152118 244424 152124
rect 244660 149954 244688 158374
rect 245844 154896 245896 154902
rect 245844 154838 245896 154844
rect 245660 154148 245712 154154
rect 245660 154090 245712 154096
rect 245672 150226 245700 154090
rect 245856 151814 245884 154838
rect 245948 154154 245976 163200
rect 246580 159724 246632 159730
rect 246580 159666 246632 159672
rect 245936 154148 245988 154154
rect 245936 154090 245988 154096
rect 245856 151786 245976 151814
rect 245672 150198 245746 150226
rect 237668 149926 238096 149954
rect 238404 149926 238740 149954
rect 239140 149926 239384 149954
rect 239692 149926 240028 149954
rect 240244 149926 240672 149954
rect 240980 149926 241316 149954
rect 241532 149926 241960 149954
rect 242084 149926 242512 149954
rect 242912 149926 243156 149954
rect 243464 149926 243800 149954
rect 244292 149926 244444 149954
rect 244660 149926 245088 149954
rect 245718 149940 245746 150198
rect 245948 149954 245976 151786
rect 246592 149954 246620 159666
rect 246776 158166 246804 163200
rect 246764 158160 246816 158166
rect 246764 158102 246816 158108
rect 247052 152658 247080 163254
rect 247604 163146 247632 163254
rect 247682 163200 247738 164400
rect 248510 163200 248566 164400
rect 248616 163254 249288 163282
rect 247696 163146 247724 163200
rect 247604 163118 247724 163146
rect 248524 159730 248552 163200
rect 248512 159724 248564 159730
rect 248512 159666 248564 159672
rect 247132 158364 247184 158370
rect 247132 158306 247184 158312
rect 247040 152652 247092 152658
rect 247040 152594 247092 152600
rect 247144 151814 247172 158306
rect 247868 155508 247920 155514
rect 247868 155450 247920 155456
rect 247144 151786 247264 151814
rect 247236 149954 247264 151786
rect 247880 149954 247908 155450
rect 248616 154086 248644 163254
rect 249260 163146 249288 163254
rect 249338 163200 249394 164400
rect 250166 163200 250222 164400
rect 250994 163200 251050 164400
rect 251192 163254 251772 163282
rect 249352 163146 249380 163200
rect 249260 163118 249380 163146
rect 249800 158636 249852 158642
rect 249800 158578 249852 158584
rect 248604 154080 248656 154086
rect 248604 154022 248656 154028
rect 248604 153536 248656 153542
rect 248604 153478 248656 153484
rect 248616 149954 248644 153478
rect 249248 152448 249300 152454
rect 249248 152390 249300 152396
rect 249260 149954 249288 152390
rect 249812 149954 249840 158578
rect 250180 155378 250208 163200
rect 251008 159594 251036 163200
rect 250996 159588 251048 159594
rect 250996 159530 251048 159536
rect 250168 155372 250220 155378
rect 250168 155314 250220 155320
rect 250536 154216 250588 154222
rect 250536 154158 250588 154164
rect 250548 149954 250576 154158
rect 251192 152726 251220 163254
rect 251744 163146 251772 163254
rect 251822 163200 251878 164400
rect 252650 163200 252706 164400
rect 253570 163200 253626 164400
rect 254398 163200 254454 164400
rect 255226 163200 255282 164400
rect 255332 163254 256004 163282
rect 251836 163146 251864 163200
rect 251744 163118 251864 163146
rect 252560 158500 252612 158506
rect 252560 158442 252612 158448
rect 251272 157616 251324 157622
rect 251272 157558 251324 157564
rect 251180 152720 251232 152726
rect 251180 152662 251232 152668
rect 251284 149954 251312 157558
rect 251824 152856 251876 152862
rect 251824 152798 251876 152804
rect 251836 149954 251864 152798
rect 252572 149954 252600 158442
rect 252664 153542 252692 163200
rect 253020 155644 253072 155650
rect 253020 155586 253072 155592
rect 252652 153536 252704 153542
rect 252652 153478 252704 153484
rect 253032 149954 253060 155586
rect 253584 155446 253612 163200
rect 254308 159792 254360 159798
rect 254308 159734 254360 159740
rect 254032 157140 254084 157146
rect 254032 157082 254084 157088
rect 253572 155440 253624 155446
rect 253572 155382 253624 155388
rect 254044 150226 254072 157082
rect 254044 150198 254118 150226
rect 245948 149926 246376 149954
rect 246592 149926 247020 149954
rect 247236 149926 247664 149954
rect 247880 149926 248308 149954
rect 248616 149926 248952 149954
rect 249260 149926 249596 149954
rect 249812 149926 250240 149954
rect 250548 149926 250884 149954
rect 251284 149926 251528 149954
rect 251836 149926 252172 149954
rect 252572 149926 252816 149954
rect 253032 149926 253460 149954
rect 254090 149940 254118 150198
rect 254320 149954 254348 159734
rect 254412 158778 254440 163200
rect 255240 159798 255268 163200
rect 255228 159792 255280 159798
rect 255228 159734 255280 159740
rect 254400 158772 254452 158778
rect 254400 158714 254452 158720
rect 255332 154222 255360 163254
rect 255976 163146 256004 163254
rect 256054 163200 256110 164400
rect 256882 163200 256938 164400
rect 257710 163200 257766 164400
rect 258538 163200 258594 164400
rect 259458 163200 259514 164400
rect 260286 163200 260342 164400
rect 261114 163200 261170 164400
rect 261942 163200 261998 164400
rect 262232 163254 262720 163282
rect 256068 163146 256096 163200
rect 255976 163118 256096 163146
rect 255412 158772 255464 158778
rect 255412 158714 255464 158720
rect 255320 154216 255372 154222
rect 255320 154158 255372 154164
rect 255424 152862 255452 158714
rect 255596 158568 255648 158574
rect 255596 158510 255648 158516
rect 255412 152856 255464 152862
rect 255412 152798 255464 152804
rect 255608 149954 255636 158510
rect 256896 158234 256924 163200
rect 257528 158704 257580 158710
rect 257528 158646 257580 158652
rect 256884 158228 256936 158234
rect 256884 158170 256936 158176
rect 255872 157548 255924 157554
rect 255872 157490 255924 157496
rect 255688 155576 255740 155582
rect 255688 155518 255740 155524
rect 254320 149926 254748 149954
rect 255392 149926 255636 149954
rect 255700 149954 255728 155518
rect 255884 151814 255912 157490
rect 256976 153128 257028 153134
rect 256976 153070 257028 153076
rect 255884 151786 256280 151814
rect 256252 149954 256280 151786
rect 256988 149954 257016 153070
rect 257540 149954 257568 158646
rect 257724 152794 257752 163200
rect 258552 158778 258580 163200
rect 258540 158772 258592 158778
rect 258540 158714 258592 158720
rect 258264 154284 258316 154290
rect 258264 154226 258316 154232
rect 257712 152788 257764 152794
rect 257712 152730 257764 152736
rect 258276 149954 258304 154226
rect 258908 153468 258960 153474
rect 258908 153410 258960 153416
rect 258920 149954 258948 153410
rect 259472 153406 259500 163200
rect 259552 159860 259604 159866
rect 259552 159802 259604 159808
rect 259460 153400 259512 153406
rect 259460 153342 259512 153348
rect 259564 149954 259592 159802
rect 260104 157956 260156 157962
rect 260104 157898 260156 157904
rect 260116 149954 260144 157898
rect 260300 155514 260328 163200
rect 261128 158846 261156 163200
rect 261956 159866 261984 163200
rect 261944 159860 261996 159866
rect 261944 159802 261996 159808
rect 261116 158840 261168 158846
rect 261116 158782 261168 158788
rect 260840 158772 260892 158778
rect 260840 158714 260892 158720
rect 260288 155508 260340 155514
rect 260288 155450 260340 155456
rect 260852 152454 260880 158714
rect 260932 155712 260984 155718
rect 260932 155654 260984 155660
rect 260840 152448 260892 152454
rect 260840 152390 260892 152396
rect 260944 149954 260972 155654
rect 261484 154964 261536 154970
rect 261484 154906 261536 154912
rect 261496 149954 261524 154906
rect 262232 154290 262260 163254
rect 262692 163146 262720 163254
rect 262770 163200 262826 164400
rect 263598 163200 263654 164400
rect 264426 163200 264482 164400
rect 264992 163254 265296 163282
rect 262784 163146 262812 163200
rect 262692 163118 262812 163146
rect 262680 157888 262732 157894
rect 262680 157830 262732 157836
rect 262220 154284 262272 154290
rect 262220 154226 262272 154232
rect 262220 152312 262272 152318
rect 262220 152254 262272 152260
rect 262232 149954 262260 152254
rect 262692 149954 262720 157830
rect 263612 155582 263640 163200
rect 264440 158778 264468 163200
rect 264888 159928 264940 159934
rect 264888 159870 264940 159876
rect 264428 158772 264480 158778
rect 264428 158714 264480 158720
rect 264060 157752 264112 157758
rect 264060 157694 264112 157700
rect 263600 155576 263652 155582
rect 263600 155518 263652 155524
rect 263692 155168 263744 155174
rect 263692 155110 263744 155116
rect 263704 150226 263732 155110
rect 263704 150198 263778 150226
rect 255700 149926 256036 149954
rect 256252 149926 256680 149954
rect 256988 149926 257324 149954
rect 257540 149926 257968 149954
rect 258276 149926 258612 149954
rect 258920 149926 259256 149954
rect 259564 149926 259900 149954
rect 260116 149926 260544 149954
rect 260944 149926 261188 149954
rect 261496 149926 261832 149954
rect 262232 149926 262476 149954
rect 262692 149926 263120 149954
rect 263750 149940 263778 150198
rect 264072 149954 264100 157694
rect 264900 151814 264928 159870
rect 264992 153134 265020 163254
rect 265268 163146 265296 163254
rect 265346 163200 265402 164400
rect 265452 163254 266124 163282
rect 265360 163146 265388 163200
rect 265268 163118 265388 163146
rect 265164 157276 265216 157282
rect 265164 157218 265216 157224
rect 264980 153128 265032 153134
rect 264980 153070 265032 153076
rect 265176 151814 265204 157218
rect 265452 153474 265480 163254
rect 266096 163146 266124 163254
rect 266174 163200 266230 164400
rect 267002 163200 267058 164400
rect 267830 163200 267886 164400
rect 268658 163200 268714 164400
rect 269224 163254 269436 163282
rect 266188 163146 266216 163200
rect 266096 163118 266216 163146
rect 266360 158772 266412 158778
rect 266360 158714 266412 158720
rect 265900 155848 265952 155854
rect 265900 155790 265952 155796
rect 265440 153468 265492 153474
rect 265440 153410 265492 153416
rect 264900 151786 265020 151814
rect 265176 151786 265296 151814
rect 264992 150226 265020 151786
rect 264992 150198 265066 150226
rect 264072 149926 264408 149954
rect 265038 149940 265066 150198
rect 265268 149954 265296 151786
rect 265912 149954 265940 155790
rect 266372 152318 266400 158714
rect 266544 156256 266596 156262
rect 266544 156198 266596 156204
rect 266360 152312 266412 152318
rect 266360 152254 266412 152260
rect 266556 149954 266584 156198
rect 267016 155650 267044 163200
rect 267844 158778 267872 163200
rect 268672 159934 268700 163200
rect 268660 159928 268712 159934
rect 268660 159870 268712 159876
rect 267832 158772 267884 158778
rect 267832 158714 267884 158720
rect 267740 157820 267792 157826
rect 267740 157762 267792 157768
rect 267004 155644 267056 155650
rect 267004 155586 267056 155592
rect 267280 153060 267332 153066
rect 267280 153002 267332 153008
rect 267292 149954 267320 153002
rect 267752 151814 267780 157762
rect 268476 155916 268528 155922
rect 268476 155858 268528 155864
rect 267752 151786 267872 151814
rect 267844 149954 267872 151786
rect 268488 149954 268516 155858
rect 269224 153270 269252 163254
rect 269408 163146 269436 163254
rect 269486 163200 269542 164400
rect 270314 163200 270370 164400
rect 271234 163200 271290 164400
rect 272062 163200 272118 164400
rect 272890 163200 272946 164400
rect 273718 163200 273774 164400
rect 274546 163200 274602 164400
rect 275374 163200 275430 164400
rect 276202 163200 276258 164400
rect 277122 163200 277178 164400
rect 277412 163254 277900 163282
rect 269500 163146 269528 163200
rect 269408 163118 269528 163146
rect 269856 159996 269908 160002
rect 269856 159938 269908 159944
rect 269304 155032 269356 155038
rect 269304 154974 269356 154980
rect 269212 153264 269264 153270
rect 269212 153206 269264 153212
rect 269316 149954 269344 154974
rect 269868 149954 269896 159938
rect 270328 155718 270356 163200
rect 271248 160002 271276 163200
rect 272076 161474 272104 163200
rect 272076 161446 272196 161474
rect 271236 159996 271288 160002
rect 271236 159938 271288 159944
rect 272064 156936 272116 156942
rect 272064 156878 272116 156884
rect 270500 156596 270552 156602
rect 270500 156538 270552 156544
rect 270316 155712 270368 155718
rect 270316 155654 270368 155660
rect 270512 149954 270540 156538
rect 271052 155100 271104 155106
rect 271052 155042 271104 155048
rect 271064 149954 271092 155042
rect 272076 150226 272104 156878
rect 272168 153066 272196 161446
rect 272524 159996 272576 160002
rect 272524 159938 272576 159944
rect 272156 153060 272208 153066
rect 272156 153002 272208 153008
rect 272536 152046 272564 159938
rect 272904 153338 272932 163200
rect 273732 157010 273760 163200
rect 274560 159497 274588 163200
rect 275388 160002 275416 163200
rect 275376 159996 275428 160002
rect 275376 159938 275428 159944
rect 274546 159488 274602 159497
rect 274546 159423 274602 159432
rect 274822 159352 274878 159361
rect 274822 159287 274878 159296
rect 273720 157004 273772 157010
rect 273720 156946 273772 156952
rect 273536 156120 273588 156126
rect 273536 156062 273588 156068
rect 273352 156052 273404 156058
rect 273352 155994 273404 156000
rect 272892 153332 272944 153338
rect 272892 153274 272944 153280
rect 272432 152040 272484 152046
rect 272432 151982 272484 151988
rect 272524 152040 272576 152046
rect 272524 151982 272576 151988
rect 272076 150198 272150 150226
rect 265268 149926 265696 149954
rect 265912 149926 266340 149954
rect 266556 149926 266984 149954
rect 267292 149926 267628 149954
rect 267844 149926 268272 149954
rect 268488 149926 268916 149954
rect 269316 149926 269560 149954
rect 269868 149926 270204 149954
rect 270512 149926 270848 149954
rect 271064 149926 271492 149954
rect 272122 149940 272150 150198
rect 272444 149954 272472 151982
rect 273364 150226 273392 155994
rect 273318 150198 273392 150226
rect 272444 149926 272780 149954
rect 273318 149940 273346 150198
rect 273548 149954 273576 156062
rect 274272 152108 274324 152114
rect 274272 152050 274324 152056
rect 274284 149954 274312 152050
rect 274836 149954 274864 159287
rect 276112 155780 276164 155786
rect 276112 155722 276164 155728
rect 275560 154420 275612 154426
rect 275560 154362 275612 154368
rect 275572 149954 275600 154362
rect 276124 149954 276152 155722
rect 276216 154426 276244 163200
rect 277136 156942 277164 163200
rect 277124 156936 277176 156942
rect 277124 156878 277176 156884
rect 276756 156188 276808 156194
rect 276756 156130 276808 156136
rect 276204 154420 276256 154426
rect 276204 154362 276256 154368
rect 276768 149954 276796 156130
rect 277412 152114 277440 163254
rect 277872 163146 277900 163254
rect 277950 163200 278006 164400
rect 278778 163200 278834 164400
rect 278884 163254 279556 163282
rect 277964 163146 277992 163200
rect 277872 163118 277992 163146
rect 278136 154352 278188 154358
rect 278136 154294 278188 154300
rect 277492 152924 277544 152930
rect 277492 152866 277544 152872
rect 277400 152108 277452 152114
rect 277400 152050 277452 152056
rect 277504 149954 277532 152866
rect 278148 149954 278176 154294
rect 278792 152930 278820 163200
rect 278884 154358 278912 163254
rect 279528 163146 279556 163254
rect 279606 163200 279662 164400
rect 280434 163200 280490 164400
rect 281262 163200 281318 164400
rect 282090 163200 282146 164400
rect 283010 163200 283066 164400
rect 283116 163254 283420 163282
rect 279620 163146 279648 163200
rect 279528 163118 279648 163146
rect 280160 160064 280212 160070
rect 280160 160006 280212 160012
rect 278964 156392 279016 156398
rect 278964 156334 279016 156340
rect 278872 154352 278924 154358
rect 278872 154294 278924 154300
rect 278780 152924 278832 152930
rect 278780 152866 278832 152872
rect 278976 149954 279004 156334
rect 279424 153196 279476 153202
rect 279424 153138 279476 153144
rect 279436 149954 279464 153138
rect 280172 149954 280200 160006
rect 280448 157078 280476 163200
rect 281276 160070 281304 163200
rect 281264 160064 281316 160070
rect 281264 160006 281316 160012
rect 282104 159322 282132 163200
rect 283024 163146 283052 163200
rect 283116 163146 283144 163254
rect 283024 163118 283144 163146
rect 282000 159316 282052 159322
rect 282000 159258 282052 159264
rect 282092 159316 282144 159322
rect 282092 159258 282144 159264
rect 281632 157344 281684 157350
rect 281632 157286 281684 157292
rect 280436 157072 280488 157078
rect 280436 157014 280488 157020
rect 280620 154556 280672 154562
rect 280620 154498 280672 154504
rect 280252 154488 280304 154494
rect 280632 154442 280660 154498
rect 280304 154436 280660 154442
rect 280252 154430 280660 154436
rect 280264 154414 280660 154430
rect 280710 153776 280766 153785
rect 280710 153711 280766 153720
rect 280724 149954 280752 153711
rect 281644 150226 281672 157286
rect 281644 150198 281718 150226
rect 273548 149926 273976 149954
rect 274284 149926 274620 149954
rect 274836 149926 275264 149954
rect 275572 149926 275908 149954
rect 276124 149926 276552 149954
rect 276768 149926 277196 149954
rect 277504 149926 277840 149954
rect 278148 149926 278484 149954
rect 278976 149926 279128 149954
rect 279436 149926 279772 149954
rect 280172 149926 280416 149954
rect 280724 149926 281060 149954
rect 281690 149940 281718 150198
rect 282012 149954 282040 159258
rect 283196 159180 283248 159186
rect 283196 159122 283248 159128
rect 283104 156664 283156 156670
rect 283104 156606 283156 156612
rect 282920 152244 282972 152250
rect 282920 152186 282972 152192
rect 282932 150226 282960 152186
rect 283116 150550 283144 156606
rect 283208 151842 283236 159122
rect 283288 154624 283340 154630
rect 283288 154566 283340 154572
rect 283196 151836 283248 151842
rect 283196 151778 283248 151784
rect 283104 150544 283156 150550
rect 283104 150486 283156 150492
rect 282932 150198 283006 150226
rect 282012 149926 282348 149954
rect 282978 149940 283006 150198
rect 283300 149954 283328 154566
rect 283392 154494 283420 163254
rect 283838 163200 283894 164400
rect 284666 163200 284722 164400
rect 285494 163200 285550 164400
rect 285692 163254 286272 163282
rect 283852 157282 283880 163200
rect 284680 159186 284708 163200
rect 285128 159248 285180 159254
rect 285128 159190 285180 159196
rect 284668 159180 284720 159186
rect 284668 159122 284720 159128
rect 283840 157276 283892 157282
rect 283840 157218 283892 157224
rect 283380 154488 283432 154494
rect 283380 154430 283432 154436
rect 284576 152992 284628 152998
rect 284576 152934 284628 152940
rect 283932 150544 283984 150550
rect 283932 150486 283984 150492
rect 283944 149954 283972 150486
rect 284588 149954 284616 152934
rect 285140 149954 285168 159190
rect 285508 153202 285536 163200
rect 285692 154562 285720 163254
rect 286244 163146 286272 163254
rect 286322 163200 286378 164400
rect 287150 163200 287206 164400
rect 287978 163200 288034 164400
rect 288898 163200 288954 164400
rect 289726 163200 289782 164400
rect 290554 163200 290610 164400
rect 291382 163200 291438 164400
rect 292210 163200 292266 164400
rect 293038 163200 293094 164400
rect 293866 163200 293922 164400
rect 294786 163200 294842 164400
rect 295614 163200 295670 164400
rect 296442 163200 296498 164400
rect 297270 163200 297326 164400
rect 298098 163200 298154 164400
rect 298664 163254 298876 163282
rect 286336 163146 286364 163200
rect 286244 163118 286364 163146
rect 285772 159180 285824 159186
rect 285772 159122 285824 159128
rect 285588 154556 285640 154562
rect 285588 154498 285640 154504
rect 285680 154556 285732 154562
rect 285680 154498 285732 154504
rect 285600 154442 285628 154498
rect 285600 154414 285720 154442
rect 285496 153196 285548 153202
rect 285496 153138 285548 153144
rect 285692 151814 285720 154414
rect 285784 152250 285812 159122
rect 287164 157146 287192 163200
rect 287992 159254 288020 163200
rect 287980 159248 288032 159254
rect 287980 159190 288032 159196
rect 288912 159186 288940 163200
rect 288164 159180 288216 159186
rect 288164 159122 288216 159128
rect 288900 159180 288952 159186
rect 288900 159122 288952 159128
rect 287152 157140 287204 157146
rect 287152 157082 287204 157088
rect 286232 156324 286284 156330
rect 286232 156266 286284 156272
rect 285772 152244 285824 152250
rect 285772 152186 285824 152192
rect 286244 151814 286272 156266
rect 288176 152998 288204 159122
rect 288992 156732 289044 156738
rect 288992 156674 289044 156680
rect 288440 154012 288492 154018
rect 288440 153954 288492 153960
rect 288164 152992 288216 152998
rect 288164 152934 288216 152940
rect 287796 152380 287848 152386
rect 287796 152322 287848 152328
rect 287152 151836 287204 151842
rect 285692 151786 285812 151814
rect 286244 151786 286456 151814
rect 285784 149954 285812 151786
rect 286428 149954 286456 151786
rect 287152 151778 287204 151784
rect 287164 149954 287192 151778
rect 287808 149954 287836 152322
rect 288452 149954 288480 153954
rect 289004 149954 289032 156674
rect 289740 155786 289768 163200
rect 290280 159384 290332 159390
rect 290280 159326 290332 159332
rect 289728 155780 289780 155786
rect 289728 155722 289780 155728
rect 289912 152992 289964 152998
rect 289912 152934 289964 152940
rect 289924 149954 289952 152934
rect 290292 149954 290320 159326
rect 290568 157214 290596 163200
rect 290556 157208 290608 157214
rect 290556 157150 290608 157156
rect 291292 153944 291344 153950
rect 291292 153886 291344 153892
rect 291304 150226 291332 153886
rect 291396 152998 291424 163200
rect 291568 156868 291620 156874
rect 291568 156810 291620 156816
rect 291384 152992 291436 152998
rect 291384 152934 291436 152940
rect 291304 150198 291378 150226
rect 283300 149926 283636 149954
rect 283944 149926 284280 149954
rect 284588 149926 284924 149954
rect 285140 149926 285568 149954
rect 285784 149926 286212 149954
rect 286428 149926 286856 149954
rect 287164 149926 287500 149954
rect 287808 149926 288144 149954
rect 288452 149926 288788 149954
rect 289004 149926 289432 149954
rect 289924 149926 290076 149954
rect 290292 149926 290720 149954
rect 291350 149940 291378 150198
rect 291580 149954 291608 156810
rect 292224 152386 292252 163200
rect 293052 155854 293080 163200
rect 293880 156738 293908 163200
rect 294800 159390 294828 163200
rect 295628 159526 295656 163200
rect 295432 159520 295484 159526
rect 295432 159462 295484 159468
rect 295616 159520 295668 159526
rect 295616 159462 295668 159468
rect 294788 159384 294840 159390
rect 294788 159326 294840 159332
rect 294788 159044 294840 159050
rect 294788 158986 294840 158992
rect 294052 156800 294104 156806
rect 294052 156742 294104 156748
rect 293868 156732 293920 156738
rect 293868 156674 293920 156680
rect 293040 155848 293092 155854
rect 293040 155790 293092 155796
rect 293592 153672 293644 153678
rect 293592 153614 293644 153620
rect 292948 152516 293000 152522
rect 292948 152458 293000 152464
rect 292578 152416 292634 152425
rect 292212 152380 292264 152386
rect 292578 152351 292634 152360
rect 292212 152322 292264 152328
rect 292592 150226 292620 152351
rect 292592 150198 292666 150226
rect 291580 149926 292008 149954
rect 292638 149940 292666 150198
rect 292960 149954 292988 152458
rect 293604 149954 293632 153614
rect 294064 151814 294092 156742
rect 294064 151786 294184 151814
rect 294156 149954 294184 151786
rect 294800 149954 294828 158986
rect 295444 149954 295472 159462
rect 296456 155922 296484 163200
rect 297284 156806 297312 163200
rect 298008 159452 298060 159458
rect 298008 159394 298060 159400
rect 297272 156800 297324 156806
rect 297272 156742 297324 156748
rect 296444 155916 296496 155922
rect 296444 155858 296496 155864
rect 296812 155304 296864 155310
rect 296812 155246 296864 155252
rect 296168 153808 296220 153814
rect 296168 153750 296220 153756
rect 296180 149954 296208 153750
rect 296824 149954 296852 155246
rect 297456 152584 297508 152590
rect 297456 152526 297508 152532
rect 297468 149954 297496 152526
rect 298020 151814 298048 159394
rect 298112 159050 298140 163200
rect 298100 159044 298152 159050
rect 298100 158986 298152 158992
rect 298664 152522 298692 163254
rect 298848 163146 298876 163254
rect 298926 163200 298982 164400
rect 299754 163200 299810 164400
rect 300674 163200 300730 164400
rect 301502 163200 301558 164400
rect 302330 163200 302386 164400
rect 303158 163200 303214 164400
rect 303632 163254 303936 163282
rect 298940 163146 298968 163200
rect 298848 163118 298968 163146
rect 299664 159044 299716 159050
rect 299664 158986 299716 158992
rect 299480 158976 299532 158982
rect 299480 158918 299532 158924
rect 298744 153740 298796 153746
rect 298744 153682 298796 153688
rect 298652 152516 298704 152522
rect 298652 152458 298704 152464
rect 298020 151786 298140 151814
rect 298112 149954 298140 151786
rect 298756 149954 298784 153682
rect 299492 150550 299520 158918
rect 299572 158024 299624 158030
rect 299572 157966 299624 157972
rect 299480 150544 299532 150550
rect 299480 150486 299532 150492
rect 299584 149954 299612 157966
rect 299676 151842 299704 158986
rect 299768 155310 299796 163200
rect 300688 156874 300716 163200
rect 301516 159458 301544 163200
rect 301504 159452 301556 159458
rect 301504 159394 301556 159400
rect 302344 159118 302372 163200
rect 302332 159112 302384 159118
rect 302332 159054 302384 159060
rect 300676 156868 300728 156874
rect 300676 156810 300728 156816
rect 299756 155304 299808 155310
rect 299756 155246 299808 155252
rect 302516 155236 302568 155242
rect 302516 155178 302568 155184
rect 301320 153604 301372 153610
rect 301320 153546 301372 153552
rect 300860 151972 300912 151978
rect 300860 151914 300912 151920
rect 299664 151836 299716 151842
rect 299664 151778 299716 151784
rect 300032 150544 300084 150550
rect 300032 150486 300084 150492
rect 300044 149954 300072 150486
rect 300872 149954 300900 151914
rect 301332 149954 301360 153546
rect 302528 149954 302556 155178
rect 303172 155106 303200 163200
rect 303252 158908 303304 158914
rect 303252 158850 303304 158856
rect 303160 155100 303212 155106
rect 303160 155042 303212 155048
rect 302608 151904 302660 151910
rect 302608 151846 302660 151852
rect 292960 149926 293296 149954
rect 293604 149926 293940 149954
rect 294156 149926 294584 149954
rect 294800 149926 295228 149954
rect 295444 149926 295872 149954
rect 296180 149926 296516 149954
rect 296824 149926 297160 149954
rect 297468 149926 297804 149954
rect 298112 149926 298448 149954
rect 298756 149926 299092 149954
rect 299584 149926 299736 149954
rect 300044 149926 300380 149954
rect 300872 149926 301024 149954
rect 301332 149926 301668 149954
rect 302312 149926 302556 149954
rect 302620 149954 302648 151846
rect 303264 149954 303292 158850
rect 303632 152590 303660 163254
rect 303908 163146 303936 163254
rect 303986 163200 304042 164400
rect 304092 163254 304764 163282
rect 304000 163146 304028 163200
rect 303908 163118 304028 163146
rect 303804 153876 303856 153882
rect 303804 153818 303856 153824
rect 303620 152584 303672 152590
rect 303620 152526 303672 152532
rect 303816 149954 303844 153818
rect 304092 151978 304120 163254
rect 304736 163146 304764 163254
rect 304814 163200 304870 164400
rect 305642 163200 305698 164400
rect 306562 163200 306618 164400
rect 307390 163200 307446 164400
rect 308218 163200 308274 164400
rect 309046 163200 309102 164400
rect 309152 163254 309824 163282
rect 304828 163146 304856 163200
rect 304736 163118 304856 163146
rect 305184 159656 305236 159662
rect 305184 159598 305236 159604
rect 304356 158092 304408 158098
rect 304356 158034 304408 158040
rect 304080 151972 304132 151978
rect 304080 151914 304132 151920
rect 304368 149954 304396 158034
rect 305196 149954 305224 159598
rect 305656 158914 305684 163200
rect 305644 158908 305696 158914
rect 305644 158850 305696 158856
rect 306576 155242 306604 163200
rect 307404 159050 307432 163200
rect 308232 159730 308260 163200
rect 308128 159724 308180 159730
rect 308128 159666 308180 159672
rect 308220 159724 308272 159730
rect 308220 159666 308272 159672
rect 307392 159044 307444 159050
rect 307392 158986 307444 158992
rect 307392 158908 307444 158914
rect 307392 158850 307444 158856
rect 306932 158160 306984 158166
rect 306932 158102 306984 158108
rect 306564 155236 306616 155242
rect 306564 155178 306616 155184
rect 306380 154148 306432 154154
rect 306380 154090 306432 154096
rect 305736 152176 305788 152182
rect 305736 152118 305788 152124
rect 305748 149954 305776 152118
rect 306392 149954 306420 154090
rect 306944 149954 306972 158102
rect 307404 151910 307432 158850
rect 307760 152652 307812 152658
rect 307760 152594 307812 152600
rect 307392 151904 307444 151910
rect 307392 151846 307444 151852
rect 307772 149954 307800 152594
rect 308140 151814 308168 159666
rect 309060 159662 309088 163200
rect 309048 159656 309100 159662
rect 309048 159598 309100 159604
rect 309152 153882 309180 163254
rect 309796 163146 309824 163254
rect 309874 163200 309930 164400
rect 310702 163200 310758 164400
rect 311530 163200 311586 164400
rect 312450 163200 312506 164400
rect 313278 163200 313334 164400
rect 314106 163200 314162 164400
rect 314934 163200 314990 164400
rect 315762 163200 315818 164400
rect 316052 163254 316540 163282
rect 309888 163146 309916 163200
rect 309796 163118 309916 163146
rect 310612 159588 310664 159594
rect 310612 159530 310664 159536
rect 309508 155372 309560 155378
rect 309508 155314 309560 155320
rect 309232 154080 309284 154086
rect 309232 154022 309284 154028
rect 309140 153876 309192 153882
rect 309140 153818 309192 153824
rect 308140 151786 308260 151814
rect 308232 149954 308260 151786
rect 309244 150226 309272 154022
rect 309244 150198 309318 150226
rect 302620 149926 302956 149954
rect 303264 149926 303600 149954
rect 303816 149926 304152 149954
rect 304368 149926 304796 149954
rect 305196 149926 305440 149954
rect 305748 149926 306084 149954
rect 306392 149926 306728 149954
rect 306944 149926 307372 149954
rect 307772 149926 308016 149954
rect 308232 149926 308660 149954
rect 309290 149940 309318 150198
rect 309520 149954 309548 155314
rect 310624 150226 310652 159530
rect 310716 158914 310744 163200
rect 311544 161474 311572 163200
rect 311544 161446 311664 161474
rect 310704 158908 310756 158914
rect 310704 158850 310756 158856
rect 311532 153536 311584 153542
rect 311532 153478 311584 153484
rect 310888 152720 310940 152726
rect 310888 152662 310940 152668
rect 310578 150198 310652 150226
rect 309520 149926 309948 149954
rect 310578 149940 310606 150198
rect 310900 149954 310928 152662
rect 311544 149954 311572 153478
rect 311636 152658 311664 161446
rect 312464 159866 312492 163200
rect 312360 159860 312412 159866
rect 312360 159802 312412 159808
rect 312452 159860 312504 159866
rect 312452 159802 312504 159808
rect 312372 158914 312400 159802
rect 311992 158908 312044 158914
rect 311992 158850 312044 158856
rect 312360 158908 312412 158914
rect 312360 158850 312412 158856
rect 312004 152726 312032 158850
rect 312084 155440 312136 155446
rect 312084 155382 312136 155388
rect 311992 152720 312044 152726
rect 311992 152662 312044 152668
rect 311624 152652 311676 152658
rect 311624 152594 311676 152600
rect 312096 149954 312124 155382
rect 313292 153950 313320 163200
rect 313372 159860 313424 159866
rect 313372 159802 313424 159808
rect 313280 153944 313332 153950
rect 313280 153886 313332 153892
rect 312820 152856 312872 152862
rect 312820 152798 312872 152804
rect 312832 149954 312860 152798
rect 313384 152425 313412 159802
rect 314120 159798 314148 163200
rect 313464 159792 313516 159798
rect 313464 159734 313516 159740
rect 314108 159792 314160 159798
rect 314108 159734 314160 159740
rect 313370 152416 313426 152425
rect 313370 152351 313426 152360
rect 313476 149954 313504 159734
rect 314948 158982 314976 163200
rect 315776 159594 315804 163200
rect 315764 159588 315816 159594
rect 315764 159530 315816 159536
rect 314936 158976 314988 158982
rect 314936 158918 314988 158924
rect 314752 158228 314804 158234
rect 314752 158170 314804 158176
rect 314108 154216 314160 154222
rect 314108 154158 314160 154164
rect 314120 149954 314148 154158
rect 314764 149954 314792 158170
rect 316052 154018 316080 163254
rect 316512 163146 316540 163254
rect 316590 163200 316646 164400
rect 317418 163200 317474 164400
rect 317524 163254 318288 163282
rect 316604 163146 316632 163200
rect 316512 163118 316632 163146
rect 316316 158840 316368 158846
rect 316316 158782 316368 158788
rect 316040 154012 316092 154018
rect 316040 153954 316092 153960
rect 316328 152862 316356 158782
rect 316776 153400 316828 153406
rect 316776 153342 316828 153348
rect 316316 152856 316368 152862
rect 316316 152798 316368 152804
rect 315396 152788 315448 152794
rect 315396 152730 315448 152736
rect 315408 149954 315436 152730
rect 316040 152448 316092 152454
rect 316040 152390 316092 152396
rect 316052 149954 316080 152390
rect 316788 149954 316816 153342
rect 317432 152794 317460 163200
rect 317420 152788 317472 152794
rect 317420 152730 317472 152736
rect 317524 152454 317552 163254
rect 318260 163146 318288 163254
rect 318338 163200 318394 164400
rect 319166 163200 319222 164400
rect 319994 163200 320050 164400
rect 320822 163200 320878 164400
rect 321650 163200 321706 164400
rect 322478 163200 322534 164400
rect 323306 163200 323362 164400
rect 324226 163200 324282 164400
rect 324332 163254 325004 163282
rect 318352 163146 318380 163200
rect 318260 163118 318380 163146
rect 318800 158908 318852 158914
rect 318800 158850 318852 158856
rect 317604 155508 317656 155514
rect 317604 155450 317656 155456
rect 317512 152448 317564 152454
rect 317512 152390 317564 152396
rect 317616 150226 317644 155450
rect 317972 152856 318024 152862
rect 317972 152798 318024 152804
rect 317616 150198 317690 150226
rect 310900 149926 311236 149954
rect 311544 149926 311880 149954
rect 312096 149926 312524 149954
rect 312832 149926 313168 149954
rect 313476 149926 313812 149954
rect 314120 149926 314456 149954
rect 314764 149926 315100 149954
rect 315408 149926 315744 149954
rect 316052 149926 316388 149954
rect 316788 149926 317032 149954
rect 317662 149940 317690 150198
rect 317984 149954 318012 152798
rect 318812 149954 318840 158850
rect 319180 158846 319208 163200
rect 319168 158840 319220 158846
rect 319168 158782 319220 158788
rect 320008 155378 320036 163200
rect 320836 158914 320864 163200
rect 320824 158908 320876 158914
rect 320824 158850 320876 158856
rect 321664 158846 321692 163200
rect 322492 159866 322520 163200
rect 322480 159860 322532 159866
rect 322480 159802 322532 159808
rect 321652 158840 321704 158846
rect 321652 158782 321704 158788
rect 320272 158772 320324 158778
rect 320272 158714 320324 158720
rect 320180 155576 320232 155582
rect 320180 155518 320232 155524
rect 319996 155372 320048 155378
rect 319996 155314 320048 155320
rect 319260 154284 319312 154290
rect 319260 154226 319312 154232
rect 319272 149954 319300 154226
rect 320192 150226 320220 155518
rect 320284 152794 320312 158714
rect 321560 158704 321612 158710
rect 321560 158646 321612 158652
rect 321192 153128 321244 153134
rect 321192 153070 321244 153076
rect 320272 152788 320324 152794
rect 320272 152730 320324 152736
rect 320732 152652 320784 152658
rect 320732 152594 320784 152600
rect 320824 152652 320876 152658
rect 320824 152594 320876 152600
rect 320548 152312 320600 152318
rect 320548 152254 320600 152260
rect 320192 150198 320266 150226
rect 317984 149926 318320 149954
rect 318812 149926 318964 149954
rect 319272 149926 319608 149954
rect 320238 149940 320266 150198
rect 320560 149954 320588 152254
rect 320744 152182 320772 152594
rect 320836 152454 320864 152594
rect 320824 152448 320876 152454
rect 320824 152390 320876 152396
rect 320824 152312 320876 152318
rect 320824 152254 320876 152260
rect 320732 152176 320784 152182
rect 320732 152118 320784 152124
rect 320836 152046 320864 152254
rect 320824 152040 320876 152046
rect 320824 151982 320876 151988
rect 321204 149954 321232 153070
rect 321572 152046 321600 158646
rect 322112 155644 322164 155650
rect 322112 155586 322164 155592
rect 321836 153468 321888 153474
rect 321836 153410 321888 153416
rect 321560 152040 321612 152046
rect 321560 151982 321612 151988
rect 321848 149954 321876 153410
rect 322124 151814 322152 155586
rect 323320 154086 323348 163200
rect 323676 159928 323728 159934
rect 323676 159870 323728 159876
rect 323308 154080 323360 154086
rect 323308 154022 323360 154028
rect 323124 152788 323176 152794
rect 323124 152730 323176 152736
rect 322124 151786 322428 151814
rect 322400 149954 322428 151786
rect 323136 149954 323164 152730
rect 323688 149954 323716 159870
rect 324240 152794 324268 163200
rect 324332 153134 324360 163254
rect 324976 163146 325004 163254
rect 325054 163200 325110 164400
rect 325882 163200 325938 164400
rect 326710 163200 326766 164400
rect 327538 163200 327594 164400
rect 328366 163200 328422 164400
rect 329194 163200 329250 164400
rect 330114 163200 330170 164400
rect 330942 163200 330998 164400
rect 331232 163254 331720 163282
rect 325068 163146 325096 163200
rect 324976 163118 325096 163146
rect 324964 155712 325016 155718
rect 324964 155654 325016 155660
rect 324412 153264 324464 153270
rect 324412 153206 324464 153212
rect 324320 153128 324372 153134
rect 324320 153070 324372 153076
rect 324228 152788 324280 152794
rect 324228 152730 324280 152736
rect 324424 149954 324452 153206
rect 324976 149954 325004 155654
rect 325896 152454 325924 163200
rect 326724 154154 326752 163200
rect 327552 158778 327580 163200
rect 328380 159934 328408 163200
rect 329208 160002 329236 163200
rect 328460 159996 328512 160002
rect 328460 159938 328512 159944
rect 329196 159996 329248 160002
rect 329196 159938 329248 159944
rect 328368 159928 328420 159934
rect 328368 159870 328420 159876
rect 327540 158772 327592 158778
rect 327540 158714 327592 158720
rect 327540 157004 327592 157010
rect 327540 156946 327592 156952
rect 326712 154148 326764 154154
rect 326712 154090 326764 154096
rect 327080 153332 327132 153338
rect 327080 153274 327132 153280
rect 326344 153060 326396 153066
rect 326344 153002 326396 153008
rect 325884 152448 325936 152454
rect 325884 152390 325936 152396
rect 325700 152312 325752 152318
rect 325700 152254 325752 152260
rect 325712 149954 325740 152254
rect 326356 149954 326384 153002
rect 327092 149954 327120 153274
rect 327552 149954 327580 156946
rect 328472 150550 328500 159938
rect 328550 159488 328606 159497
rect 328550 159423 328606 159432
rect 328460 150544 328512 150550
rect 328460 150486 328512 150492
rect 328564 150226 328592 159423
rect 330024 156936 330076 156942
rect 330024 156878 330076 156884
rect 329932 154420 329984 154426
rect 329932 154362 329984 154368
rect 328920 150544 328972 150550
rect 328920 150486 328972 150492
rect 328564 150198 328638 150226
rect 320560 149926 320896 149954
rect 321204 149926 321540 149954
rect 321848 149926 322184 149954
rect 322400 149926 322828 149954
rect 323136 149926 323472 149954
rect 323688 149926 324116 149954
rect 324424 149926 324760 149954
rect 324976 149926 325404 149954
rect 325712 149926 326048 149954
rect 326356 149926 326692 149954
rect 327092 149926 327336 149954
rect 327552 149926 327980 149954
rect 328610 149940 328638 150198
rect 328932 149954 328960 150486
rect 329944 150226 329972 154362
rect 330036 151814 330064 156878
rect 330128 155446 330156 163200
rect 330116 155440 330168 155446
rect 330116 155382 330168 155388
rect 330956 153066 330984 163200
rect 330944 153060 330996 153066
rect 330944 153002 330996 153008
rect 331232 152318 331260 163254
rect 331692 163146 331720 163254
rect 331770 163200 331826 164400
rect 332598 163200 332654 164400
rect 333426 163200 333482 164400
rect 334254 163200 334310 164400
rect 335082 163200 335138 164400
rect 335372 163254 335952 163282
rect 331784 163146 331812 163200
rect 331692 163118 331812 163146
rect 332140 154352 332192 154358
rect 332140 154294 332192 154300
rect 331496 152924 331548 152930
rect 331496 152866 331548 152872
rect 331220 152312 331272 152318
rect 331220 152254 331272 152260
rect 330852 152108 330904 152114
rect 330852 152050 330904 152056
rect 330036 151786 330156 151814
rect 329898 150198 329972 150226
rect 328932 149926 329268 149954
rect 329898 149940 329926 150198
rect 330128 149954 330156 151786
rect 330864 149954 330892 152050
rect 331508 149954 331536 152866
rect 332152 149954 332180 154294
rect 332612 152930 332640 163200
rect 332692 160064 332744 160070
rect 332692 160006 332744 160012
rect 332600 152924 332652 152930
rect 332600 152866 332652 152872
rect 332704 150550 332732 160006
rect 332876 157072 332928 157078
rect 332876 157014 332928 157020
rect 332692 150544 332744 150550
rect 332692 150486 332744 150492
rect 332888 149954 332916 157014
rect 333440 155514 333468 163200
rect 334268 159322 334296 163200
rect 335096 160070 335124 163200
rect 335084 160064 335136 160070
rect 335084 160006 335136 160012
rect 333980 159316 334032 159322
rect 333980 159258 334032 159264
rect 334256 159316 334308 159322
rect 334256 159258 334308 159264
rect 333428 155508 333480 155514
rect 333428 155450 333480 155456
rect 333428 150544 333480 150550
rect 333428 150486 333480 150492
rect 333440 149954 333468 150486
rect 333992 149954 334020 159258
rect 334624 154488 334676 154494
rect 334624 154430 334676 154436
rect 334636 149954 334664 154430
rect 335372 152114 335400 163254
rect 335924 163146 335952 163254
rect 336002 163200 336058 164400
rect 336830 163200 336886 164400
rect 337658 163200 337714 164400
rect 338486 163200 338542 164400
rect 339314 163200 339370 164400
rect 339512 163254 340092 163282
rect 336016 163146 336044 163200
rect 335924 163118 336044 163146
rect 335820 159520 335872 159526
rect 336188 159520 336240 159526
rect 335872 159480 336136 159508
rect 335820 159462 335872 159468
rect 336108 159390 336136 159480
rect 336188 159462 336240 159468
rect 336004 159384 336056 159390
rect 336004 159326 336056 159332
rect 336096 159384 336148 159390
rect 336096 159326 336148 159332
rect 336016 159236 336044 159326
rect 336200 159236 336228 159462
rect 336016 159208 336228 159236
rect 335452 157276 335504 157282
rect 335452 157218 335504 157224
rect 335360 152108 335412 152114
rect 335360 152050 335412 152056
rect 335464 149954 335492 157218
rect 336844 154222 336872 163200
rect 337672 155582 337700 163200
rect 338500 160070 338528 163200
rect 338488 160064 338540 160070
rect 338488 160006 338540 160012
rect 339328 159254 339356 163200
rect 338396 159248 338448 159254
rect 338396 159190 338448 159196
rect 339316 159248 339368 159254
rect 339316 159190 339368 159196
rect 338120 157140 338172 157146
rect 338120 157082 338172 157088
rect 337660 155576 337712 155582
rect 337660 155518 337712 155524
rect 337200 154556 337252 154562
rect 337200 154498 337252 154504
rect 336832 154216 336884 154222
rect 336832 154158 336884 154164
rect 336740 153196 336792 153202
rect 336740 153138 336792 153144
rect 335912 152244 335964 152250
rect 335912 152186 335964 152192
rect 335924 149954 335952 152186
rect 336752 149954 336780 153138
rect 337212 149954 337240 154498
rect 338132 150226 338160 157082
rect 338132 150198 338206 150226
rect 330128 149926 330556 149954
rect 330864 149926 331200 149954
rect 331508 149926 331844 149954
rect 332152 149926 332488 149954
rect 332888 149926 333132 149954
rect 333440 149926 333776 149954
rect 333992 149926 334420 149954
rect 334636 149926 334972 149954
rect 335464 149926 335616 149954
rect 335924 149926 336260 149954
rect 336752 149926 336904 149954
rect 337212 149926 337548 149954
rect 338178 149940 338206 150198
rect 338408 149954 338436 159190
rect 339040 159180 339092 159186
rect 339040 159122 339092 159128
rect 339052 149954 339080 159122
rect 339512 154358 339540 163254
rect 340064 163146 340092 163254
rect 340142 163200 340198 164400
rect 340970 163200 341026 164400
rect 341890 163200 341946 164400
rect 341996 163254 342208 163282
rect 340156 163146 340184 163200
rect 340064 163118 340184 163146
rect 339684 160064 339736 160070
rect 339684 160006 339736 160012
rect 339592 155780 339644 155786
rect 339592 155722 339644 155728
rect 339500 154352 339552 154358
rect 339500 154294 339552 154300
rect 339604 151814 339632 155722
rect 339696 153202 339724 160006
rect 340052 157208 340104 157214
rect 340052 157150 340104 157156
rect 339684 153196 339736 153202
rect 339684 153138 339736 153144
rect 340064 151814 340092 157150
rect 340984 155718 341012 163200
rect 341904 163146 341932 163200
rect 341996 163146 342024 163254
rect 341904 163118 342024 163146
rect 342180 159474 342208 163254
rect 342718 163200 342774 164400
rect 343546 163200 343602 164400
rect 344374 163200 344430 164400
rect 345202 163200 345258 164400
rect 346030 163200 346086 164400
rect 346412 163254 346808 163282
rect 342732 159730 342760 163200
rect 342720 159724 342772 159730
rect 342720 159666 342772 159672
rect 342272 159594 342484 159610
rect 342260 159588 342496 159594
rect 342312 159582 342444 159588
rect 342260 159530 342312 159536
rect 342444 159530 342496 159536
rect 341432 159452 341484 159458
rect 342180 159446 342392 159474
rect 341432 159394 341484 159400
rect 341444 159186 341472 159394
rect 342364 159390 342392 159446
rect 343456 159452 343508 159458
rect 343456 159394 343508 159400
rect 342260 159384 342312 159390
rect 342260 159326 342312 159332
rect 342352 159384 342404 159390
rect 342352 159326 342404 159332
rect 341432 159180 341484 159186
rect 341432 159122 341484 159128
rect 340972 155712 341024 155718
rect 340972 155654 341024 155660
rect 342272 152998 342300 159326
rect 342812 156732 342864 156738
rect 342812 156674 342864 156680
rect 342352 155848 342404 155854
rect 342352 155790 342404 155796
rect 341064 152992 341116 152998
rect 341064 152934 341116 152940
rect 342260 152992 342312 152998
rect 342260 152934 342312 152940
rect 339604 151786 339724 151814
rect 340064 151786 340368 151814
rect 339696 149954 339724 151786
rect 340340 149954 340368 151786
rect 341076 149954 341104 152934
rect 341708 152380 341760 152386
rect 341708 152322 341760 152328
rect 341720 149954 341748 152322
rect 342364 149954 342392 155790
rect 342824 151814 342852 156674
rect 343468 151814 343496 159394
rect 343560 154290 343588 163200
rect 343824 159724 343876 159730
rect 343824 159666 343876 159672
rect 343548 154284 343600 154290
rect 343548 154226 343600 154232
rect 343836 152386 343864 159666
rect 344388 155650 344416 163200
rect 345216 157334 345244 163200
rect 346044 159390 346072 163200
rect 346032 159384 346084 159390
rect 346032 159326 346084 159332
rect 345216 157306 345336 157334
rect 345204 155916 345256 155922
rect 345204 155858 345256 155864
rect 344376 155644 344428 155650
rect 344376 155586 344428 155592
rect 344284 152992 344336 152998
rect 344284 152934 344336 152940
rect 343824 152380 343876 152386
rect 343824 152322 343876 152328
rect 342824 151786 342944 151814
rect 343468 151786 343680 151814
rect 342916 149954 342944 151786
rect 343652 149954 343680 151786
rect 344296 149954 344324 152934
rect 345216 150226 345244 155858
rect 345308 152998 345336 157306
rect 345572 156800 345624 156806
rect 345572 156742 345624 156748
rect 345296 152992 345348 152998
rect 345296 152934 345348 152940
rect 345216 150198 345290 150226
rect 338408 149926 338836 149954
rect 339052 149926 339480 149954
rect 339696 149926 340124 149954
rect 340340 149926 340768 149954
rect 341076 149926 341412 149954
rect 341720 149926 342056 149954
rect 342364 149926 342700 149954
rect 342916 149926 343344 149954
rect 343652 149926 343988 149954
rect 344296 149926 344632 149954
rect 345262 149940 345290 150198
rect 345584 149954 345612 156742
rect 346412 154426 346440 163254
rect 346780 163146 346808 163254
rect 346858 163200 346914 164400
rect 347778 163200 347834 164400
rect 348160 163254 348556 163282
rect 346872 163146 346900 163200
rect 346780 163118 346900 163146
rect 347792 159730 347820 163200
rect 347780 159724 347832 159730
rect 347780 159666 347832 159672
rect 348056 156868 348108 156874
rect 348056 156810 348108 156816
rect 347964 155304 348016 155310
rect 347964 155246 348016 155252
rect 346400 154420 346452 154426
rect 346400 154362 346452 154368
rect 346860 152516 346912 152522
rect 346860 152458 346912 152464
rect 346400 151836 346452 151842
rect 346452 151786 346532 151814
rect 346400 151778 346452 151784
rect 346504 150226 346532 151786
rect 346504 150198 346578 150226
rect 345584 149926 345920 149954
rect 346550 149940 346578 150198
rect 346872 149954 346900 152458
rect 347976 149954 348004 155246
rect 346872 149926 347208 149954
rect 347852 149926 348004 149954
rect 348068 149954 348096 156810
rect 348160 152522 348188 163254
rect 348528 163146 348556 163254
rect 348606 163200 348662 164400
rect 349172 163254 349384 163282
rect 348620 163146 348648 163200
rect 348528 163118 348648 163146
rect 348792 159452 348844 159458
rect 348792 159394 348844 159400
rect 348804 159186 348832 159394
rect 348700 159180 348752 159186
rect 348700 159122 348752 159128
rect 348792 159180 348844 159186
rect 348792 159122 348844 159128
rect 348148 152516 348200 152522
rect 348148 152458 348200 152464
rect 348712 149954 348740 159122
rect 349172 152250 349200 163254
rect 349356 163146 349384 163254
rect 349434 163200 349490 164400
rect 349540 163254 350212 163282
rect 349448 163146 349476 163200
rect 349356 163118 349476 163146
rect 349252 159112 349304 159118
rect 349252 159054 349304 159060
rect 349160 152244 349212 152250
rect 349160 152186 349212 152192
rect 349264 151814 349292 159054
rect 349540 154494 349568 163254
rect 350184 163146 350212 163254
rect 350262 163200 350318 164400
rect 351090 163200 351146 164400
rect 351918 163200 351974 164400
rect 352024 163254 352696 163282
rect 350276 163146 350304 163200
rect 350184 163118 350304 163146
rect 351104 159050 351132 163200
rect 351932 159118 351960 163200
rect 351828 159112 351880 159118
rect 351828 159054 351880 159060
rect 351920 159112 351972 159118
rect 351920 159054 351972 159060
rect 351092 159044 351144 159050
rect 351092 158986 351144 158992
rect 351840 158930 351868 159054
rect 351840 158902 351960 158930
rect 349988 155100 350040 155106
rect 349988 155042 350040 155048
rect 349528 154488 349580 154494
rect 349528 154430 349580 154436
rect 349804 152380 349856 152386
rect 349804 152322 349856 152328
rect 349896 152380 349948 152386
rect 349896 152322 349948 152328
rect 349816 151842 349844 152322
rect 349908 152250 349936 152322
rect 349896 152244 349948 152250
rect 349896 152186 349948 152192
rect 349804 151836 349856 151842
rect 349264 151786 349384 151814
rect 349356 149954 349384 151786
rect 349804 151778 349856 151784
rect 350000 149954 350028 155042
rect 351932 152590 351960 158902
rect 350724 152584 350776 152590
rect 350724 152526 350776 152532
rect 351920 152584 351972 152590
rect 351920 152526 351972 152532
rect 350736 149954 350764 152526
rect 352024 152250 352052 163254
rect 352668 163146 352696 163254
rect 352746 163200 352802 164400
rect 353666 163200 353722 164400
rect 354494 163200 354550 164400
rect 354692 163254 355272 163282
rect 352760 163146 352788 163200
rect 352668 163118 352788 163146
rect 353392 159656 353444 159662
rect 353392 159598 353444 159604
rect 352472 155236 352524 155242
rect 352472 155178 352524 155184
rect 352012 152244 352064 152250
rect 352012 152186 352064 152192
rect 351368 151972 351420 151978
rect 351368 151914 351420 151920
rect 351380 149954 351408 151914
rect 352012 151904 352064 151910
rect 352012 151846 352064 151852
rect 352024 149954 352052 151846
rect 352484 151814 352512 155178
rect 353300 152584 353352 152590
rect 353300 152526 353352 152532
rect 352484 151786 352604 151814
rect 352576 149954 352604 151786
rect 353312 149954 353340 152526
rect 353404 151814 353432 159598
rect 353680 154562 353708 163200
rect 353668 154556 353720 154562
rect 353668 154498 353720 154504
rect 354508 152590 354536 163200
rect 354496 152584 354548 152590
rect 354496 152526 354548 152532
rect 354692 151978 354720 163254
rect 355244 163146 355272 163254
rect 355322 163200 355378 164400
rect 356150 163200 356206 164400
rect 356256 163254 356928 163282
rect 355336 163146 355364 163200
rect 355244 163118 355364 163146
rect 354772 159520 354824 159526
rect 354772 159462 354824 159468
rect 354680 151972 354732 151978
rect 354680 151914 354732 151920
rect 353404 151786 353892 151814
rect 353864 149954 353892 151786
rect 354784 149954 354812 159462
rect 356164 159458 356192 163200
rect 356152 159452 356204 159458
rect 356152 159394 356204 159400
rect 356256 153882 356284 163254
rect 356900 163146 356928 163254
rect 356978 163200 357034 164400
rect 357806 163200 357862 164400
rect 358634 163200 358690 164400
rect 358832 163254 359504 163282
rect 356992 163146 357020 163200
rect 356900 163118 357020 163146
rect 357440 159656 357492 159662
rect 357440 159598 357492 159604
rect 357452 158846 357480 159598
rect 357820 158982 357848 163200
rect 357992 159792 358044 159798
rect 357992 159734 358044 159740
rect 357532 158976 357584 158982
rect 357532 158918 357584 158924
rect 357808 158976 357860 158982
rect 357808 158918 357860 158924
rect 357440 158840 357492 158846
rect 357440 158782 357492 158788
rect 355232 153876 355284 153882
rect 355232 153818 355284 153824
rect 356244 153876 356296 153882
rect 356244 153818 356296 153824
rect 355244 149954 355272 153818
rect 356060 152720 356112 152726
rect 356060 152662 356112 152668
rect 356072 149954 356100 152662
rect 357438 152416 357494 152425
rect 357438 152351 357494 152360
rect 356520 152176 356572 152182
rect 356520 152118 356572 152124
rect 356532 149954 356560 152118
rect 357452 150226 357480 152351
rect 357544 152182 357572 158918
rect 357808 153944 357860 153950
rect 357808 153886 357860 153892
rect 357532 152176 357584 152182
rect 357532 152118 357584 152124
rect 357452 150198 357526 150226
rect 348068 149926 348496 149954
rect 348712 149926 349140 149954
rect 349356 149926 349784 149954
rect 350000 149926 350428 149954
rect 350736 149926 351072 149954
rect 351380 149926 351716 149954
rect 352024 149926 352360 149954
rect 352576 149926 353004 149954
rect 353312 149926 353648 149954
rect 353864 149926 354292 149954
rect 354784 149926 354936 149954
rect 355244 149926 355580 149954
rect 356072 149926 356224 149954
rect 356532 149926 356868 149954
rect 357498 149940 357526 150198
rect 357820 149954 357848 153886
rect 358004 151814 358032 159734
rect 358648 159526 358676 163200
rect 358636 159520 358688 159526
rect 358636 159462 358688 159468
rect 358832 152726 358860 163254
rect 359476 163146 359504 163254
rect 359554 163200 359610 164400
rect 360382 163200 360438 164400
rect 361210 163200 361266 164400
rect 361592 163254 361988 163282
rect 359568 163146 359596 163200
rect 359476 163118 359596 163146
rect 360396 161474 360424 163200
rect 360396 161446 360516 161474
rect 359648 159588 359700 159594
rect 359648 159530 359700 159536
rect 358820 152720 358872 152726
rect 358820 152662 358872 152668
rect 359096 152176 359148 152182
rect 359096 152118 359148 152124
rect 358004 151786 358400 151814
rect 358372 149954 358400 151786
rect 359108 149954 359136 152118
rect 359660 149954 359688 159530
rect 360384 154012 360436 154018
rect 360384 153954 360436 153960
rect 360396 149954 360424 153954
rect 360488 153814 360516 161446
rect 361224 158914 361252 163200
rect 361212 158908 361264 158914
rect 361212 158850 361264 158856
rect 360476 153808 360528 153814
rect 360476 153750 360528 153756
rect 361592 152862 361620 163254
rect 361960 163146 361988 163254
rect 362038 163200 362094 164400
rect 362866 163200 362922 164400
rect 363064 163254 363644 163282
rect 362052 163146 362080 163200
rect 361960 163118 362080 163146
rect 362880 159594 362908 163200
rect 362868 159588 362920 159594
rect 362868 159530 362920 159536
rect 362960 158840 363012 158846
rect 362960 158782 363012 158788
rect 361028 152856 361080 152862
rect 361028 152798 361080 152804
rect 361580 152856 361632 152862
rect 361580 152798 361632 152804
rect 361040 149954 361068 152798
rect 361672 152652 361724 152658
rect 361672 152594 361724 152600
rect 361684 149954 361712 152594
rect 362316 152040 362368 152046
rect 362316 151982 362368 151988
rect 362328 149954 362356 151982
rect 362972 150550 363000 158782
rect 363064 153950 363092 163254
rect 363616 163146 363644 163254
rect 363694 163200 363750 164400
rect 364522 163200 364578 164400
rect 365442 163200 365498 164400
rect 365732 163254 366220 163282
rect 363708 163146 363736 163200
rect 363616 163118 363736 163146
rect 363236 159656 363288 159662
rect 363236 159598 363288 159604
rect 363144 155372 363196 155378
rect 363144 155314 363196 155320
rect 363052 153944 363104 153950
rect 363052 153886 363104 153892
rect 362960 150544 363012 150550
rect 362960 150486 363012 150492
rect 363156 149954 363184 155314
rect 363248 151910 363276 159598
rect 364536 152658 364564 163200
rect 364800 159860 364852 159866
rect 364800 159802 364852 159808
rect 364524 152652 364576 152658
rect 364524 152594 364576 152600
rect 363236 151904 363288 151910
rect 363236 151846 363288 151852
rect 364340 151904 364392 151910
rect 364340 151846 364392 151852
rect 363604 150544 363656 150550
rect 363604 150486 363656 150492
rect 363616 149954 363644 150486
rect 364352 149954 364380 151846
rect 364812 149954 364840 159802
rect 365456 159798 365484 163200
rect 365444 159792 365496 159798
rect 365444 159734 365496 159740
rect 365732 152182 365760 163254
rect 366192 163146 366220 163254
rect 366270 163200 366326 164400
rect 367098 163200 367154 164400
rect 367926 163200 367982 164400
rect 368492 163254 368704 163282
rect 366284 163146 366312 163200
rect 366192 163118 366312 163146
rect 365812 154080 365864 154086
rect 365812 154022 365864 154028
rect 365720 152176 365772 152182
rect 365720 152118 365772 152124
rect 365824 150226 365852 154022
rect 367112 154018 367140 163200
rect 367940 158846 367968 163200
rect 367928 158840 367980 158846
rect 367928 158782 367980 158788
rect 368388 158772 368440 158778
rect 368388 158714 368440 158720
rect 368020 154148 368072 154154
rect 368020 154090 368072 154096
rect 367100 154012 367152 154018
rect 367100 153954 367152 153960
rect 366732 153128 366784 153134
rect 366732 153070 366784 153076
rect 366088 152788 366140 152794
rect 366088 152730 366140 152736
rect 365778 150198 365852 150226
rect 357820 149926 358156 149954
rect 358372 149926 358800 149954
rect 359108 149926 359444 149954
rect 359660 149926 360088 149954
rect 360396 149926 360732 149954
rect 361040 149926 361376 149954
rect 361684 149926 362020 149954
rect 362328 149926 362664 149954
rect 363156 149926 363308 149954
rect 363616 149926 363952 149954
rect 364352 149926 364596 149954
rect 364812 149926 365240 149954
rect 365778 149940 365806 150198
rect 366100 149954 366128 152730
rect 366744 149954 366772 153070
rect 367376 152448 367428 152454
rect 367376 152390 367428 152396
rect 367388 149954 367416 152390
rect 368032 149954 368060 154090
rect 368400 151814 368428 158714
rect 368492 152794 368520 163254
rect 368676 163146 368704 163254
rect 368754 163200 368810 164400
rect 369582 163200 369638 164400
rect 370410 163200 370466 164400
rect 371330 163200 371386 164400
rect 372158 163200 372214 164400
rect 372632 163254 372936 163282
rect 368768 163146 368796 163200
rect 368676 163118 368796 163146
rect 369216 159928 369268 159934
rect 369216 159870 369268 159876
rect 368480 152788 368532 152794
rect 368480 152730 368532 152736
rect 368400 151786 368612 151814
rect 368584 149954 368612 151786
rect 369228 149954 369256 159870
rect 369596 159662 369624 163200
rect 369860 159996 369912 160002
rect 369860 159938 369912 159944
rect 369584 159656 369636 159662
rect 369584 159598 369636 159604
rect 369872 149954 369900 159938
rect 370424 155242 370452 163200
rect 370504 155440 370556 155446
rect 370504 155382 370556 155388
rect 370412 155236 370464 155242
rect 370412 155178 370464 155184
rect 370516 149954 370544 155382
rect 371240 153060 371292 153066
rect 371240 153002 371292 153008
rect 371252 149954 371280 153002
rect 371344 152454 371372 163200
rect 372172 159934 372200 163200
rect 372160 159928 372212 159934
rect 372160 159870 372212 159876
rect 372632 153066 372660 163254
rect 372908 163146 372936 163254
rect 372986 163200 373042 164400
rect 373814 163200 373870 164400
rect 374642 163200 374698 164400
rect 375470 163200 375526 164400
rect 376298 163200 376354 164400
rect 376864 163254 377168 163282
rect 373000 163146 373028 163200
rect 372908 163118 373028 163146
rect 373080 155508 373132 155514
rect 373080 155450 373132 155456
rect 372620 153060 372672 153066
rect 372620 153002 372672 153008
rect 372620 152924 372672 152930
rect 372620 152866 372672 152872
rect 371332 152448 371384 152454
rect 371332 152390 371384 152396
rect 371884 152312 371936 152318
rect 371884 152254 371936 152260
rect 371896 149954 371924 152254
rect 372632 149954 372660 152866
rect 373092 149954 373120 155450
rect 373828 155310 373856 163200
rect 374368 160064 374420 160070
rect 374368 160006 374420 160012
rect 374000 159316 374052 159322
rect 374000 159258 374052 159264
rect 373816 155304 373868 155310
rect 373816 155246 373868 155252
rect 374012 149954 374040 159258
rect 374092 159180 374144 159186
rect 374092 159122 374144 159128
rect 374104 159066 374132 159122
rect 374104 159038 374224 159066
rect 374196 158778 374224 159038
rect 374184 158772 374236 158778
rect 374184 158714 374236 158720
rect 374380 149954 374408 160006
rect 374656 160002 374684 163200
rect 374644 159996 374696 160002
rect 374644 159938 374696 159944
rect 375484 152930 375512 163200
rect 376312 159866 376340 163200
rect 376300 159860 376352 159866
rect 376300 159802 376352 159808
rect 376300 155576 376352 155582
rect 376300 155518 376352 155524
rect 375748 154216 375800 154222
rect 375748 154158 375800 154164
rect 375472 152924 375524 152930
rect 375472 152866 375524 152872
rect 375380 152108 375432 152114
rect 375380 152050 375432 152056
rect 375392 150226 375420 152050
rect 375392 150198 375466 150226
rect 366100 149926 366436 149954
rect 366744 149926 367080 149954
rect 367388 149926 367724 149954
rect 368032 149926 368368 149954
rect 368584 149926 369012 149954
rect 369228 149926 369656 149954
rect 369872 149926 370300 149954
rect 370516 149926 370944 149954
rect 371252 149926 371588 149954
rect 371896 149926 372232 149954
rect 372632 149926 372876 149954
rect 373092 149926 373520 149954
rect 374012 149926 374164 149954
rect 374380 149926 374808 149954
rect 375438 149940 375466 150198
rect 375760 149954 375788 154158
rect 376312 149954 376340 155518
rect 376864 154154 376892 163254
rect 377140 163146 377168 163254
rect 377218 163200 377274 164400
rect 378046 163200 378102 164400
rect 378874 163200 378930 164400
rect 379702 163200 379758 164400
rect 380176 163254 380480 163282
rect 377232 163146 377260 163200
rect 377140 163118 377260 163146
rect 377588 159248 377640 159254
rect 377588 159190 377640 159196
rect 376852 154148 376904 154154
rect 376852 154090 376904 154096
rect 377036 153196 377088 153202
rect 377036 153138 377088 153144
rect 377048 149954 377076 153138
rect 377600 149954 377628 159190
rect 378060 159118 378088 163200
rect 378888 160070 378916 163200
rect 378876 160064 378928 160070
rect 378876 160006 378928 160012
rect 379716 159730 379744 163200
rect 378600 159724 378652 159730
rect 378600 159666 378652 159672
rect 379704 159724 379756 159730
rect 379704 159666 379756 159672
rect 378048 159112 378100 159118
rect 378048 159054 378100 159060
rect 378324 154352 378376 154358
rect 378324 154294 378376 154300
rect 378336 149954 378364 154294
rect 378612 152046 378640 159666
rect 379428 158772 379480 158778
rect 379428 158714 379480 158720
rect 378692 155712 378744 155718
rect 378692 155654 378744 155660
rect 378600 152040 378652 152046
rect 378600 151982 378652 151988
rect 378704 151814 378732 155654
rect 379440 151814 379468 158714
rect 380176 154086 380204 163254
rect 380452 163146 380480 163254
rect 380530 163200 380586 164400
rect 381096 163254 381308 163282
rect 380544 163146 380572 163200
rect 380452 163118 380572 163146
rect 380992 154284 381044 154290
rect 380992 154226 381044 154232
rect 380164 154080 380216 154086
rect 380164 154022 380216 154028
rect 380256 151836 380308 151842
rect 378704 151786 378916 151814
rect 379440 151786 379560 151814
rect 378888 149954 378916 151786
rect 379532 149954 379560 151786
rect 380256 151778 380308 151784
rect 380268 149954 380296 151778
rect 381004 149954 381032 154226
rect 381096 152318 381124 163254
rect 381280 163146 381308 163254
rect 381358 163200 381414 164400
rect 382186 163200 382242 164400
rect 383106 163200 383162 164400
rect 383672 163254 383884 163282
rect 381372 163146 381400 163200
rect 381280 163118 381400 163146
rect 381452 155644 381504 155650
rect 381452 155586 381504 155592
rect 381084 152312 381136 152318
rect 381084 152254 381136 152260
rect 381464 149954 381492 155586
rect 382200 153134 382228 163200
rect 383120 159390 383148 163200
rect 382740 159384 382792 159390
rect 382740 159326 382792 159332
rect 383108 159384 383160 159390
rect 383108 159326 383160 159332
rect 382372 159044 382424 159050
rect 382372 158986 382424 158992
rect 382188 153128 382240 153134
rect 382188 153070 382240 153076
rect 382384 152998 382412 158986
rect 382280 152992 382332 152998
rect 382280 152934 382332 152940
rect 382372 152992 382424 152998
rect 382372 152934 382424 152940
rect 382292 149954 382320 152934
rect 382752 149954 382780 159326
rect 383672 154222 383700 163254
rect 383856 163146 383884 163254
rect 383934 163200 383990 164400
rect 384762 163200 384818 164400
rect 385590 163200 385646 164400
rect 386418 163200 386474 164400
rect 386524 163254 387196 163282
rect 383948 163146 383976 163200
rect 383856 163118 383976 163146
rect 384776 158778 384804 163200
rect 385604 159254 385632 163200
rect 385592 159248 385644 159254
rect 385592 159190 385644 159196
rect 385408 159180 385460 159186
rect 385408 159122 385460 159128
rect 384948 158976 385000 158982
rect 384948 158918 385000 158924
rect 384764 158772 384816 158778
rect 384764 158714 384816 158720
rect 383752 154420 383804 154426
rect 383752 154362 383804 154368
rect 383660 154216 383712 154222
rect 383660 154158 383712 154164
rect 383764 150226 383792 154362
rect 384960 152114 384988 158918
rect 385132 158908 385184 158914
rect 385132 158850 385184 158856
rect 385040 152516 385092 152522
rect 385040 152458 385092 152464
rect 384948 152108 385000 152114
rect 384948 152050 385000 152056
rect 384120 152040 384172 152046
rect 384120 151982 384172 151988
rect 383764 150198 383838 150226
rect 375760 149926 376096 149954
rect 376312 149926 376740 149954
rect 377048 149926 377384 149954
rect 377600 149926 378028 149954
rect 378336 149926 378672 149954
rect 378888 149926 379316 149954
rect 379532 149926 379960 149954
rect 380268 149926 380604 149954
rect 381004 149926 381248 149954
rect 381464 149926 381892 149954
rect 382292 149926 382536 149954
rect 382752 149926 383180 149954
rect 383810 149940 383838 150198
rect 384132 149954 384160 151982
rect 385052 150226 385080 152458
rect 385144 151910 385172 158850
rect 385420 153202 385448 159122
rect 386328 158840 386380 158846
rect 386328 158782 386380 158788
rect 386052 154488 386104 154494
rect 386052 154430 386104 154436
rect 385408 153196 385460 153202
rect 385408 153138 385460 153144
rect 385408 152380 385460 152386
rect 385408 152322 385460 152328
rect 385132 151904 385184 151910
rect 385132 151846 385184 151852
rect 385052 150198 385126 150226
rect 384132 149926 384468 149954
rect 385098 149940 385126 150198
rect 385420 149954 385448 152322
rect 386064 149954 386092 154430
rect 386340 152046 386368 158782
rect 386432 152522 386460 163200
rect 386524 154290 386552 163254
rect 387168 163146 387196 163254
rect 387246 163200 387302 164400
rect 388074 163200 388130 164400
rect 388994 163200 389050 164400
rect 389822 163200 389878 164400
rect 390650 163200 390706 164400
rect 391478 163200 391534 164400
rect 392306 163200 392362 164400
rect 393134 163200 393190 164400
rect 393332 163254 393912 163282
rect 387260 163146 387288 163200
rect 387168 163118 387288 163146
rect 388088 158778 388116 163200
rect 388352 159996 388404 160002
rect 388352 159938 388404 159944
rect 388076 158772 388128 158778
rect 388076 158714 388128 158720
rect 386512 154284 386564 154290
rect 386512 154226 386564 154232
rect 387340 153196 387392 153202
rect 387340 153138 387392 153144
rect 386696 152992 386748 152998
rect 386696 152934 386748 152940
rect 386420 152516 386472 152522
rect 386420 152458 386472 152464
rect 386328 152040 386380 152046
rect 386328 151982 386380 151988
rect 386708 149954 386736 152934
rect 387352 149954 387380 153138
rect 388364 152386 388392 159938
rect 389008 159322 389036 163200
rect 389836 160002 389864 163200
rect 389824 159996 389876 160002
rect 389824 159938 389876 159944
rect 390560 159452 390612 159458
rect 390560 159394 390612 159400
rect 388996 159316 389048 159322
rect 388996 159258 389048 159264
rect 388444 159112 388496 159118
rect 388444 159054 388496 159060
rect 388352 152380 388404 152386
rect 388352 152322 388404 152328
rect 388456 152250 388484 159054
rect 389180 158840 389232 158846
rect 389180 158782 389232 158788
rect 388628 154556 388680 154562
rect 388628 154498 388680 154504
rect 387984 152244 388036 152250
rect 387984 152186 388036 152192
rect 388444 152244 388496 152250
rect 388444 152186 388496 152192
rect 387996 149954 388024 152186
rect 388640 149954 388668 154498
rect 389192 153202 389220 158782
rect 390376 158772 390428 158778
rect 390376 158714 390428 158720
rect 389180 153196 389232 153202
rect 389180 153138 389232 153144
rect 390388 152998 390416 158714
rect 390376 152992 390428 152998
rect 390376 152934 390428 152940
rect 389272 152584 389324 152590
rect 389272 152526 389324 152532
rect 389284 149954 389312 152526
rect 389916 151972 389968 151978
rect 389916 151914 389968 151920
rect 389928 149954 389956 151914
rect 390572 149954 390600 159394
rect 390664 154494 390692 163200
rect 391492 158914 391520 163200
rect 392320 159186 392348 163200
rect 392400 159520 392452 159526
rect 392400 159462 392452 159468
rect 392308 159180 392360 159186
rect 392308 159122 392360 159128
rect 391480 158908 391532 158914
rect 391480 158850 391532 158856
rect 390652 154488 390704 154494
rect 390652 154430 390704 154436
rect 391204 153876 391256 153882
rect 391204 153818 391256 153824
rect 391216 149954 391244 153818
rect 392032 152380 392084 152386
rect 392032 152322 392084 152328
rect 392044 152114 392072 152322
rect 391940 152108 391992 152114
rect 391940 152050 391992 152056
rect 392032 152108 392084 152114
rect 392032 152050 392084 152056
rect 391952 149954 391980 152050
rect 392412 149954 392440 159462
rect 393148 152590 393176 163200
rect 393332 154426 393360 163254
rect 393884 163146 393912 163254
rect 393962 163200 394018 164400
rect 394882 163200 394938 164400
rect 395710 163200 395766 164400
rect 396538 163200 396594 164400
rect 397366 163200 397422 164400
rect 397472 163254 398144 163282
rect 393976 163146 394004 163200
rect 393884 163118 394004 163146
rect 394608 158908 394660 158914
rect 394608 158850 394660 158856
rect 393320 154420 393372 154426
rect 393320 154362 393372 154368
rect 393780 153808 393832 153814
rect 393780 153750 393832 153756
rect 393320 152720 393372 152726
rect 393320 152662 393372 152668
rect 393136 152584 393188 152590
rect 393136 152526 393188 152532
rect 393332 149954 393360 152662
rect 393792 149954 393820 153750
rect 394620 152386 394648 158850
rect 394896 152726 394924 163200
rect 395436 159792 395488 159798
rect 395436 159734 395488 159740
rect 395252 159588 395304 159594
rect 395252 159530 395304 159536
rect 395068 152856 395120 152862
rect 395068 152798 395120 152804
rect 394884 152720 394936 152726
rect 394884 152662 394936 152668
rect 394608 152380 394660 152386
rect 394608 152322 394660 152328
rect 394700 151904 394752 151910
rect 394700 151846 394752 151852
rect 394712 150226 394740 151846
rect 394712 150198 394786 150226
rect 385420 149926 385756 149954
rect 386064 149926 386400 149954
rect 386708 149926 387044 149954
rect 387352 149926 387688 149954
rect 387996 149926 388332 149954
rect 388640 149926 388976 149954
rect 389284 149926 389620 149954
rect 389928 149926 390264 149954
rect 390572 149926 390908 149954
rect 391216 149926 391552 149954
rect 391952 149926 392196 149954
rect 392412 149926 392840 149954
rect 393332 149926 393484 149954
rect 393792 149926 394128 149954
rect 394758 149940 394786 150198
rect 395080 149954 395108 152798
rect 395264 151814 395292 159530
rect 395448 152862 395476 159734
rect 395724 159118 395752 163200
rect 396264 159928 396316 159934
rect 396264 159870 396316 159876
rect 395712 159112 395764 159118
rect 395712 159054 395764 159060
rect 395436 152856 395488 152862
rect 395436 152798 395488 152804
rect 396276 151910 396304 159870
rect 396552 159798 396580 163200
rect 396540 159792 396592 159798
rect 396540 159734 396592 159740
rect 397380 154358 397408 163200
rect 397368 154352 397420 154358
rect 397368 154294 397420 154300
rect 396356 153944 396408 153950
rect 396356 153886 396408 153892
rect 396264 151904 396316 151910
rect 396264 151846 396316 151852
rect 395264 151786 395660 151814
rect 395632 149954 395660 151786
rect 396368 149954 396396 153886
rect 397472 153882 397500 163254
rect 398116 163146 398144 163254
rect 398194 163200 398250 164400
rect 399022 163200 399078 164400
rect 399128 163254 399800 163282
rect 398208 163146 398236 163200
rect 398116 163118 398236 163146
rect 398104 160064 398156 160070
rect 398104 160006 398156 160012
rect 397460 153876 397512 153882
rect 397460 153818 397512 153824
rect 397552 152856 397604 152862
rect 397552 152798 397604 152804
rect 396908 152652 396960 152658
rect 396908 152594 396960 152600
rect 396920 149954 396948 152594
rect 397564 149954 397592 152798
rect 398116 151842 398144 160006
rect 399036 159594 399064 163200
rect 399024 159588 399076 159594
rect 399024 159530 399076 159536
rect 398932 159248 398984 159254
rect 398932 159190 398984 159196
rect 398840 154012 398892 154018
rect 398840 153954 398892 153960
rect 398196 152176 398248 152182
rect 398196 152118 398248 152124
rect 398104 151836 398156 151842
rect 398104 151778 398156 151784
rect 398208 149954 398236 152118
rect 398852 149954 398880 153954
rect 398944 151978 398972 159190
rect 399128 152658 399156 163254
rect 399772 163146 399800 163254
rect 399850 163200 399906 164400
rect 400770 163200 400826 164400
rect 401598 163200 401654 164400
rect 402426 163200 402482 164400
rect 403254 163200 403310 164400
rect 404082 163200 404138 164400
rect 404372 163254 404860 163282
rect 399864 163146 399892 163200
rect 399772 163118 399892 163146
rect 400680 159656 400732 159662
rect 400680 159598 400732 159604
rect 400220 152788 400272 152794
rect 400220 152730 400272 152736
rect 399116 152652 399168 152658
rect 399116 152594 399168 152600
rect 399484 152040 399536 152046
rect 399484 151982 399536 151988
rect 398932 151972 398984 151978
rect 398932 151914 398984 151920
rect 399496 149954 399524 151982
rect 400232 149954 400260 152730
rect 400692 149954 400720 159598
rect 400784 159254 400812 163200
rect 400772 159248 400824 159254
rect 400772 159190 400824 159196
rect 401612 153950 401640 163200
rect 401784 155236 401836 155242
rect 401784 155178 401836 155184
rect 401600 153944 401652 153950
rect 401600 153886 401652 153892
rect 401796 150226 401824 155178
rect 402440 152794 402468 163200
rect 403268 159934 403296 163200
rect 403256 159928 403308 159934
rect 403256 159870 403308 159876
rect 404096 159458 404124 163200
rect 404084 159452 404136 159458
rect 404084 159394 404136 159400
rect 404176 159316 404228 159322
rect 404176 159258 404228 159264
rect 403532 155304 403584 155310
rect 403532 155246 403584 155252
rect 403348 153060 403400 153066
rect 403348 153002 403400 153008
rect 402428 152788 402480 152794
rect 402428 152730 402480 152736
rect 402060 152448 402112 152454
rect 402060 152390 402112 152396
rect 401750 150198 401824 150226
rect 395080 149926 395416 149954
rect 395632 149926 396060 149954
rect 396368 149926 396612 149954
rect 396920 149926 397256 149954
rect 397564 149926 397900 149954
rect 398208 149926 398544 149954
rect 398852 149926 399188 149954
rect 399496 149926 399832 149954
rect 400232 149926 400476 149954
rect 400692 149926 401120 149954
rect 401750 149940 401778 150198
rect 402072 149954 402100 152390
rect 402980 151904 403032 151910
rect 402980 151846 403032 151852
rect 402992 150226 403020 151846
rect 402992 150198 403066 150226
rect 402072 149926 402408 149954
rect 403038 149940 403066 150198
rect 403360 149954 403388 153002
rect 403544 151814 403572 155246
rect 404188 152454 404216 159258
rect 404268 159180 404320 159186
rect 404268 159122 404320 159128
rect 404176 152448 404228 152454
rect 404176 152390 404228 152396
rect 404280 151910 404308 159122
rect 404372 153066 404400 163254
rect 404832 163146 404860 163254
rect 404910 163200 404966 164400
rect 405738 163200 405794 164400
rect 406658 163200 406714 164400
rect 407486 163200 407542 164400
rect 407684 163254 408264 163282
rect 404924 163146 404952 163200
rect 404832 163118 404952 163146
rect 405464 159112 405516 159118
rect 405464 159054 405516 159060
rect 404360 153060 404412 153066
rect 404360 153002 404412 153008
rect 405280 152924 405332 152930
rect 405280 152866 405332 152872
rect 404636 152108 404688 152114
rect 404636 152050 404688 152056
rect 404268 151904 404320 151910
rect 404268 151846 404320 151852
rect 403544 151786 403940 151814
rect 403912 149954 403940 151786
rect 404648 149954 404676 152050
rect 405292 149954 405320 152866
rect 405476 152182 405504 159054
rect 405752 158846 405780 163200
rect 405832 159860 405884 159866
rect 405832 159802 405884 159808
rect 405740 158840 405792 158846
rect 405740 158782 405792 158788
rect 405464 152176 405516 152182
rect 405464 152118 405516 152124
rect 405844 149954 405872 159802
rect 405924 159724 405976 159730
rect 405924 159666 405976 159672
rect 405936 152930 405964 159666
rect 406568 154148 406620 154154
rect 406568 154090 406620 154096
rect 405924 152924 405976 152930
rect 405924 152866 405976 152872
rect 406580 149954 406608 154090
rect 406672 152862 406700 163200
rect 407500 159662 407528 163200
rect 407488 159656 407540 159662
rect 407488 159598 407540 159604
rect 406660 152856 406712 152862
rect 406660 152798 406712 152804
rect 407684 152425 407712 163254
rect 408236 163146 408264 163254
rect 408314 163200 408370 164400
rect 409142 163200 409198 164400
rect 409970 163200 410026 164400
rect 410798 163200 410854 164400
rect 411272 163254 411576 163282
rect 408328 163146 408356 163200
rect 408236 163118 408356 163146
rect 408592 159588 408644 159594
rect 408592 159530 408644 159536
rect 408500 152924 408552 152930
rect 408500 152866 408552 152872
rect 407948 152448 408000 152454
rect 407670 152416 407726 152425
rect 407948 152390 408000 152396
rect 407670 152351 407726 152360
rect 407212 152244 407264 152250
rect 407212 152186 407264 152192
rect 407224 149954 407252 152186
rect 407960 151910 407988 152390
rect 407948 151904 408000 151910
rect 407948 151846 408000 151852
rect 407856 151836 407908 151842
rect 407856 151778 407908 151784
rect 407868 149954 407896 151778
rect 408512 149954 408540 152866
rect 408604 151978 408632 159530
rect 409156 158982 409184 163200
rect 409984 160070 410012 163200
rect 409972 160064 410024 160070
rect 409972 160006 410024 160012
rect 410812 159594 410840 163200
rect 410800 159588 410852 159594
rect 410800 159530 410852 159536
rect 409144 158976 409196 158982
rect 409144 158918 409196 158924
rect 410892 158976 410944 158982
rect 410892 158918 410944 158924
rect 409236 158840 409288 158846
rect 409236 158782 409288 158788
rect 409144 154080 409196 154086
rect 409144 154022 409196 154028
rect 408592 151972 408644 151978
rect 408592 151914 408644 151920
rect 409156 149954 409184 154022
rect 409248 152250 409276 158782
rect 410432 153128 410484 153134
rect 410432 153070 410484 153076
rect 409880 152312 409932 152318
rect 409880 152254 409932 152260
rect 409236 152244 409288 152250
rect 409236 152186 409288 152192
rect 409892 149954 409920 152254
rect 410444 149954 410472 153070
rect 410904 152454 410932 158918
rect 411272 152930 411300 163254
rect 411548 163146 411576 163254
rect 411626 163200 411682 164400
rect 412546 163200 412602 164400
rect 413374 163200 413430 164400
rect 414202 163200 414258 164400
rect 414308 163254 414980 163282
rect 411640 163146 411668 163200
rect 411548 163118 411668 163146
rect 411352 159384 411404 159390
rect 411352 159326 411404 159332
rect 411260 152924 411312 152930
rect 411260 152866 411312 152872
rect 410892 152448 410944 152454
rect 410892 152390 410944 152396
rect 411364 150226 411392 159326
rect 412560 158914 412588 163200
rect 413388 158982 413416 163200
rect 413928 159996 413980 160002
rect 413928 159938 413980 159944
rect 413836 159792 413888 159798
rect 413836 159734 413888 159740
rect 413376 158976 413428 158982
rect 413376 158918 413428 158924
rect 412548 158908 412600 158914
rect 412548 158850 412600 158856
rect 413100 158908 413152 158914
rect 413100 158850 413152 158856
rect 411720 154216 411772 154222
rect 411720 154158 411772 154164
rect 411364 150198 411438 150226
rect 403360 149926 403696 149954
rect 403912 149926 404340 149954
rect 404648 149926 404984 149954
rect 405292 149926 405628 149954
rect 405844 149926 406272 149954
rect 406580 149926 406916 149954
rect 407224 149926 407560 149954
rect 407868 149926 408204 149954
rect 408512 149926 408848 149954
rect 409156 149926 409492 149954
rect 409892 149926 410136 149954
rect 410444 149926 410780 149954
rect 411410 149940 411438 150198
rect 411732 149954 411760 154158
rect 413112 153202 413140 158850
rect 412640 153196 412692 153202
rect 412640 153138 412692 153144
rect 413100 153196 413152 153202
rect 413100 153138 413152 153144
rect 412652 150226 412680 153138
rect 413652 152516 413704 152522
rect 413652 152458 413704 152464
rect 412916 152312 412968 152318
rect 412744 152272 412916 152300
rect 412744 152182 412772 152272
rect 412916 152254 412968 152260
rect 412732 152176 412784 152182
rect 412732 152118 412784 152124
rect 413008 152176 413060 152182
rect 413008 152118 413060 152124
rect 412652 150198 412726 150226
rect 411732 149926 412068 149954
rect 412698 149940 412726 150198
rect 413020 149954 413048 152118
rect 413560 152040 413612 152046
rect 413560 151982 413612 151988
rect 413572 151842 413600 151982
rect 413560 151836 413612 151842
rect 413560 151778 413612 151784
rect 413664 149954 413692 152458
rect 413848 151978 413876 159734
rect 413940 152182 413968 159938
rect 414216 159730 414244 163200
rect 414204 159724 414256 159730
rect 414204 159666 414256 159672
rect 414204 154284 414256 154290
rect 414204 154226 414256 154232
rect 413928 152176 413980 152182
rect 413928 152118 413980 152124
rect 413836 151972 413888 151978
rect 413836 151914 413888 151920
rect 414216 149954 414244 154226
rect 414308 153134 414336 163254
rect 414952 163146 414980 163254
rect 415030 163200 415086 164400
rect 415412 163254 415808 163282
rect 415044 163146 415072 163200
rect 414952 163118 415072 163146
rect 414296 153128 414348 153134
rect 414296 153070 414348 153076
rect 414940 152992 414992 152998
rect 414940 152934 414992 152940
rect 414952 149954 414980 152934
rect 415412 152522 415440 163254
rect 415780 163146 415808 163254
rect 415858 163200 415914 164400
rect 416686 163200 416742 164400
rect 417514 163200 417570 164400
rect 418172 163254 418384 163282
rect 415872 163146 415900 163200
rect 415780 163118 415900 163146
rect 416596 159928 416648 159934
rect 416596 159870 416648 159876
rect 415400 152516 415452 152522
rect 415400 152458 415452 152464
rect 416608 152182 416636 159870
rect 416700 158846 416728 163200
rect 417528 159390 417556 163200
rect 417608 160064 417660 160070
rect 417608 160006 417660 160012
rect 417516 159384 417568 159390
rect 417516 159326 417568 159332
rect 416688 158840 416740 158846
rect 416688 158782 416740 158788
rect 416872 154488 416924 154494
rect 416872 154430 416924 154436
rect 416228 152176 416280 152182
rect 416228 152118 416280 152124
rect 416596 152176 416648 152182
rect 416596 152118 416648 152124
rect 415676 151904 415728 151910
rect 415676 151846 415728 151852
rect 415688 149954 415716 151846
rect 416240 149954 416268 152118
rect 416884 149954 416912 154430
rect 417424 152652 417476 152658
rect 417424 152594 417476 152600
rect 417436 151842 417464 152594
rect 417620 152386 417648 160006
rect 418172 152998 418200 163254
rect 418356 163146 418384 163254
rect 418434 163200 418490 164400
rect 418632 163254 419212 163282
rect 418448 163146 418476 163200
rect 418356 163118 418476 163146
rect 418160 152992 418212 152998
rect 418160 152934 418212 152940
rect 418632 152658 418660 163254
rect 419184 163146 419212 163254
rect 419262 163200 419318 164400
rect 420090 163200 420146 164400
rect 420918 163200 420974 164400
rect 421024 163254 421696 163282
rect 419276 163146 419304 163200
rect 419184 163118 419304 163146
rect 419724 158976 419776 158982
rect 419724 158918 419776 158924
rect 419632 158840 419684 158846
rect 419632 158782 419684 158788
rect 419540 154420 419592 154426
rect 419540 154362 419592 154368
rect 418620 152652 418672 152658
rect 418620 152594 418672 152600
rect 418804 152584 418856 152590
rect 418804 152526 418856 152532
rect 418896 152584 418948 152590
rect 418896 152526 418948 152532
rect 417516 152380 417568 152386
rect 417516 152322 417568 152328
rect 417608 152380 417660 152386
rect 417608 152322 417660 152328
rect 417424 151836 417476 151842
rect 417424 151778 417476 151784
rect 417528 149954 417556 152322
rect 418160 151904 418212 151910
rect 418160 151846 418212 151852
rect 418172 149954 418200 151846
rect 418816 149954 418844 152526
rect 418908 152386 418936 152526
rect 418896 152380 418948 152386
rect 418896 152322 418948 152328
rect 419552 149954 419580 154362
rect 419644 151910 419672 158782
rect 419736 152046 419764 158918
rect 420104 158914 420132 163200
rect 420932 159798 420960 163200
rect 420920 159792 420972 159798
rect 420920 159734 420972 159740
rect 420092 158908 420144 158914
rect 420092 158850 420144 158856
rect 421024 152726 421052 163254
rect 421668 163146 421696 163254
rect 421746 163200 421802 164400
rect 422312 163254 422524 163282
rect 421760 163146 421788 163200
rect 421668 163118 421788 163146
rect 420092 152720 420144 152726
rect 420092 152662 420144 152668
rect 421012 152720 421064 152726
rect 421012 152662 421064 152668
rect 419724 152040 419776 152046
rect 419724 151982 419776 151988
rect 419632 151904 419684 151910
rect 419632 151846 419684 151852
rect 420104 149954 420132 152662
rect 422312 152318 422340 163254
rect 422496 163146 422524 163254
rect 422574 163200 422630 164400
rect 422772 163254 423352 163282
rect 422588 163146 422616 163200
rect 422496 163118 422616 163146
rect 422484 154352 422536 154358
rect 422484 154294 422536 154300
rect 420920 152312 420972 152318
rect 420920 152254 420972 152260
rect 422300 152312 422352 152318
rect 422300 152254 422352 152260
rect 420932 149954 420960 152254
rect 421380 151972 421432 151978
rect 421380 151914 421432 151920
rect 421392 149954 421420 151914
rect 422496 149954 422524 154294
rect 422668 153876 422720 153882
rect 422668 153818 422720 153824
rect 413020 149926 413356 149954
rect 413664 149926 414000 149954
rect 414216 149926 414644 149954
rect 414952 149926 415288 149954
rect 415688 149926 415932 149954
rect 416240 149926 416576 149954
rect 416884 149926 417220 149954
rect 417528 149926 417864 149954
rect 418172 149926 418508 149954
rect 418816 149926 419152 149954
rect 419552 149926 419796 149954
rect 420104 149926 420440 149954
rect 420932 149926 421084 149954
rect 421392 149926 421728 149954
rect 422372 149926 422524 149954
rect 422680 149954 422708 153818
rect 422772 151978 422800 163254
rect 423324 163146 423352 163254
rect 423402 163200 423458 164400
rect 424322 163200 424378 164400
rect 425150 163200 425206 164400
rect 425978 163200 426034 164400
rect 426452 163254 426756 163282
rect 423416 163146 423444 163200
rect 423324 163118 423444 163146
rect 424336 159526 424364 163200
rect 424324 159520 424376 159526
rect 424324 159462 424376 159468
rect 424508 159248 424560 159254
rect 424508 159190 424560 159196
rect 423588 158908 423640 158914
rect 423588 158850 423640 158856
rect 423600 153270 423628 158850
rect 423588 153264 423640 153270
rect 423588 153206 423640 153212
rect 424048 152312 424100 152318
rect 424048 152254 424100 152260
rect 423312 152108 423364 152114
rect 423312 152050 423364 152056
rect 422760 151972 422812 151978
rect 422760 151914 422812 151920
rect 423324 149954 423352 152050
rect 424060 151842 424088 152254
rect 423956 151836 424008 151842
rect 423956 151778 424008 151784
rect 424048 151836 424100 151842
rect 424048 151778 424100 151784
rect 423968 149954 423996 151778
rect 424520 149954 424548 159190
rect 425164 152318 425192 163200
rect 425336 153944 425388 153950
rect 425336 153886 425388 153892
rect 425152 152312 425204 152318
rect 425152 152254 425204 152260
rect 425348 149954 425376 153886
rect 425888 152788 425940 152794
rect 425888 152730 425940 152736
rect 425900 149954 425928 152730
rect 425992 152114 426020 163200
rect 426452 152794 426480 163254
rect 426728 163146 426756 163254
rect 426806 163200 426862 164400
rect 427634 163200 427690 164400
rect 427832 163254 428412 163282
rect 426820 163146 426848 163200
rect 426728 163118 426848 163146
rect 427648 159458 427676 163200
rect 426992 159452 427044 159458
rect 426992 159394 427044 159400
rect 427636 159452 427688 159458
rect 427636 159394 427688 159400
rect 426440 152788 426492 152794
rect 426440 152730 426492 152736
rect 426900 152584 426952 152590
rect 426900 152526 426952 152532
rect 426912 152386 426940 152526
rect 426900 152380 426952 152386
rect 426900 152322 426952 152328
rect 426532 152176 426584 152182
rect 426532 152118 426584 152124
rect 425980 152108 426032 152114
rect 425980 152050 426032 152056
rect 426544 149954 426572 152118
rect 427004 149954 427032 159394
rect 427832 153814 427860 163254
rect 428384 163146 428412 163254
rect 428462 163200 428518 164400
rect 429290 163200 429346 164400
rect 429396 163254 430160 163282
rect 428476 163146 428504 163200
rect 428384 163118 428504 163146
rect 427820 153808 427872 153814
rect 427820 153750 427872 153756
rect 428004 153264 428056 153270
rect 428004 153206 428056 153212
rect 427912 153060 427964 153066
rect 427912 153002 427964 153008
rect 427726 152688 427782 152697
rect 427726 152623 427728 152632
rect 427780 152623 427782 152632
rect 427728 152594 427780 152600
rect 427096 152114 427492 152130
rect 427096 152108 427504 152114
rect 427096 152102 427452 152108
rect 427096 152046 427124 152102
rect 427452 152050 427504 152056
rect 427084 152040 427136 152046
rect 427084 151982 427136 151988
rect 427924 149954 427952 153002
rect 428016 152182 428044 153206
rect 429200 152856 429252 152862
rect 429200 152798 429252 152804
rect 428372 152244 428424 152250
rect 428372 152186 428424 152192
rect 428004 152176 428056 152182
rect 428004 152118 428056 152124
rect 428384 149954 428412 152186
rect 429212 149954 429240 152798
rect 429304 152182 429332 163200
rect 429396 152862 429424 163254
rect 430132 163146 430160 163254
rect 430210 163200 430266 164400
rect 430684 163254 430988 163282
rect 430224 163146 430252 163200
rect 430132 163118 430252 163146
rect 429568 159656 429620 159662
rect 429568 159598 429620 159604
rect 429384 152856 429436 152862
rect 429384 152798 429436 152804
rect 429292 152176 429344 152182
rect 429292 152118 429344 152124
rect 429580 149954 429608 159598
rect 430684 153134 430712 163254
rect 430960 163146 430988 163254
rect 431038 163200 431094 164400
rect 431236 163254 431816 163282
rect 431052 163146 431080 163200
rect 430960 163118 431080 163146
rect 430672 153128 430724 153134
rect 430672 153070 430724 153076
rect 431236 152561 431264 163254
rect 431788 163146 431816 163254
rect 431866 163200 431922 164400
rect 431972 163254 432644 163282
rect 431880 163146 431908 163200
rect 431788 163118 431908 163146
rect 431972 153066 432000 163254
rect 432616 163146 432644 163254
rect 432694 163200 432750 164400
rect 433522 163200 433578 164400
rect 434350 163200 434406 164400
rect 434732 163254 435128 163282
rect 432708 163146 432736 163200
rect 432616 163118 432736 163146
rect 432144 159588 432196 159594
rect 432144 159530 432196 159536
rect 431868 153060 431920 153066
rect 431868 153002 431920 153008
rect 431960 153060 432012 153066
rect 431960 153002 432012 153008
rect 431222 152552 431278 152561
rect 430856 152516 430908 152522
rect 431222 152487 431278 152496
rect 430856 152458 430908 152464
rect 430868 152425 430896 152458
rect 430948 152448 431000 152454
rect 430302 152416 430358 152425
rect 430302 152351 430358 152360
rect 430854 152416 430910 152425
rect 430948 152390 431000 152396
rect 430854 152351 430910 152360
rect 422680 149926 423016 149954
rect 423324 149926 423660 149954
rect 423968 149926 424304 149954
rect 424520 149926 424948 149954
rect 425348 149926 425592 149954
rect 425900 149926 426236 149954
rect 426544 149926 426880 149954
rect 427004 149926 427432 149954
rect 427924 149926 428076 149954
rect 428384 149926 428720 149954
rect 429212 149926 429364 149954
rect 429580 149926 430008 149954
rect 200192 149790 200344 149818
rect 430316 149818 430344 152351
rect 430960 149954 430988 152390
rect 431880 152386 431908 153002
rect 431592 152380 431644 152386
rect 431592 152322 431644 152328
rect 431868 152380 431920 152386
rect 431868 152322 431920 152328
rect 431604 149954 431632 152322
rect 432156 149954 432184 159530
rect 432696 153808 432748 153814
rect 432696 153750 432748 153756
rect 432604 152924 432656 152930
rect 432604 152866 432656 152872
rect 432616 152538 432644 152866
rect 432708 152658 432736 153750
rect 433536 153202 433564 163200
rect 433432 153196 433484 153202
rect 433432 153138 433484 153144
rect 433524 153196 433576 153202
rect 433524 153138 433576 153144
rect 432880 152992 432932 152998
rect 432880 152934 432932 152940
rect 432892 152726 432920 152934
rect 432880 152720 432932 152726
rect 432880 152662 432932 152668
rect 432970 152688 433026 152697
rect 432696 152652 432748 152658
rect 432970 152623 433026 152632
rect 432696 152594 432748 152600
rect 432984 152590 433012 152623
rect 432972 152584 433024 152590
rect 432616 152510 432828 152538
rect 432972 152526 433024 152532
rect 432512 152380 432564 152386
rect 432512 152322 432564 152328
rect 432604 152380 432656 152386
rect 432604 152322 432656 152328
rect 432420 152312 432472 152318
rect 432418 152280 432420 152289
rect 432472 152280 432474 152289
rect 432418 152215 432474 152224
rect 432326 152144 432382 152153
rect 432326 152079 432382 152088
rect 432420 152108 432472 152114
rect 432340 152046 432368 152079
rect 432420 152050 432472 152056
rect 432328 152040 432380 152046
rect 432328 151982 432380 151988
rect 432432 151774 432460 152050
rect 432524 151858 432552 152322
rect 432616 151978 432644 152322
rect 432604 151972 432656 151978
rect 432604 151914 432656 151920
rect 432696 151972 432748 151978
rect 432696 151914 432748 151920
rect 432708 151858 432736 151914
rect 432524 151830 432736 151858
rect 432420 151768 432472 151774
rect 432420 151710 432472 151716
rect 432800 149954 432828 152510
rect 433062 152416 433118 152425
rect 433062 152351 433118 152360
rect 432878 152280 432934 152289
rect 433076 152250 433104 152351
rect 432878 152215 432934 152224
rect 433064 152244 433116 152250
rect 432892 152046 432920 152215
rect 433064 152186 433116 152192
rect 432972 152176 433024 152182
rect 432970 152144 432972 152153
rect 433024 152144 433026 152153
rect 432970 152079 433026 152088
rect 432880 152040 432932 152046
rect 432880 151982 432932 151988
rect 433444 149954 433472 153138
rect 434364 152930 434392 163200
rect 434352 152924 434404 152930
rect 434352 152866 434404 152872
rect 434732 152454 434760 163254
rect 435100 163146 435128 163254
rect 435178 163200 435234 164400
rect 436098 163200 436154 164400
rect 436926 163200 436982 164400
rect 437754 163200 437810 164400
rect 438582 163200 438638 164400
rect 438872 163254 439360 163282
rect 435192 163146 435220 163200
rect 435100 163118 435220 163146
rect 434812 159724 434864 159730
rect 434812 159666 434864 159672
rect 434720 152448 434772 152454
rect 434720 152390 434772 152396
rect 434168 151768 434220 151774
rect 434168 151710 434220 151716
rect 434180 149954 434208 151710
rect 434824 149954 434852 159666
rect 436112 152318 436140 163200
rect 436940 153134 436968 163200
rect 437664 159384 437716 159390
rect 437664 159326 437716 159332
rect 436284 153128 436336 153134
rect 436284 153070 436336 153076
rect 436928 153128 436980 153134
rect 436928 153070 436980 153076
rect 435548 152312 435600 152318
rect 435548 152254 435600 152260
rect 436100 152312 436152 152318
rect 436100 152254 436152 152260
rect 435560 151978 435588 152254
rect 436296 152250 436324 153070
rect 436192 152244 436244 152250
rect 436192 152186 436244 152192
rect 436284 152244 436336 152250
rect 436284 152186 436336 152192
rect 435456 151972 435508 151978
rect 435456 151914 435508 151920
rect 435548 151972 435600 151978
rect 435548 151914 435600 151920
rect 435468 149954 435496 151914
rect 436204 149954 436232 152186
rect 436744 151904 436796 151910
rect 436744 151846 436796 151852
rect 436756 149954 436784 151846
rect 437676 150226 437704 159326
rect 437768 151842 437796 163200
rect 438032 152720 438084 152726
rect 438032 152662 438084 152668
rect 438124 152720 438176 152726
rect 438124 152662 438176 152668
rect 437756 151836 437808 151842
rect 437756 151778 437808 151784
rect 437676 150198 437750 150226
rect 430960 149926 431296 149954
rect 431604 149926 431940 149954
rect 432156 149926 432584 149954
rect 432800 149926 433228 149954
rect 433444 149926 433872 149954
rect 434180 149926 434516 149954
rect 434824 149926 435160 149954
rect 435468 149926 435804 149954
rect 436204 149926 436448 149954
rect 436756 149926 437092 149954
rect 437722 149940 437750 150198
rect 438044 149954 438072 152662
rect 438136 152522 438164 152662
rect 438596 152522 438624 163200
rect 438872 152998 438900 163254
rect 439332 163146 439360 163254
rect 439410 163200 439466 164400
rect 440238 163200 440294 164400
rect 440344 163254 441016 163282
rect 439424 163146 439452 163200
rect 439332 163118 439452 163146
rect 438860 152992 438912 152998
rect 438860 152934 438912 152940
rect 438780 152658 439084 152674
rect 438768 152652 439096 152658
rect 438820 152646 439044 152652
rect 438768 152594 438820 152600
rect 439044 152594 439096 152600
rect 438860 152584 438912 152590
rect 438860 152526 438912 152532
rect 438124 152516 438176 152522
rect 438124 152458 438176 152464
rect 438584 152516 438636 152522
rect 438584 152458 438636 152464
rect 438872 149954 438900 152526
rect 440252 151978 440280 163200
rect 440344 152726 440372 163254
rect 440988 163146 441016 163254
rect 441066 163200 441122 164400
rect 441724 163254 441936 163282
rect 441080 163146 441108 163200
rect 440988 163118 441108 163146
rect 440424 159792 440476 159798
rect 440424 159734 440476 159740
rect 440332 152720 440384 152726
rect 440332 152662 440384 152668
rect 439320 151972 439372 151978
rect 439320 151914 439372 151920
rect 440240 151972 440292 151978
rect 440240 151914 440292 151920
rect 439332 149954 439360 151914
rect 440436 149954 440464 159734
rect 441620 153400 441672 153406
rect 441620 153342 441672 153348
rect 441632 152930 441660 153342
rect 441724 152930 441752 163254
rect 441908 163146 441936 163254
rect 441986 163200 442042 164400
rect 442814 163200 442870 164400
rect 443012 163254 443592 163282
rect 442000 163146 442028 163200
rect 441908 163118 442028 163146
rect 442448 159520 442500 159526
rect 442448 159462 442500 159468
rect 441804 153196 441856 153202
rect 441804 153138 441856 153144
rect 441620 152924 441672 152930
rect 441620 152866 441672 152872
rect 441712 152924 441764 152930
rect 441712 152866 441764 152872
rect 440608 152584 440660 152590
rect 440608 152526 440660 152532
rect 438044 149926 438380 149954
rect 438872 149926 439024 149954
rect 439332 149926 439668 149954
rect 440312 149926 440464 149954
rect 440620 149954 440648 152526
rect 441816 151910 441844 153138
rect 441896 152380 441948 152386
rect 441896 152322 441948 152328
rect 441252 151904 441304 151910
rect 441252 151846 441304 151852
rect 441804 151904 441856 151910
rect 441804 151846 441856 151852
rect 441264 149954 441292 151846
rect 441908 149954 441936 152322
rect 442460 149954 442488 159462
rect 442828 152590 442856 163200
rect 443012 153202 443040 163254
rect 443564 163146 443592 163254
rect 443642 163200 443698 164400
rect 444470 163200 444526 164400
rect 445298 163200 445354 164400
rect 446126 163200 446182 164400
rect 446324 163254 446904 163282
rect 443656 163146 443684 163200
rect 443564 163118 443684 163146
rect 443000 153196 443052 153202
rect 443000 153138 443052 153144
rect 443920 153196 443972 153202
rect 443920 153138 443972 153144
rect 442816 152584 442868 152590
rect 442816 152526 442868 152532
rect 443932 152182 443960 153138
rect 443828 152176 443880 152182
rect 443828 152118 443880 152124
rect 443920 152176 443972 152182
rect 443920 152118 443972 152124
rect 443184 152040 443236 152046
rect 443184 151982 443236 151988
rect 443196 149954 443224 151982
rect 443840 149954 443868 152118
rect 444484 152046 444512 163200
rect 445024 159452 445076 159458
rect 445024 159394 445076 159400
rect 444564 152788 444616 152794
rect 444564 152730 444616 152736
rect 444472 152040 444524 152046
rect 444472 151982 444524 151988
rect 444576 149954 444604 152730
rect 445036 149954 445064 159394
rect 445312 152386 445340 163200
rect 446140 159730 446168 163200
rect 446128 159724 446180 159730
rect 446128 159666 446180 159672
rect 446324 152794 446352 163254
rect 446876 163146 446904 163254
rect 446954 163200 447010 164400
rect 447874 163200 447930 164400
rect 448702 163200 448758 164400
rect 449530 163200 449586 164400
rect 450358 163200 450414 164400
rect 451186 163200 451242 164400
rect 452014 163200 452070 164400
rect 452842 163200 452898 164400
rect 453762 163200 453818 164400
rect 454590 163200 454646 164400
rect 455418 163200 455474 164400
rect 456246 163200 456302 164400
rect 457074 163200 457130 164400
rect 457902 163200 457958 164400
rect 458730 163200 458786 164400
rect 459650 163200 459706 164400
rect 460478 163200 460534 164400
rect 461306 163200 461362 164400
rect 462134 163200 462190 164400
rect 462962 163200 463018 164400
rect 463790 163200 463846 164400
rect 464618 163200 464674 164400
rect 465538 163200 465594 164400
rect 466366 163200 466422 164400
rect 467194 163200 467250 164400
rect 468022 163200 468078 164400
rect 468850 163200 468906 164400
rect 469678 163200 469734 164400
rect 470506 163200 470562 164400
rect 471426 163200 471482 164400
rect 472254 163200 472310 164400
rect 473082 163200 473138 164400
rect 473910 163200 473966 164400
rect 474738 163200 474794 164400
rect 475566 163200 475622 164400
rect 476394 163200 476450 164400
rect 477314 163200 477370 164400
rect 478142 163200 478198 164400
rect 478970 163200 479026 164400
rect 479798 163200 479854 164400
rect 480626 163200 480682 164400
rect 481454 163200 481510 164400
rect 482282 163200 482338 164400
rect 483202 163200 483258 164400
rect 484030 163200 484086 164400
rect 484504 163254 484808 163282
rect 446968 163146 446996 163200
rect 446876 163118 446996 163146
rect 447888 159458 447916 163200
rect 447876 159452 447928 159458
rect 447876 159394 447928 159400
rect 448716 159390 448744 163200
rect 449544 159866 449572 163200
rect 449532 159860 449584 159866
rect 449532 159802 449584 159808
rect 450372 159662 450400 163200
rect 450360 159656 450412 159662
rect 450360 159598 450412 159604
rect 451200 159594 451228 163200
rect 451188 159588 451240 159594
rect 451188 159530 451240 159536
rect 452028 159526 452056 163200
rect 452856 160002 452884 163200
rect 452844 159996 452896 160002
rect 452844 159938 452896 159944
rect 453776 159798 453804 163200
rect 454604 160070 454632 163200
rect 454592 160064 454644 160070
rect 454592 160006 454644 160012
rect 455432 159934 455460 163200
rect 455420 159928 455472 159934
rect 455420 159870 455472 159876
rect 453764 159792 453816 159798
rect 453764 159734 453816 159740
rect 452016 159520 452068 159526
rect 452016 159462 452068 159468
rect 448704 159384 448756 159390
rect 448704 159326 448756 159332
rect 456260 159186 456288 163200
rect 456800 159724 456852 159730
rect 456800 159666 456852 159672
rect 456248 159180 456300 159186
rect 456248 159122 456300 159128
rect 456812 153202 456840 159666
rect 457088 159254 457116 163200
rect 457916 159322 457944 163200
rect 458744 159730 458772 163200
rect 459560 159860 459612 159866
rect 459560 159802 459612 159808
rect 458732 159724 458784 159730
rect 458732 159666 458784 159672
rect 457904 159316 457956 159322
rect 457904 159258 457956 159264
rect 457076 159248 457128 159254
rect 457076 159190 457128 159196
rect 450268 153196 450320 153202
rect 450268 153138 450320 153144
rect 456800 153196 456852 153202
rect 456800 153138 456852 153144
rect 459192 153196 459244 153202
rect 459192 153138 459244 153144
rect 448980 153060 449032 153066
rect 448980 153002 449032 153008
rect 447876 152924 447928 152930
rect 447876 152866 447928 152872
rect 447140 152856 447192 152862
rect 447140 152798 447192 152804
rect 446312 152788 446364 152794
rect 446312 152730 446364 152736
rect 445760 152652 445812 152658
rect 445760 152594 445812 152600
rect 445300 152380 445352 152386
rect 445300 152322 445352 152328
rect 445772 149954 445800 152594
rect 446496 152312 446548 152318
rect 446232 152238 446444 152266
rect 446496 152254 446548 152260
rect 446232 151910 446260 152238
rect 446416 152114 446444 152238
rect 446312 152108 446364 152114
rect 446312 152050 446364 152056
rect 446404 152108 446456 152114
rect 446404 152050 446456 152056
rect 446220 151904 446272 151910
rect 446220 151846 446272 151852
rect 446324 149954 446352 152050
rect 446508 151910 446536 152254
rect 446496 151904 446548 151910
rect 446496 151846 446548 151852
rect 447152 149954 447180 152798
rect 447692 152244 447744 152250
rect 447692 152186 447744 152192
rect 447704 149954 447732 152186
rect 447888 152182 447916 152866
rect 448518 152552 448574 152561
rect 448518 152487 448574 152496
rect 447876 152176 447928 152182
rect 447876 152118 447928 152124
rect 448532 149954 448560 152487
rect 448992 149954 449020 153002
rect 449900 152108 449952 152114
rect 449900 152050 449952 152056
rect 449912 150226 449940 152050
rect 449912 150198 449986 150226
rect 440620 149926 440956 149954
rect 441264 149926 441600 149954
rect 441908 149926 442244 149954
rect 442460 149926 442888 149954
rect 443196 149926 443532 149954
rect 443840 149926 444176 149954
rect 444576 149926 444820 149954
rect 445036 149926 445464 149954
rect 445772 149926 446108 149954
rect 446324 149926 446752 149954
rect 447152 149926 447396 149954
rect 447704 149926 448040 149954
rect 448532 149926 448684 149954
rect 448992 149926 449328 149954
rect 449958 149940 449986 150198
rect 450280 149954 450308 153138
rect 452200 153128 452252 153134
rect 452200 153070 452252 153076
rect 450912 152448 450964 152454
rect 450912 152390 450964 152396
rect 450924 149954 450952 152390
rect 451556 151904 451608 151910
rect 451556 151846 451608 151852
rect 451568 149954 451596 151846
rect 452212 149954 452240 153070
rect 454224 152992 454276 152998
rect 454224 152934 454276 152940
rect 453488 152516 453540 152522
rect 453488 152458 453540 152464
rect 452844 151836 452896 151842
rect 452844 151778 452896 151784
rect 452856 149954 452884 151778
rect 453500 149954 453528 152458
rect 454236 149954 454264 152934
rect 455420 152720 455472 152726
rect 455420 152662 455472 152668
rect 454776 151972 454828 151978
rect 454776 151914 454828 151920
rect 454788 149954 454816 151914
rect 455432 149954 455460 152662
rect 456800 152584 456852 152590
rect 456800 152526 456852 152532
rect 456064 152176 456116 152182
rect 456064 152118 456116 152124
rect 456076 149954 456104 152118
rect 456812 149954 456840 152526
rect 458548 152380 458600 152386
rect 458548 152322 458600 152328
rect 457352 152312 457404 152318
rect 457352 152254 457404 152260
rect 457364 149954 457392 152254
rect 458180 152040 458232 152046
rect 458180 151982 458232 151988
rect 458192 150226 458220 151982
rect 458192 150198 458266 150226
rect 450280 149926 450616 149954
rect 450924 149926 451260 149954
rect 451568 149926 451904 149954
rect 452212 149926 452548 149954
rect 452856 149926 453192 149954
rect 453500 149926 453836 149954
rect 454236 149926 454480 149954
rect 454788 149926 455124 149954
rect 455432 149926 455768 149954
rect 456076 149926 456412 149954
rect 456812 149926 457056 149954
rect 457364 149926 457700 149954
rect 458238 149940 458266 150198
rect 458560 149954 458588 152322
rect 459204 149954 459232 153138
rect 459572 152046 459600 159802
rect 459664 159050 459692 163200
rect 460112 159452 460164 159458
rect 460112 159394 460164 159400
rect 459652 159044 459704 159050
rect 459652 158986 459704 158992
rect 459836 152788 459888 152794
rect 459836 152730 459888 152736
rect 459560 152040 459612 152046
rect 459560 151982 459612 151988
rect 459848 149954 459876 152730
rect 460124 151814 460152 159394
rect 460492 159118 460520 163200
rect 461320 159390 461348 163200
rect 461492 159588 461544 159594
rect 461492 159530 461544 159536
rect 461216 159384 461268 159390
rect 461216 159326 461268 159332
rect 461308 159384 461360 159390
rect 461308 159326 461360 159332
rect 460480 159112 460532 159118
rect 460480 159054 460532 159060
rect 460124 151786 460428 151814
rect 460400 149954 460428 151786
rect 461228 149954 461256 159326
rect 461504 153202 461532 159530
rect 462148 158982 462176 163200
rect 462228 159656 462280 159662
rect 462228 159598 462280 159604
rect 462136 158976 462188 158982
rect 462136 158918 462188 158924
rect 461492 153196 461544 153202
rect 461492 153138 461544 153144
rect 461768 152040 461820 152046
rect 461768 151982 461820 151988
rect 461780 149954 461808 151982
rect 462240 151814 462268 159598
rect 462976 158914 463004 163200
rect 463804 159594 463832 163200
rect 464252 159996 464304 160002
rect 464252 159938 464304 159944
rect 463792 159588 463844 159594
rect 463792 159530 463844 159536
rect 463608 159520 463660 159526
rect 463608 159462 463660 159468
rect 462964 158908 463016 158914
rect 462964 158850 463016 158856
rect 463056 153196 463108 153202
rect 463056 153138 463108 153144
rect 462240 151786 462360 151814
rect 462332 149954 462360 151786
rect 463068 149954 463096 153138
rect 463620 151814 463648 159462
rect 463620 151786 463740 151814
rect 463712 149954 463740 151786
rect 464264 149954 464292 159938
rect 464632 158778 464660 163200
rect 465448 160064 465500 160070
rect 465448 160006 465500 160012
rect 464988 159792 465040 159798
rect 464988 159734 465040 159740
rect 464620 158772 464672 158778
rect 464620 158714 464672 158720
rect 465000 151814 465028 159734
rect 465080 159724 465132 159730
rect 465080 159666 465132 159672
rect 465092 153066 465120 159666
rect 465080 153060 465132 153066
rect 465080 153002 465132 153008
rect 465460 151814 465488 160006
rect 465552 159526 465580 163200
rect 465540 159520 465592 159526
rect 465540 159462 465592 159468
rect 466380 158846 466408 163200
rect 467208 159934 467236 163200
rect 468036 160002 468064 163200
rect 468024 159996 468076 160002
rect 468024 159938 468076 159944
rect 466644 159928 466696 159934
rect 466644 159870 466696 159876
rect 467196 159928 467248 159934
rect 467196 159870 467248 159876
rect 466552 159112 466604 159118
rect 466552 159054 466604 159060
rect 466460 159044 466512 159050
rect 466460 158986 466512 158992
rect 466368 158840 466420 158846
rect 466368 158782 466420 158788
rect 466472 153202 466500 158986
rect 466460 153196 466512 153202
rect 466460 153138 466512 153144
rect 466564 153134 466592 159054
rect 466552 153128 466604 153134
rect 466552 153070 466604 153076
rect 465000 151786 465120 151814
rect 465460 151786 465580 151814
rect 465092 149954 465120 151786
rect 465552 149954 465580 151786
rect 466656 150226 466684 159870
rect 468864 159662 468892 163200
rect 468852 159656 468904 159662
rect 468852 159598 468904 159604
rect 469692 159390 469720 163200
rect 470520 159730 470548 163200
rect 470508 159724 470560 159730
rect 470508 159666 470560 159672
rect 468024 159384 468076 159390
rect 468024 159326 468076 159332
rect 469680 159384 469732 159390
rect 469680 159326 469732 159332
rect 467840 159248 467892 159254
rect 467840 159190 467892 159196
rect 466920 159180 466972 159186
rect 466920 159122 466972 159128
rect 466610 150198 466684 150226
rect 458560 149926 458896 149954
rect 459204 149926 459540 149954
rect 459848 149926 460184 149954
rect 460400 149926 460828 149954
rect 461228 149926 461472 149954
rect 461780 149926 462116 149954
rect 462332 149926 462760 149954
rect 463068 149926 463404 149954
rect 463712 149926 464048 149954
rect 464264 149926 464692 149954
rect 465092 149926 465336 149954
rect 465552 149926 465980 149954
rect 466610 149940 466638 150198
rect 466932 149954 466960 159122
rect 467852 150226 467880 159190
rect 467932 158976 467984 158982
rect 467932 158918 467984 158924
rect 467944 151842 467972 158918
rect 468036 151910 468064 159326
rect 468116 159316 468168 159322
rect 468116 159258 468168 159264
rect 468024 151904 468076 151910
rect 468024 151846 468076 151852
rect 467932 151836 467984 151842
rect 467932 151778 467984 151784
rect 467852 150198 467926 150226
rect 466932 149926 467268 149954
rect 467898 149940 467926 150198
rect 468128 149954 468156 159258
rect 471440 159118 471468 163200
rect 472268 159866 472296 163200
rect 472256 159860 472308 159866
rect 472256 159802 472308 159808
rect 471520 159588 471572 159594
rect 471520 159530 471572 159536
rect 471428 159112 471480 159118
rect 471428 159054 471480 159060
rect 469220 158908 469272 158914
rect 469220 158850 469272 158856
rect 468852 153060 468904 153066
rect 468852 153002 468904 153008
rect 468864 149954 468892 153002
rect 469232 151978 469260 158850
rect 471244 158772 471296 158778
rect 471244 158714 471296 158720
rect 471256 153202 471284 158714
rect 469496 153196 469548 153202
rect 469496 153138 469548 153144
rect 471244 153196 471296 153202
rect 471244 153138 471296 153144
rect 469220 151972 469272 151978
rect 469220 151914 469272 151920
rect 469508 149954 469536 153138
rect 471532 153134 471560 159530
rect 472256 159520 472308 159526
rect 472256 159462 472308 159468
rect 470140 153128 470192 153134
rect 470140 153070 470192 153076
rect 471520 153128 471572 153134
rect 471520 153070 471572 153076
rect 470152 149954 470180 153070
rect 472268 152998 472296 159462
rect 472440 158840 472492 158846
rect 472440 158782 472492 158788
rect 472452 153066 472480 158782
rect 473096 158778 473124 163200
rect 473360 159928 473412 159934
rect 473360 159870 473412 159876
rect 473084 158772 473136 158778
rect 473084 158714 473136 158720
rect 473372 153134 473400 159870
rect 473924 159050 473952 163200
rect 473912 159044 473964 159050
rect 473912 158986 473964 158992
rect 474752 158914 474780 163200
rect 474832 159656 474884 159662
rect 474832 159598 474884 159604
rect 474740 158908 474792 158914
rect 474740 158850 474792 158856
rect 474844 153202 474872 159598
rect 475580 158982 475608 163200
rect 476028 159996 476080 160002
rect 476028 159938 476080 159944
rect 475568 158976 475620 158982
rect 475568 158918 475620 158924
rect 473544 153196 473596 153202
rect 473544 153138 473596 153144
rect 474832 153196 474884 153202
rect 474832 153138 474884 153144
rect 472716 153128 472768 153134
rect 472716 153070 472768 153076
rect 473360 153128 473412 153134
rect 473360 153070 473412 153076
rect 472440 153060 472492 153066
rect 472440 153002 472492 153008
rect 472256 152992 472308 152998
rect 472256 152934 472308 152940
rect 472072 151972 472124 151978
rect 472072 151914 472124 151920
rect 470784 151904 470836 151910
rect 470784 151846 470836 151852
rect 470796 149954 470824 151846
rect 471428 151836 471480 151842
rect 471428 151778 471480 151784
rect 471440 149954 471468 151778
rect 472084 149954 472112 151914
rect 472728 149954 472756 153070
rect 473556 149954 473584 153138
rect 475292 153128 475344 153134
rect 475292 153070 475344 153076
rect 474740 153060 474792 153066
rect 474740 153002 474792 153008
rect 474004 152992 474056 152998
rect 474004 152934 474056 152940
rect 474016 149954 474044 152934
rect 474752 149954 474780 153002
rect 475304 149954 475332 153070
rect 476040 151814 476068 159938
rect 476120 159724 476172 159730
rect 476120 159666 476172 159672
rect 476132 153134 476160 159666
rect 476408 158846 476436 163200
rect 477328 159662 477356 163200
rect 477316 159656 477368 159662
rect 477316 159598 477368 159604
rect 478156 159390 478184 163200
rect 478984 159730 479012 163200
rect 479064 159860 479116 159866
rect 479064 159802 479116 159808
rect 478972 159724 479024 159730
rect 478972 159666 479024 159672
rect 477408 159384 477460 159390
rect 477408 159326 477460 159332
rect 478144 159384 478196 159390
rect 478144 159326 478196 159332
rect 476396 158840 476448 158846
rect 476396 158782 476448 158788
rect 476580 153196 476632 153202
rect 476580 153138 476632 153144
rect 476120 153128 476172 153134
rect 476120 153070 476172 153076
rect 476040 151786 476160 151814
rect 476132 149954 476160 151786
rect 476592 149954 476620 153138
rect 477420 151814 477448 159326
rect 478420 159112 478472 159118
rect 478420 159054 478472 159060
rect 477868 153128 477920 153134
rect 477868 153070 477920 153076
rect 477420 151786 477540 151814
rect 477512 150226 477540 151786
rect 477512 150198 477586 150226
rect 468128 149926 468556 149954
rect 468864 149926 469200 149954
rect 469508 149926 469844 149954
rect 470152 149926 470488 149954
rect 470796 149926 471132 149954
rect 471440 149926 471776 149954
rect 472084 149926 472420 149954
rect 472728 149926 473064 149954
rect 473556 149926 473708 149954
rect 474016 149926 474352 149954
rect 474752 149926 474996 149954
rect 475304 149926 475640 149954
rect 476132 149926 476284 149954
rect 476592 149926 476928 149954
rect 477558 149940 477586 150198
rect 477880 149954 477908 153070
rect 478432 149954 478460 159054
rect 479076 149954 479104 159802
rect 479812 159594 479840 163200
rect 479800 159588 479852 159594
rect 479800 159530 479852 159536
rect 480640 159050 480668 163200
rect 480352 159044 480404 159050
rect 480352 158986 480404 158992
rect 480628 159044 480680 159050
rect 480628 158986 480680 158992
rect 479708 158772 479760 158778
rect 479708 158714 479760 158720
rect 479720 149954 479748 158714
rect 480364 149954 480392 158986
rect 481088 158908 481140 158914
rect 481088 158850 481140 158856
rect 481100 149954 481128 158850
rect 481468 158778 481496 163200
rect 481732 158976 481784 158982
rect 481732 158918 481784 158924
rect 481456 158772 481508 158778
rect 481456 158714 481508 158720
rect 481744 149954 481772 158918
rect 482296 158914 482324 163200
rect 482284 158908 482336 158914
rect 482284 158850 482336 158856
rect 482376 158840 482428 158846
rect 482376 158782 482428 158788
rect 482388 149954 482416 158782
rect 483216 152998 483244 163200
rect 483296 159656 483348 159662
rect 483296 159598 483348 159604
rect 483204 152992 483256 152998
rect 483204 152934 483256 152940
rect 483308 150226 483336 159598
rect 483664 159384 483716 159390
rect 483664 159326 483716 159332
rect 483308 150198 483382 150226
rect 477880 149926 478216 149954
rect 478432 149926 478860 149954
rect 479076 149926 479504 149954
rect 479720 149926 480148 149954
rect 480364 149926 480792 149954
rect 481100 149926 481436 149954
rect 481744 149926 482080 149954
rect 482388 149926 482724 149954
rect 483354 149940 483382 150198
rect 483676 149954 483704 159326
rect 484044 153134 484072 163200
rect 484032 153128 484084 153134
rect 484032 153070 484084 153076
rect 484504 153066 484532 163254
rect 484780 163146 484808 163254
rect 484858 163200 484914 164400
rect 485686 163200 485742 164400
rect 485792 163254 486464 163282
rect 484872 163146 484900 163200
rect 484780 163118 484900 163146
rect 484676 159724 484728 159730
rect 484676 159666 484728 159672
rect 484492 153060 484544 153066
rect 484492 153002 484544 153008
rect 484688 150226 484716 159666
rect 484860 159588 484912 159594
rect 484860 159530 484912 159536
rect 484642 150198 484716 150226
rect 483676 149926 484012 149954
rect 484642 149940 484670 150198
rect 484872 149954 484900 159530
rect 485700 153202 485728 163200
rect 485688 153196 485740 153202
rect 485688 153138 485740 153144
rect 485792 152046 485820 163254
rect 486436 163146 486464 163254
rect 486514 163200 486570 164400
rect 487342 163200 487398 164400
rect 488170 163200 488226 164400
rect 488552 163254 489040 163282
rect 486528 163146 486556 163200
rect 486436 163118 486556 163146
rect 485964 159044 486016 159050
rect 485964 158986 486016 158992
rect 485780 152040 485832 152046
rect 485780 151982 485832 151988
rect 485976 150226 486004 158986
rect 487252 158908 487304 158914
rect 487252 158850 487304 158856
rect 486148 158772 486200 158778
rect 486148 158714 486200 158720
rect 485930 150198 486004 150226
rect 484872 149926 485300 149954
rect 485930 149940 485958 150198
rect 486160 149954 486188 158714
rect 487264 150226 487292 158850
rect 487356 151978 487384 163200
rect 488080 153128 488132 153134
rect 488080 153070 488132 153076
rect 487528 152992 487580 152998
rect 487528 152934 487580 152940
rect 487344 151972 487396 151978
rect 487344 151914 487396 151920
rect 487218 150198 487292 150226
rect 486160 149926 486588 149954
rect 487218 149940 487246 150198
rect 487540 149954 487568 152934
rect 488092 149954 488120 153070
rect 488184 151910 488212 163200
rect 488552 151910 488580 163254
rect 489012 163146 489040 163254
rect 489090 163200 489146 164400
rect 489918 163200 489974 164400
rect 490746 163200 490802 164400
rect 491312 163254 491524 163282
rect 489104 163146 489132 163200
rect 489012 163118 489132 163146
rect 489368 153196 489420 153202
rect 489368 153138 489420 153144
rect 488724 153060 488776 153066
rect 488724 153002 488776 153008
rect 488172 151904 488224 151910
rect 488172 151846 488224 151852
rect 488540 151904 488592 151910
rect 488540 151846 488592 151852
rect 488736 149954 488764 153002
rect 489380 149954 489408 153138
rect 489932 153134 489960 163200
rect 490760 153202 490788 163200
rect 490748 153196 490800 153202
rect 490748 153138 490800 153144
rect 489920 153128 489972 153134
rect 489920 153070 489972 153076
rect 491312 152998 491340 163254
rect 491496 163146 491524 163254
rect 491574 163200 491630 164400
rect 491680 163254 492352 163282
rect 491588 163146 491616 163200
rect 491496 163118 491616 163146
rect 491300 152992 491352 152998
rect 491300 152934 491352 152940
rect 491680 152930 491708 163254
rect 492324 163146 492352 163254
rect 492402 163200 492458 164400
rect 492692 163254 493180 163282
rect 492416 163146 492444 163200
rect 492324 163118 492444 163146
rect 492692 153066 492720 163254
rect 493152 163146 493180 163254
rect 493230 163200 493286 164400
rect 494058 163200 494114 164400
rect 494164 163254 494928 163282
rect 493244 163146 493272 163200
rect 493152 163118 493272 163146
rect 493232 153196 493284 153202
rect 493232 153138 493284 153144
rect 492772 153128 492824 153134
rect 492772 153070 492824 153076
rect 492680 153060 492732 153066
rect 492680 153002 492732 153008
rect 491668 152924 491720 152930
rect 491668 152866 491720 152872
rect 490012 152040 490064 152046
rect 490012 151982 490064 151988
rect 490024 149954 490052 151982
rect 490656 151972 490708 151978
rect 490656 151914 490708 151920
rect 490668 149954 490696 151914
rect 491944 151904 491996 151910
rect 491944 151846 491996 151852
rect 491300 151836 491352 151842
rect 491300 151778 491352 151784
rect 491312 149954 491340 151778
rect 491956 149954 491984 151846
rect 492784 149954 492812 153070
rect 493244 149954 493272 153138
rect 494072 153134 494100 163200
rect 494164 153202 494192 163254
rect 494900 163146 494928 163254
rect 494978 163200 495034 164400
rect 495544 163254 495756 163282
rect 494992 163146 495020 163200
rect 494900 163118 495020 163146
rect 494152 153196 494204 153202
rect 494152 153138 494204 153144
rect 494060 153128 494112 153134
rect 494060 153070 494112 153076
rect 495544 153066 495572 163254
rect 495728 163146 495756 163254
rect 495806 163200 495862 164400
rect 496634 163200 496690 164400
rect 496832 163254 497412 163282
rect 495820 163146 495848 163200
rect 495728 163118 495848 163146
rect 496648 153202 496676 163200
rect 496452 153196 496504 153202
rect 496452 153138 496504 153144
rect 496636 153196 496688 153202
rect 496636 153138 496688 153144
rect 495808 153128 495860 153134
rect 495808 153070 495860 153076
rect 495440 153060 495492 153066
rect 495440 153002 495492 153008
rect 495532 153060 495584 153066
rect 495532 153002 495584 153008
rect 494060 152992 494112 152998
rect 494060 152934 494112 152940
rect 494072 149954 494100 152934
rect 494520 152924 494572 152930
rect 494520 152866 494572 152872
rect 494532 149954 494560 152866
rect 495452 150226 495480 153002
rect 495452 150198 495526 150226
rect 487540 149926 487876 149954
rect 488092 149926 488520 149954
rect 488736 149926 489072 149954
rect 489380 149926 489716 149954
rect 490024 149926 490360 149954
rect 490668 149926 491004 149954
rect 491312 149926 491648 149954
rect 491956 149926 492292 149954
rect 492784 149926 492936 149954
rect 493244 149926 493580 149954
rect 494072 149926 494224 149954
rect 494532 149926 494868 149954
rect 495498 149940 495526 150198
rect 495820 149954 495848 153070
rect 496464 149954 496492 153138
rect 496832 153134 496860 163254
rect 497384 163146 497412 163254
rect 497462 163200 497518 164400
rect 498290 163200 498346 164400
rect 498396 163254 498976 163282
rect 497476 163146 497504 163200
rect 497384 163118 497504 163146
rect 498304 163146 498332 163200
rect 498396 163146 498424 163254
rect 498304 163118 498424 163146
rect 497740 153196 497792 153202
rect 497740 153138 497792 153144
rect 496820 153128 496872 153134
rect 496820 153070 496872 153076
rect 497096 153060 497148 153066
rect 497096 153002 497148 153008
rect 497108 149954 497136 153002
rect 497752 149954 497780 153138
rect 498384 153128 498436 153134
rect 498384 153070 498436 153076
rect 498396 149954 498424 153070
rect 498948 149954 498976 163254
rect 499118 163200 499174 164400
rect 499946 163200 500002 164400
rect 500052 163254 500264 163282
rect 499132 151842 499160 163200
rect 499960 163146 499988 163200
rect 500052 163146 500080 163254
rect 499960 163118 500080 163146
rect 499120 151836 499172 151842
rect 499120 151778 499172 151784
rect 499764 151836 499816 151842
rect 499764 151778 499816 151784
rect 499776 149954 499804 151778
rect 500236 149954 500264 163254
rect 500866 163200 500922 164400
rect 501694 163200 501750 164400
rect 502522 163200 502578 164400
rect 503350 163200 503406 164400
rect 503732 163254 504128 163282
rect 500880 151814 500908 163200
rect 501708 161474 501736 163200
rect 501524 161446 501736 161474
rect 500880 151786 501000 151814
rect 500972 149954 501000 151786
rect 501524 149954 501552 161446
rect 502536 150226 502564 163200
rect 502536 150198 502610 150226
rect 495820 149926 496156 149954
rect 496464 149926 496800 149954
rect 497108 149926 497444 149954
rect 497752 149926 498088 149954
rect 498396 149926 498732 149954
rect 498948 149926 499376 149954
rect 499776 149926 500020 149954
rect 500236 149926 500664 149954
rect 500972 149926 501308 149954
rect 501524 149926 501952 149954
rect 502582 149940 502610 150198
rect 503364 149954 503392 163200
rect 503240 149926 503392 149954
rect 503732 149954 503760 163254
rect 504100 163146 504128 163254
rect 504178 163200 504234 164400
rect 504284 163254 504956 163282
rect 504192 163146 504220 163200
rect 504100 163118 504220 163146
rect 504284 149954 504312 163254
rect 504928 163146 504956 163254
rect 505006 163200 505062 164400
rect 505112 163254 505784 163282
rect 505020 163146 505048 163200
rect 504928 163118 505048 163146
rect 505112 150226 505140 163254
rect 505756 163146 505784 163254
rect 505834 163200 505890 164400
rect 506754 163200 506810 164400
rect 507582 163200 507638 164400
rect 508410 163200 508466 164400
rect 509238 163200 509294 164400
rect 509344 163254 509556 163282
rect 505848 163146 505876 163200
rect 505756 163118 505876 163146
rect 506664 158976 506716 158982
rect 506664 158918 506716 158924
rect 506112 158840 506164 158846
rect 506112 158782 506164 158788
rect 505376 158772 505428 158778
rect 505376 158714 505428 158720
rect 505112 150198 505186 150226
rect 503732 149926 503884 149954
rect 504284 149926 504528 149954
rect 505158 149940 505186 150198
rect 505388 149954 505416 158714
rect 506124 149954 506152 158782
rect 506676 149954 506704 158918
rect 506768 158778 506796 163200
rect 507596 158846 507624 163200
rect 508424 158982 508452 163200
rect 509252 163146 509280 163200
rect 509344 163146 509372 163254
rect 509252 163118 509372 163146
rect 508412 158976 508464 158982
rect 508412 158918 508464 158924
rect 507952 158908 508004 158914
rect 507952 158850 508004 158856
rect 507584 158840 507636 158846
rect 507584 158782 507636 158788
rect 506756 158772 506808 158778
rect 506756 158714 506808 158720
rect 507768 151904 507820 151910
rect 507768 151846 507820 151852
rect 507780 150226 507808 151846
rect 507734 150198 507808 150226
rect 505388 149926 505816 149954
rect 506124 149926 506460 149954
rect 506676 149926 507104 149954
rect 507734 149940 507762 150198
rect 507964 149954 507992 158850
rect 509332 158772 509384 158778
rect 509332 158714 509384 158720
rect 509148 151972 509200 151978
rect 509148 151914 509200 151920
rect 509160 149954 509188 151914
rect 507964 149926 508392 149954
rect 509036 149926 509188 149954
rect 509344 149954 509372 158714
rect 509528 151910 509556 163254
rect 510066 163200 510122 164400
rect 510894 163200 510950 164400
rect 511722 163200 511778 164400
rect 512012 163254 512592 163282
rect 510080 158914 510108 163200
rect 510068 158908 510120 158914
rect 510068 158850 510120 158856
rect 510528 152788 510580 152794
rect 510528 152730 510580 152736
rect 509516 151904 509568 151910
rect 509516 151846 509568 151852
rect 510540 149954 510568 152730
rect 510908 151978 510936 163200
rect 511736 158778 511764 163200
rect 511724 158772 511776 158778
rect 511724 158714 511776 158720
rect 511264 153128 511316 153134
rect 511264 153070 511316 153076
rect 510896 151972 510948 151978
rect 510896 151914 510948 151920
rect 511276 149954 511304 153070
rect 511724 153060 511776 153066
rect 511724 153002 511776 153008
rect 511736 149954 511764 153002
rect 512012 152794 512040 163254
rect 512564 163146 512592 163254
rect 512642 163200 512698 164400
rect 513470 163200 513526 164400
rect 514298 163200 514354 164400
rect 514864 163254 515076 163282
rect 512656 163146 512684 163200
rect 512564 163118 512684 163146
rect 512552 153196 512604 153202
rect 512552 153138 512604 153144
rect 512000 152788 512052 152794
rect 512000 152730 512052 152736
rect 512564 149954 512592 153138
rect 513484 153134 513512 163200
rect 513472 153128 513524 153134
rect 513472 153070 513524 153076
rect 514312 153066 514340 163200
rect 514864 153202 514892 163254
rect 515048 163146 515076 163254
rect 515126 163200 515182 164400
rect 515954 163200 516010 164400
rect 516152 163254 516732 163282
rect 515140 163146 515168 163200
rect 515048 163118 515168 163146
rect 514944 158772 514996 158778
rect 514944 158714 514996 158720
rect 514852 153196 514904 153202
rect 514852 153138 514904 153144
rect 514484 153128 514536 153134
rect 514484 153070 514536 153076
rect 514300 153060 514352 153066
rect 514300 153002 514352 153008
rect 513196 152992 513248 152998
rect 513196 152934 513248 152940
rect 513208 149954 513236 152934
rect 513840 152924 513892 152930
rect 513840 152866 513892 152872
rect 513852 149954 513880 152866
rect 514496 149954 514524 153070
rect 514956 149954 514984 158714
rect 515968 152998 515996 163200
rect 515956 152992 516008 152998
rect 515956 152934 516008 152940
rect 516152 152930 516180 163254
rect 516704 163146 516732 163254
rect 516782 163200 516838 164400
rect 517610 163200 517666 164400
rect 518530 163200 518586 164400
rect 519004 163254 519308 163282
rect 516796 163146 516824 163200
rect 516704 163118 516824 163146
rect 517624 161474 517652 163200
rect 517532 161446 517652 161474
rect 517532 158794 517560 161446
rect 518348 159452 518400 159458
rect 518348 159394 518400 159400
rect 517612 159384 517664 159390
rect 517612 159326 517664 159332
rect 517440 158766 517560 158794
rect 517440 153134 517468 158766
rect 517428 153128 517480 153134
rect 517428 153070 517480 153076
rect 516140 152924 516192 152930
rect 516140 152866 516192 152872
rect 515772 152108 515824 152114
rect 515772 152050 515824 152056
rect 515784 149954 515812 152050
rect 516048 152040 516100 152046
rect 516048 151982 516100 151988
rect 516060 150226 516088 151982
rect 517428 151972 517480 151978
rect 517428 151914 517480 151920
rect 517060 151836 517112 151842
rect 517060 151778 517112 151784
rect 516060 150198 516134 150226
rect 509344 149926 509680 149954
rect 510324 149926 510568 149954
rect 510968 149926 511304 149954
rect 511612 149926 511764 149954
rect 512256 149926 512592 149954
rect 512900 149926 513236 149954
rect 513544 149926 513880 149954
rect 514188 149926 514524 149954
rect 514832 149926 514984 149954
rect 515476 149926 515812 149954
rect 516106 149940 516134 150198
rect 517072 149954 517100 151778
rect 517440 150226 517468 151914
rect 516764 149926 517100 149954
rect 517394 150198 517468 150226
rect 517394 149940 517422 150198
rect 517624 149954 517652 159326
rect 518360 149954 518388 159394
rect 518544 158778 518572 163200
rect 518532 158772 518584 158778
rect 518532 158714 518584 158720
rect 519004 152114 519032 163254
rect 519280 163146 519308 163254
rect 519358 163200 519414 164400
rect 520186 163200 520242 164400
rect 520292 163254 520964 163282
rect 519372 163146 519400 163200
rect 519280 163118 519400 163146
rect 519726 163160 519782 163169
rect 519726 163095 519782 163104
rect 519542 161664 519598 161673
rect 519542 161599 519598 161608
rect 518992 152108 519044 152114
rect 518992 152050 519044 152056
rect 517624 149926 518052 149954
rect 518360 149926 518696 149954
rect 430316 149790 430652 149818
rect 519556 147937 519584 161599
rect 519634 160168 519690 160177
rect 519634 160103 519690 160112
rect 519542 147928 519598 147937
rect 519542 147863 519598 147872
rect 519648 146577 519676 160103
rect 519740 149297 519768 163095
rect 519818 158672 519874 158681
rect 519818 158607 519874 158616
rect 519726 149288 519782 149297
rect 519726 149223 519782 149232
rect 519726 148064 519782 148073
rect 519726 147999 519782 148008
rect 519634 146568 519690 146577
rect 519634 146503 519690 146512
rect 519450 143440 519506 143449
rect 519450 143375 519506 143384
rect 519358 141944 519414 141953
rect 519358 141879 519414 141888
rect 519266 140448 519322 140457
rect 519266 140383 519322 140392
rect 117240 132518 117360 132546
rect 117332 132410 117360 132518
rect 117240 132382 117360 132410
rect 117240 127945 117268 132382
rect 519280 128897 519308 140383
rect 519372 130257 519400 141879
rect 519464 131617 519492 143375
rect 519740 135697 519768 147999
rect 519832 145217 519860 158607
rect 520002 157176 520058 157185
rect 520002 157111 520058 157120
rect 519910 151056 519966 151065
rect 519910 150991 519966 151000
rect 519818 145208 519874 145217
rect 519818 145143 519874 145152
rect 519924 138417 519952 150991
rect 520016 143857 520044 157111
rect 520094 154048 520150 154057
rect 520094 153983 520150 153992
rect 520002 143848 520058 143857
rect 520002 143783 520058 143792
rect 520108 141137 520136 153983
rect 520200 152046 520228 163200
rect 520188 152040 520240 152046
rect 520188 151982 520240 151988
rect 520292 151842 520320 163254
rect 520936 163146 520964 163254
rect 521014 163200 521070 164400
rect 521842 163200 521898 164400
rect 522670 163200 522726 164400
rect 523498 163200 523554 164400
rect 521028 163146 521056 163200
rect 520936 163118 521056 163146
rect 521856 161474 521884 163200
rect 521672 161446 521884 161474
rect 521672 158794 521700 161446
rect 522684 159390 522712 163200
rect 523512 159458 523540 163200
rect 523500 159452 523552 159458
rect 523500 159394 523552 159400
rect 522672 159384 522724 159390
rect 522672 159326 522724 159332
rect 521580 158766 521700 158794
rect 521106 155680 521162 155689
rect 521106 155615 521162 155624
rect 521014 152552 521070 152561
rect 521014 152487 521070 152496
rect 520280 151836 520332 151842
rect 520280 151778 520332 151784
rect 520186 149560 520242 149569
rect 520186 149495 520242 149504
rect 520094 141128 520150 141137
rect 520094 141063 520150 141072
rect 520094 138952 520150 138961
rect 520094 138887 520150 138896
rect 519910 138408 519966 138417
rect 519910 138343 519966 138352
rect 520002 137456 520058 137465
rect 520002 137391 520058 137400
rect 519910 135824 519966 135833
rect 519910 135759 519966 135768
rect 519726 135688 519782 135697
rect 519726 135623 519782 135632
rect 519818 134328 519874 134337
rect 519818 134263 519874 134272
rect 519542 132832 519598 132841
rect 519542 132767 519598 132776
rect 519450 131608 519506 131617
rect 519450 131543 519506 131552
rect 519358 130248 519414 130257
rect 519358 130183 519414 130192
rect 519266 128888 519322 128897
rect 519266 128823 519322 128832
rect 519450 128344 519506 128353
rect 519450 128279 519506 128288
rect 117226 127936 117282 127945
rect 117226 127871 117282 127880
rect 519358 120592 519414 120601
rect 519358 120527 519414 120536
rect 519372 111217 519400 120527
rect 519464 118017 519492 128279
rect 519556 122097 519584 132767
rect 519726 131336 519782 131345
rect 519726 131271 519782 131280
rect 519634 129840 519690 129849
rect 519634 129775 519690 129784
rect 519542 122088 519598 122097
rect 519542 122023 519598 122032
rect 519648 119377 519676 129775
rect 519740 120737 519768 131271
rect 519832 123457 519860 134263
rect 519924 124817 519952 135759
rect 520016 126177 520044 137391
rect 520108 127537 520136 138887
rect 520200 137057 520228 149495
rect 520922 144936 520978 144945
rect 520922 144871 520978 144880
rect 520186 137048 520242 137057
rect 520186 136983 520242 136992
rect 520936 132977 520964 144871
rect 521028 139777 521056 152487
rect 521120 142497 521148 155615
rect 521580 151978 521608 158766
rect 521568 151972 521620 151978
rect 521568 151914 521620 151920
rect 521198 146568 521254 146577
rect 521198 146503 521254 146512
rect 521106 142488 521162 142497
rect 521106 142423 521162 142432
rect 521014 139768 521070 139777
rect 521014 139703 521070 139712
rect 521212 134473 521240 146503
rect 521198 134464 521254 134473
rect 521198 134399 521254 134408
rect 520922 132968 520978 132977
rect 520922 132903 520978 132912
rect 520094 127528 520150 127537
rect 520094 127463 520150 127472
rect 520186 126712 520242 126721
rect 520186 126647 520242 126656
rect 520002 126168 520058 126177
rect 520002 126103 520058 126112
rect 520094 125216 520150 125225
rect 520094 125151 520150 125160
rect 519910 124808 519966 124817
rect 519910 124743 519966 124752
rect 520002 123720 520058 123729
rect 520002 123655 520058 123664
rect 519818 123448 519874 123457
rect 519818 123383 519874 123392
rect 519910 122224 519966 122233
rect 519910 122159 519966 122168
rect 519726 120728 519782 120737
rect 519726 120663 519782 120672
rect 519634 119368 519690 119377
rect 519634 119303 519690 119312
rect 519818 119232 519874 119241
rect 519818 119167 519874 119176
rect 519450 118008 519506 118017
rect 519450 117943 519506 117952
rect 519726 117600 519782 117609
rect 519726 117535 519782 117544
rect 519542 116104 519598 116113
rect 519542 116039 519598 116048
rect 519358 111208 519414 111217
rect 519358 111143 519414 111152
rect 519556 107137 519584 116039
rect 519634 114608 519690 114617
rect 519634 114543 519690 114552
rect 519542 107128 519598 107137
rect 519542 107063 519598 107072
rect 519648 105777 519676 114543
rect 519740 108497 519768 117535
rect 519832 109857 519860 119167
rect 519924 112577 519952 122159
rect 520016 113937 520044 123655
rect 520108 115297 520136 125151
rect 520200 116657 520228 126647
rect 520186 116648 520242 116657
rect 520186 116583 520242 116592
rect 520094 115288 520150 115297
rect 520094 115223 520150 115232
rect 520002 113928 520058 113937
rect 520002 113863 520058 113872
rect 521106 113112 521162 113121
rect 521106 113047 521162 113056
rect 519910 112568 519966 112577
rect 519910 112503 519966 112512
rect 519818 109848 519874 109857
rect 519818 109783 519874 109792
rect 519726 108488 519782 108497
rect 519726 108423 519782 108432
rect 521014 108488 521070 108497
rect 521014 108423 521070 108432
rect 520922 106992 520978 107001
rect 520922 106927 520978 106936
rect 519634 105768 519690 105777
rect 519634 105703 519690 105712
rect 520278 105496 520334 105505
rect 520278 105431 520334 105440
rect 117134 104816 117190 104825
rect 117134 104751 117190 104760
rect 117042 101008 117098 101017
rect 117042 100943 117098 100952
rect 519818 99376 519874 99385
rect 519818 99311 519874 99320
rect 116858 99104 116914 99113
rect 116858 99039 116914 99048
rect 519726 97880 519782 97889
rect 519726 97815 519782 97824
rect 116766 97200 116822 97209
rect 116766 97135 116822 97144
rect 519266 96384 519322 96393
rect 519266 96319 519322 96328
rect 116674 95296 116730 95305
rect 116674 95231 116730 95240
rect 116582 93392 116638 93401
rect 116582 93327 116638 93336
rect 116124 92472 116176 92478
rect 116124 92414 116176 92420
rect 116136 91361 116164 92414
rect 116122 91352 116178 91361
rect 116122 91287 116178 91296
rect 116124 89684 116176 89690
rect 116124 89626 116176 89632
rect 116136 89457 116164 89626
rect 519280 89457 519308 96319
rect 519740 90817 519768 97815
rect 519832 92177 519860 99311
rect 520292 97617 520320 105431
rect 520936 98977 520964 106927
rect 521028 100337 521056 108423
rect 521120 104417 521148 113047
rect 521566 111616 521622 111625
rect 521566 111551 521622 111560
rect 521290 110120 521346 110129
rect 521290 110055 521346 110064
rect 521106 104408 521162 104417
rect 521106 104343 521162 104352
rect 521198 104000 521254 104009
rect 521198 103935 521254 103944
rect 521106 102504 521162 102513
rect 521106 102439 521162 102448
rect 521014 100328 521070 100337
rect 521014 100263 521070 100272
rect 520922 98968 520978 98977
rect 520922 98903 520978 98912
rect 520278 97608 520334 97617
rect 520278 97543 520334 97552
rect 521120 95033 521148 102439
rect 521212 96257 521240 103935
rect 521304 101697 521332 110055
rect 521580 103057 521608 111551
rect 521566 103048 521622 103057
rect 521566 102983 521622 102992
rect 521290 101688 521346 101697
rect 521290 101623 521346 101632
rect 521474 101008 521530 101017
rect 521474 100943 521530 100952
rect 521198 96248 521254 96257
rect 521198 96183 521254 96192
rect 521106 95024 521162 95033
rect 521106 94959 521162 94968
rect 519910 94888 519966 94897
rect 519910 94823 519966 94832
rect 519818 92168 519874 92177
rect 519818 92103 519874 92112
rect 519726 90808 519782 90817
rect 519726 90743 519782 90752
rect 116122 89448 116178 89457
rect 116122 89383 116178 89392
rect 519266 89448 519322 89457
rect 519266 89383 519322 89392
rect 116032 88324 116084 88330
rect 116032 88266 116084 88272
rect 116044 87553 116072 88266
rect 519924 88097 519952 94823
rect 521488 93537 521516 100943
rect 521474 93528 521530 93537
rect 521474 93463 521530 93472
rect 520186 93392 520242 93401
rect 520186 93327 520242 93336
rect 519910 88088 519966 88097
rect 519910 88023 519966 88032
rect 116030 87544 116086 87553
rect 116030 87479 116086 87488
rect 520200 86737 520228 93327
rect 521290 91896 521346 91905
rect 521290 91831 521346 91840
rect 520922 90264 520978 90273
rect 520922 90199 520978 90208
rect 520186 86728 520242 86737
rect 520186 86663 520242 86672
rect 520278 85776 520334 85785
rect 520278 85711 520334 85720
rect 115202 85640 115258 85649
rect 115202 85575 115258 85584
rect 116584 83972 116636 83978
rect 116584 83914 116636 83920
rect 116596 83745 116624 83914
rect 116582 83736 116638 83745
rect 116582 83671 116638 83680
rect 116216 82816 116268 82822
rect 116216 82758 116268 82764
rect 520186 82784 520242 82793
rect 116228 81841 116256 82758
rect 520186 82719 520242 82728
rect 116214 81832 116270 81841
rect 116214 81767 116270 81776
rect 519634 81152 519690 81161
rect 519634 81087 519690 81096
rect 115940 80028 115992 80034
rect 115940 79970 115992 79976
rect 115952 79937 115980 79970
rect 115938 79928 115994 79937
rect 115938 79863 115994 79872
rect 114192 78668 114244 78674
rect 114192 78610 114244 78616
rect 116124 78668 116176 78674
rect 116124 78610 116176 78616
rect 116136 78033 116164 78610
rect 116122 78024 116178 78033
rect 116122 77959 116178 77968
rect 519648 74633 519676 81087
rect 519818 79656 519874 79665
rect 519818 79591 519874 79600
rect 519726 76664 519782 76673
rect 519726 76599 519782 76608
rect 519634 74624 519690 74633
rect 519634 74559 519690 74568
rect 116674 74080 116730 74089
rect 116674 74015 116730 74024
rect 116582 72176 116638 72185
rect 116582 72111 116638 72120
rect 116596 71806 116624 72111
rect 114192 71800 114244 71806
rect 114192 71742 114244 71748
rect 116584 71800 116636 71806
rect 116584 71742 116636 71748
rect 114100 69080 114152 69086
rect 114100 69022 114152 69028
rect 114008 67652 114060 67658
rect 114008 67594 114060 67600
rect 113916 66292 113968 66298
rect 113916 66234 113968 66240
rect 113364 64728 113416 64734
rect 113364 64670 113416 64676
rect 113376 64569 113404 64670
rect 113362 64560 113418 64569
rect 113362 64495 113418 64504
rect 113824 63572 113876 63578
rect 113824 63514 113876 63520
rect 112444 62144 112496 62150
rect 112444 62086 112496 62092
rect 110326 58032 110382 58041
rect 109696 57990 110326 58018
rect 109696 45554 109724 57990
rect 110326 57967 110382 57976
rect 110326 56808 110382 56817
rect 110326 56743 110382 56752
rect 110340 55214 110368 56743
rect 109512 45526 109724 45554
rect 109788 55186 110368 55214
rect 109512 39522 109540 45526
rect 109788 39658 109816 55186
rect 110326 53952 110382 53961
rect 109880 53910 110326 53938
rect 109880 41562 109908 53910
rect 110326 53887 110382 53896
rect 110326 52592 110382 52601
rect 110326 52527 110382 52536
rect 110340 51218 110368 52527
rect 110340 51190 110460 51218
rect 110326 51096 110382 51105
rect 109972 51054 110326 51082
rect 109972 42378 110000 51054
rect 110326 51031 110382 51040
rect 110432 50946 110460 51190
rect 110064 50918 110460 50946
rect 110064 44690 110092 50918
rect 110326 48376 110382 48385
rect 110156 48334 110326 48362
rect 110156 45554 110184 48334
rect 110326 48311 110382 48320
rect 110326 47152 110382 47161
rect 110326 47087 110382 47096
rect 110156 45526 110276 45554
rect 110248 44962 110276 45526
rect 110340 45121 110368 47087
rect 110326 45112 110382 45121
rect 110326 45047 110382 45056
rect 110878 45112 110934 45121
rect 110878 45047 110934 45056
rect 110326 44976 110382 44985
rect 110248 44934 110326 44962
rect 110326 44911 110382 44920
rect 110064 44662 110460 44690
rect 110432 44174 110460 44662
rect 110432 44146 110736 44174
rect 109972 42350 110644 42378
rect 109880 41534 110552 41562
rect 110418 41440 110474 41449
rect 110418 41375 110474 41384
rect 109788 39630 110368 39658
rect 109512 39494 110092 39522
rect 110064 38654 110092 39494
rect 110064 38626 110276 38654
rect 110248 35306 110276 38626
rect 110340 37369 110368 39630
rect 110326 37360 110382 37369
rect 110326 37295 110382 37304
rect 110326 35320 110382 35329
rect 110248 35278 110326 35306
rect 110326 35255 110382 35264
rect 110326 35184 110382 35193
rect 109512 35142 110326 35170
rect 109512 3641 109540 35142
rect 110326 35119 110382 35128
rect 110432 34898 110460 41375
rect 109604 34870 110460 34898
rect 109604 29866 109632 34870
rect 110326 33824 110382 33833
rect 109972 33782 110326 33810
rect 109604 29838 109724 29866
rect 109696 29594 109724 29838
rect 109604 29566 109724 29594
rect 109498 3632 109554 3641
rect 109498 3567 109554 3576
rect 109406 3496 109462 3505
rect 109406 3431 109462 3440
rect 109420 2961 109448 3431
rect 109498 3360 109554 3369
rect 109498 3295 109554 3304
rect 109406 2952 109462 2961
rect 109406 2887 109462 2896
rect 33046 2680 33102 2689
rect 33046 2615 33102 2624
rect 42062 2680 42118 2689
rect 42706 2680 42762 2689
rect 42642 2638 42706 2666
rect 42062 2615 42118 2624
rect 42706 2615 42762 2624
rect 44730 2680 44786 2689
rect 44730 2615 44786 2624
rect 62394 2680 62450 2689
rect 63038 2680 63094 2689
rect 62698 2638 63038 2666
rect 62394 2615 62450 2624
rect 63038 2615 63094 2624
rect 64050 2680 64106 2689
rect 64050 2615 64106 2624
rect 68282 2680 68338 2689
rect 68282 2615 68338 2624
rect 78770 2680 78826 2689
rect 78770 2615 78826 2624
rect 87050 2680 87106 2689
rect 87050 2615 87106 2624
rect 90086 2680 90142 2689
rect 90086 2615 90142 2624
rect 90362 2680 90418 2689
rect 90362 2615 90418 2624
rect 91558 2680 91614 2689
rect 91558 2615 91614 2624
rect 91926 2680 91982 2689
rect 93030 2680 93086 2689
rect 92690 2638 93030 2666
rect 91926 2615 91982 2624
rect 93030 2615 93086 2624
rect 93858 2680 93914 2689
rect 93858 2615 93914 2624
rect 95698 2680 95754 2689
rect 95698 2615 95754 2624
rect 97722 2680 97778 2689
rect 97722 2615 97778 2624
rect 97906 2680 97962 2689
rect 97906 2615 97962 2624
rect 99194 2680 99250 2689
rect 99194 2615 99250 2624
rect 103702 2680 103758 2689
rect 103702 2615 103758 2624
rect 104438 2680 104494 2689
rect 104990 2680 105046 2689
rect 104494 2638 104990 2666
rect 104438 2615 104494 2624
rect 104990 2615 105046 2624
rect 106186 2680 106242 2689
rect 106370 2680 106426 2689
rect 106242 2638 106370 2666
rect 106186 2615 106242 2624
rect 106370 2615 106426 2624
rect 29550 2544 29606 2553
rect 29302 2502 29550 2530
rect 29550 2479 29606 2488
rect 26054 2408 26110 2417
rect 25990 2366 26054 2394
rect 26054 2343 26110 2352
rect 22926 2272 22982 2281
rect 22678 2230 22926 2258
rect 22926 2207 22982 2216
rect 19614 2136 19670 2145
rect 2700 1358 2728 2108
rect 6012 1873 6040 2108
rect 5998 1864 6054 1873
rect 5998 1799 6054 1808
rect 9324 1601 9352 2108
rect 12636 1737 12664 2108
rect 15962 2094 16252 2122
rect 19366 2094 19614 2122
rect 16224 2009 16252 2094
rect 19614 2071 19670 2080
rect 16210 2000 16266 2009
rect 16210 1935 16266 1944
rect 12622 1728 12678 1737
rect 12622 1663 12678 1672
rect 9310 1592 9366 1601
rect 9310 1527 9366 1536
rect 32692 1426 32720 2108
rect 32680 1420 32732 1426
rect 32680 1362 32732 1368
rect 2688 1352 2740 1358
rect 2688 1294 2740 1300
rect 32784 870 32904 898
rect 32784 800 32812 870
rect 32770 -400 32826 800
rect 32876 762 32904 870
rect 33060 762 33088 2615
rect 36004 1290 36032 2108
rect 35992 1284 36044 1290
rect 35992 1226 36044 1232
rect 39316 1222 39344 2108
rect 42076 1902 42104 2615
rect 44744 1902 44772 2615
rect 42064 1896 42116 1902
rect 42064 1838 42116 1844
rect 44732 1896 44784 1902
rect 44732 1838 44784 1844
rect 46032 1494 46060 2108
rect 46020 1488 46072 1494
rect 46020 1430 46072 1436
rect 39304 1216 39356 1222
rect 39304 1158 39356 1164
rect 49344 1154 49372 2108
rect 49332 1148 49384 1154
rect 49332 1090 49384 1096
rect 52656 1086 52684 2108
rect 55968 1465 55996 2108
rect 59372 1766 59400 2108
rect 62408 1902 62436 2615
rect 62396 1896 62448 1902
rect 62396 1838 62448 1844
rect 59360 1760 59412 1766
rect 59360 1702 59412 1708
rect 64064 1494 64092 2615
rect 64052 1488 64104 1494
rect 55954 1456 56010 1465
rect 64052 1430 64104 1436
rect 55954 1391 56010 1400
rect 52644 1080 52696 1086
rect 52644 1022 52696 1028
rect 65996 1018 66024 2108
rect 68296 1902 68324 2615
rect 68284 1896 68336 1902
rect 68284 1838 68336 1844
rect 69308 1630 69336 2108
rect 69296 1624 69348 1630
rect 69296 1566 69348 1572
rect 72712 1494 72740 2108
rect 72700 1488 72752 1494
rect 72700 1430 72752 1436
rect 65984 1012 66036 1018
rect 65984 954 66036 960
rect 76024 950 76052 2108
rect 78784 1766 78812 2615
rect 78772 1760 78824 1766
rect 78772 1702 78824 1708
rect 79336 1562 79364 2108
rect 82648 1698 82676 2108
rect 86052 1766 86080 2108
rect 86040 1760 86092 1766
rect 86040 1702 86092 1708
rect 82636 1692 82688 1698
rect 82636 1634 82688 1640
rect 79324 1556 79376 1562
rect 79324 1498 79376 1504
rect 87064 1329 87092 2615
rect 89364 1834 89392 2108
rect 89352 1828 89404 1834
rect 89352 1770 89404 1776
rect 87050 1320 87106 1329
rect 87050 1255 87106 1264
rect 90100 1057 90128 2615
rect 90376 1193 90404 2615
rect 90362 1184 90418 1193
rect 90362 1119 90418 1128
rect 90086 1048 90142 1057
rect 90086 983 90142 992
rect 76012 944 76064 950
rect 76012 886 76064 892
rect 91572 882 91600 2615
rect 91940 1902 91968 2615
rect 91928 1896 91980 1902
rect 91928 1838 91980 1844
rect 93872 882 93900 2615
rect 95712 1329 95740 2615
rect 95988 1329 96016 2108
rect 95698 1320 95754 1329
rect 95698 1255 95754 1264
rect 95974 1320 96030 1329
rect 95974 1255 96030 1264
rect 97736 1193 97764 2615
rect 97920 1329 97948 2615
rect 99208 1902 99236 2615
rect 99196 1896 99248 1902
rect 99196 1838 99248 1844
rect 97906 1320 97962 1329
rect 97906 1255 97962 1264
rect 98274 1320 98330 1329
rect 98274 1255 98330 1264
rect 97722 1184 97778 1193
rect 97722 1119 97778 1128
rect 97264 1012 97316 1018
rect 97264 954 97316 960
rect 97276 882 97304 954
rect 91560 876 91612 882
rect 91560 818 91612 824
rect 93860 876 93912 882
rect 93860 818 93912 824
rect 97264 876 97316 882
rect 97264 818 97316 824
rect 98288 800 98316 1255
rect 99392 1193 99420 2108
rect 102704 1902 102732 2108
rect 102600 1896 102652 1902
rect 102600 1838 102652 1844
rect 102692 1896 102744 1902
rect 102692 1838 102744 1844
rect 102612 1193 102640 1838
rect 103716 1193 103744 2615
rect 104438 2408 104494 2417
rect 104622 2408 104678 2417
rect 104494 2366 104622 2394
rect 104438 2343 104494 2352
rect 104622 2343 104678 2352
rect 104438 2272 104494 2281
rect 104622 2272 104678 2281
rect 104494 2230 104622 2258
rect 104438 2207 104494 2216
rect 104622 2207 104678 2216
rect 104346 2136 104402 2145
rect 104622 2136 104678 2145
rect 104402 2094 104622 2122
rect 104346 2071 104402 2080
rect 104622 2071 104678 2080
rect 105912 1896 105964 1902
rect 105912 1838 105964 1844
rect 103980 1692 104032 1698
rect 103980 1634 104032 1640
rect 103796 1624 103848 1630
rect 103796 1566 103848 1572
rect 99378 1184 99434 1193
rect 99378 1119 99434 1128
rect 102598 1184 102654 1193
rect 102598 1119 102654 1128
rect 103702 1184 103758 1193
rect 103702 1119 103758 1128
rect 32876 734 33088 762
rect 98274 -400 98330 800
rect 103808 746 103836 1566
rect 103992 1562 104020 1634
rect 105924 1630 105952 1838
rect 106016 1630 106044 2108
rect 109132 1896 109184 1902
rect 109184 1844 109264 1850
rect 109132 1838 109264 1844
rect 109144 1822 109264 1838
rect 109328 1834 109356 2108
rect 109236 1698 109264 1822
rect 109316 1828 109368 1834
rect 109316 1770 109368 1776
rect 109224 1692 109276 1698
rect 109224 1634 109276 1640
rect 105912 1624 105964 1630
rect 105912 1566 105964 1572
rect 106004 1624 106056 1630
rect 106004 1566 106056 1572
rect 109040 1624 109092 1630
rect 109092 1572 109264 1578
rect 109040 1566 109264 1572
rect 103980 1556 104032 1562
rect 109052 1550 109264 1566
rect 103980 1498 104032 1504
rect 109236 1426 109264 1550
rect 109132 1420 109184 1426
rect 109132 1362 109184 1368
rect 109224 1420 109276 1426
rect 109224 1362 109276 1368
rect 109144 1306 109172 1362
rect 109408 1352 109460 1358
rect 109144 1300 109408 1306
rect 109144 1294 109460 1300
rect 109144 1278 109448 1294
rect 109040 1216 109092 1222
rect 109512 1193 109540 3295
rect 109604 1494 109632 29566
rect 109972 28994 110000 33782
rect 110326 33759 110382 33768
rect 110418 29744 110474 29753
rect 110418 29679 110474 29688
rect 110432 29458 110460 29679
rect 109696 28966 110000 28994
rect 110064 29430 110460 29458
rect 109696 1902 109724 28966
rect 110064 28914 110092 29430
rect 110524 29322 110552 41534
rect 110616 29889 110644 42350
rect 110602 29880 110658 29889
rect 110602 29815 110658 29824
rect 110708 29594 110736 44146
rect 110786 37360 110842 37369
rect 110786 37295 110842 37304
rect 110800 29753 110828 37295
rect 110786 29744 110842 29753
rect 110786 29679 110842 29688
rect 110248 29294 110552 29322
rect 110616 29566 110736 29594
rect 110248 29186 110276 29294
rect 109788 28886 110092 28914
rect 110156 29158 110276 29186
rect 109788 1902 109816 28886
rect 110156 28778 110184 29158
rect 109880 28750 110184 28778
rect 110510 28792 110566 28801
rect 109880 2689 109908 28750
rect 110510 28727 110566 28736
rect 110326 28656 110382 28665
rect 110064 28614 110326 28642
rect 110064 28370 110092 28614
rect 110326 28591 110382 28600
rect 109972 28342 110092 28370
rect 109866 2680 109922 2689
rect 109866 2615 109922 2624
rect 109684 1896 109736 1902
rect 109684 1838 109736 1844
rect 109776 1896 109828 1902
rect 109776 1838 109828 1844
rect 109868 1896 109920 1902
rect 109868 1838 109920 1844
rect 109592 1488 109644 1494
rect 109592 1430 109644 1436
rect 109880 1329 109908 1838
rect 109972 1766 110000 28342
rect 110326 28112 110382 28121
rect 110326 28047 110382 28056
rect 110340 27826 110368 28047
rect 110064 27798 110368 27826
rect 110064 3913 110092 27798
rect 110326 27704 110382 27713
rect 110326 27639 110382 27648
rect 110340 27418 110368 27639
rect 110156 27390 110368 27418
rect 110050 3904 110106 3913
rect 110050 3839 110106 3848
rect 110050 3768 110106 3777
rect 110050 3703 110106 3712
rect 110064 3097 110092 3703
rect 110050 3088 110106 3097
rect 110050 3023 110106 3032
rect 109960 1760 110012 1766
rect 109960 1702 110012 1708
rect 110052 1760 110104 1766
rect 110052 1702 110104 1708
rect 110064 1426 110092 1702
rect 110156 1630 110184 27390
rect 110326 27160 110382 27169
rect 110248 27118 110326 27146
rect 110144 1624 110196 1630
rect 110144 1566 110196 1572
rect 110248 1562 110276 27118
rect 110326 27095 110382 27104
rect 110524 25922 110552 28727
rect 110616 28121 110644 29566
rect 110602 28112 110658 28121
rect 110602 28047 110658 28056
rect 110892 27169 110920 45047
rect 110970 44976 111026 44985
rect 110970 44911 111026 44920
rect 110984 27713 111012 44911
rect 111798 44296 111854 44305
rect 111798 44231 111854 44240
rect 111062 35320 111118 35329
rect 111062 35255 111118 35264
rect 111076 33833 111104 35255
rect 111062 33824 111118 33833
rect 111062 33759 111118 33768
rect 111062 29880 111118 29889
rect 111062 29815 111118 29824
rect 111076 28665 111104 29815
rect 111812 28801 111840 44231
rect 111798 28792 111854 28801
rect 111798 28727 111854 28736
rect 111062 28656 111118 28665
rect 111062 28591 111118 28600
rect 110970 27704 111026 27713
rect 110970 27639 111026 27648
rect 110878 27160 110934 27169
rect 110878 27095 110934 27104
rect 110340 25894 110552 25922
rect 110340 3074 110368 25894
rect 110694 4176 110750 4185
rect 110694 4111 110750 4120
rect 110340 3046 110644 3074
rect 110326 2952 110382 2961
rect 110326 2887 110382 2896
rect 110340 1873 110368 2887
rect 110326 1864 110382 1873
rect 110326 1799 110382 1808
rect 110616 1698 110644 3046
rect 110708 2961 110736 4111
rect 110786 3224 110842 3233
rect 110786 3159 110842 3168
rect 110694 2952 110750 2961
rect 110694 2887 110750 2896
rect 110604 1692 110656 1698
rect 110604 1634 110656 1640
rect 110236 1556 110288 1562
rect 110236 1498 110288 1504
rect 110052 1420 110104 1426
rect 110052 1362 110104 1368
rect 109866 1320 109922 1329
rect 109866 1255 109922 1264
rect 109040 1158 109092 1164
rect 109498 1184 109554 1193
rect 109052 814 109080 1158
rect 109498 1119 109554 1128
rect 109040 808 109092 814
rect 109040 750 109092 756
rect 110800 746 110828 3159
rect 111064 2848 111116 2854
rect 111064 2790 111116 2796
rect 111076 1057 111104 2790
rect 112456 1834 112484 62086
rect 112536 42832 112588 42838
rect 112536 42774 112588 42780
rect 112444 1828 112496 1834
rect 112444 1770 112496 1776
rect 111062 1048 111118 1057
rect 111062 983 111118 992
rect 112548 950 112576 42774
rect 113836 7721 113864 63514
rect 113928 19009 113956 66234
rect 114020 30433 114048 67594
rect 114112 41857 114140 69022
rect 114204 53145 114232 71742
rect 116306 70272 116362 70281
rect 116306 70207 116362 70216
rect 116320 69086 116348 70207
rect 116308 69080 116360 69086
rect 116308 69022 116360 69028
rect 116122 68368 116178 68377
rect 116122 68303 116178 68312
rect 116136 67658 116164 68303
rect 116124 67652 116176 67658
rect 116124 67594 116176 67600
rect 116582 66464 116638 66473
rect 116582 66399 116638 66408
rect 116596 66298 116624 66399
rect 116584 66292 116636 66298
rect 116584 66234 116636 66240
rect 116688 64874 116716 74015
rect 519634 73672 519690 73681
rect 519634 73607 519690 73616
rect 519542 69048 519598 69057
rect 519542 68983 519598 68992
rect 116596 64846 116716 64874
rect 116596 64734 116624 64846
rect 116584 64728 116636 64734
rect 116584 64670 116636 64676
rect 116214 64560 116270 64569
rect 116214 64495 116270 64504
rect 116228 63578 116256 64495
rect 519556 63753 519584 68983
rect 519648 67833 519676 73607
rect 519740 70553 519768 76599
rect 519832 73273 519860 79591
rect 520002 78160 520058 78169
rect 520002 78095 520058 78104
rect 519818 73264 519874 73273
rect 519818 73199 519874 73208
rect 520016 72457 520044 78095
rect 520200 75993 520228 82719
rect 520292 78577 520320 85711
rect 520936 82657 520964 90199
rect 521198 87272 521254 87281
rect 521198 87207 521254 87216
rect 521106 84280 521162 84289
rect 521106 84215 521162 84224
rect 520922 82648 520978 82657
rect 520922 82583 520978 82592
rect 520278 78568 520334 78577
rect 520278 78503 520334 78512
rect 521120 77217 521148 84215
rect 521212 79937 521240 87207
rect 521304 84017 521332 91831
rect 521382 88768 521438 88777
rect 521382 88703 521438 88712
rect 521290 84008 521346 84017
rect 521290 83943 521346 83952
rect 521396 81297 521424 88703
rect 521382 81288 521438 81297
rect 521382 81223 521438 81232
rect 521198 79928 521254 79937
rect 521198 79863 521254 79872
rect 521106 77208 521162 77217
rect 521106 77143 521162 77152
rect 520186 75984 520242 75993
rect 520186 75919 520242 75928
rect 520094 75168 520150 75177
rect 520094 75103 520150 75112
rect 520002 72448 520058 72457
rect 520002 72383 520058 72392
rect 519726 70544 519782 70553
rect 519726 70479 519782 70488
rect 519910 70544 519966 70553
rect 519910 70479 519966 70488
rect 519634 67824 519690 67833
rect 519634 67759 519690 67768
rect 519818 66056 519874 66065
rect 519818 65991 519874 66000
rect 519542 63744 519598 63753
rect 519542 63679 519598 63688
rect 116216 63572 116268 63578
rect 116216 63514 116268 63520
rect 116122 62656 116178 62665
rect 116122 62591 116178 62600
rect 116136 62150 116164 62591
rect 116124 62144 116176 62150
rect 116124 62086 116176 62092
rect 116582 60616 116638 60625
rect 116582 60551 116638 60560
rect 114190 53136 114246 53145
rect 114190 53071 114246 53080
rect 116122 43344 116178 43353
rect 116122 43279 116178 43288
rect 116136 42838 116164 43279
rect 116124 42832 116176 42838
rect 116124 42774 116176 42780
rect 114098 41848 114154 41857
rect 114098 41783 114154 41792
rect 114006 30424 114062 30433
rect 114006 30359 114062 30368
rect 116398 26072 116454 26081
rect 116398 26007 116454 26016
rect 116306 20360 116362 20369
rect 116306 20295 116362 20304
rect 113914 19000 113970 19009
rect 113914 18935 113970 18944
rect 116214 18456 116270 18465
rect 116214 18391 116270 18400
rect 116030 16416 116086 16425
rect 116030 16351 116086 16360
rect 115938 12608 115994 12617
rect 115938 12543 115994 12552
rect 113822 7712 113878 7721
rect 113822 7647 113878 7656
rect 115952 2145 115980 12543
rect 116044 2417 116072 16351
rect 116122 14512 116178 14521
rect 116122 14447 116178 14456
rect 116030 2408 116086 2417
rect 116030 2343 116086 2352
rect 116136 2281 116164 14447
rect 116228 2553 116256 18391
rect 116320 7562 116348 20295
rect 116412 7682 116440 26007
rect 116490 22264 116546 22273
rect 116490 22199 116546 22208
rect 116400 7676 116452 7682
rect 116400 7618 116452 7624
rect 116320 7534 116440 7562
rect 116308 7472 116360 7478
rect 116308 7414 116360 7420
rect 116320 3369 116348 7414
rect 116306 3360 116362 3369
rect 116306 3295 116362 3304
rect 116306 3088 116362 3097
rect 116306 3023 116362 3032
rect 116214 2544 116270 2553
rect 116214 2479 116270 2488
rect 116122 2272 116178 2281
rect 116122 2207 116178 2216
rect 115938 2136 115994 2145
rect 115938 2071 115994 2080
rect 116320 1290 116348 3023
rect 116412 1426 116440 7534
rect 116400 1420 116452 1426
rect 116400 1362 116452 1368
rect 116308 1284 116360 1290
rect 116308 1226 116360 1232
rect 116504 1222 116532 22199
rect 116596 1766 116624 60551
rect 519832 59673 519860 65991
rect 519924 65113 519952 70479
rect 520108 69193 520136 75103
rect 520186 72040 520242 72049
rect 520186 71975 520242 71984
rect 520094 69184 520150 69193
rect 520094 69119 520150 69128
rect 520002 67552 520058 67561
rect 520002 67487 520058 67496
rect 519910 65104 519966 65113
rect 519910 65039 519966 65048
rect 520016 61033 520044 67487
rect 520200 66473 520228 71975
rect 520186 66464 520242 66473
rect 520186 66399 520242 66408
rect 521106 64560 521162 64569
rect 521106 64495 521162 64504
rect 520738 62928 520794 62937
rect 520738 62863 520794 62872
rect 520278 61432 520334 61441
rect 520278 61367 520334 61376
rect 520002 61024 520058 61033
rect 520002 60959 520058 60968
rect 519818 59664 519874 59673
rect 519818 59599 519874 59608
rect 520186 56944 520242 56953
rect 520292 56930 520320 61367
rect 520752 58313 520780 62863
rect 521120 62393 521148 64495
rect 521106 62384 521162 62393
rect 521106 62319 521162 62328
rect 521014 59936 521070 59945
rect 521014 59871 521070 59880
rect 520738 58304 520794 58313
rect 520738 58239 520794 58248
rect 520242 56902 520320 56930
rect 520370 56944 520426 56953
rect 520186 56879 520242 56888
rect 520370 56879 520426 56888
rect 520278 55448 520334 55457
rect 520278 55383 520334 55392
rect 519266 53816 519322 53825
rect 519266 53751 519322 53760
rect 519280 50153 519308 53751
rect 520094 52320 520150 52329
rect 520094 52255 520150 52264
rect 520002 50824 520058 50833
rect 520002 50759 520058 50768
rect 519266 50144 519322 50153
rect 519266 50079 519322 50088
rect 519450 47832 519506 47841
rect 519450 47767 519506 47776
rect 519464 44713 519492 47767
rect 520016 47433 520044 50759
rect 520108 48793 520136 52255
rect 520292 51513 520320 55383
rect 520384 52873 520412 56879
rect 521028 55593 521056 59871
rect 521106 58440 521162 58449
rect 521106 58375 521162 58384
rect 521014 55584 521070 55593
rect 521014 55519 521070 55528
rect 521120 54233 521148 58375
rect 521106 54224 521162 54233
rect 521106 54159 521162 54168
rect 520370 52864 520426 52873
rect 520370 52799 520426 52808
rect 520278 51504 520334 51513
rect 520278 51439 520334 51448
rect 520186 49328 520242 49337
rect 520186 49263 520242 49272
rect 520094 48784 520150 48793
rect 520094 48719 520150 48728
rect 520002 47424 520058 47433
rect 520002 47359 520058 47368
rect 519910 46336 519966 46345
rect 519910 46271 519966 46280
rect 519450 44704 519506 44713
rect 519450 44639 519506 44648
rect 519818 44704 519874 44713
rect 519818 44639 519874 44648
rect 519832 41993 519860 44639
rect 519924 43353 519952 46271
rect 520200 46073 520228 49263
rect 520186 46064 520242 46073
rect 520186 45999 520242 46008
rect 519910 43344 519966 43353
rect 519910 43279 519966 43288
rect 520186 43208 520242 43217
rect 520186 43143 520242 43152
rect 519818 41984 519874 41993
rect 519818 41919 519874 41928
rect 520094 41712 520150 41721
rect 520094 41647 520150 41656
rect 116766 39536 116822 39545
rect 116766 39471 116822 39480
rect 116674 37632 116730 37641
rect 116674 37567 116730 37576
rect 116584 1760 116636 1766
rect 116584 1702 116636 1708
rect 116492 1216 116544 1222
rect 116492 1158 116544 1164
rect 112536 944 112588 950
rect 112536 886 112588 892
rect 116688 882 116716 37567
rect 116780 3233 116808 39471
rect 520108 39273 520136 41647
rect 520200 40633 520228 43143
rect 520186 40624 520242 40633
rect 520186 40559 520242 40568
rect 520186 40216 520242 40225
rect 520186 40151 520242 40160
rect 520094 39264 520150 39273
rect 520094 39199 520150 39208
rect 519818 38720 519874 38729
rect 519818 38655 519874 38664
rect 519832 36553 519860 38655
rect 520200 37913 520228 40151
rect 520186 37904 520242 37913
rect 520186 37839 520242 37848
rect 521566 37224 521622 37233
rect 521566 37159 521622 37168
rect 519818 36544 519874 36553
rect 519818 36479 519874 36488
rect 521580 36009 521608 37159
rect 521566 36000 521622 36009
rect 521566 35935 521622 35944
rect 521106 35592 521162 35601
rect 521106 35527 521162 35536
rect 521120 34513 521148 35527
rect 521106 34504 521162 34513
rect 521106 34439 521162 34448
rect 520922 34096 520978 34105
rect 520922 34031 520978 34040
rect 116950 33824 117006 33833
rect 116950 33759 117006 33768
rect 116858 31784 116914 31793
rect 116858 31719 116914 31728
rect 116766 3224 116822 3233
rect 116766 3159 116822 3168
rect 116872 1018 116900 31719
rect 116964 3777 116992 33759
rect 520936 33153 520964 34031
rect 520922 33144 520978 33153
rect 520922 33079 520978 33088
rect 520922 32600 520978 32609
rect 520922 32535 520978 32544
rect 520936 31657 520964 32535
rect 520922 31648 520978 31657
rect 520922 31583 520978 31592
rect 520922 31104 520978 31113
rect 520922 31039 520978 31048
rect 520936 30297 520964 31039
rect 520922 30288 520978 30297
rect 520922 30223 520978 30232
rect 117042 29880 117098 29889
rect 117042 29815 117098 29824
rect 116950 3768 117006 3777
rect 116950 3703 117006 3712
rect 117056 1154 117084 29815
rect 521106 29608 521162 29617
rect 521106 29543 521162 29552
rect 521120 28393 521148 29543
rect 521106 28384 521162 28393
rect 521106 28319 521162 28328
rect 117134 27976 117190 27985
rect 117134 27911 117190 27920
rect 117148 3505 117176 27911
rect 117226 24168 117282 24177
rect 117226 24103 117282 24112
rect 117134 3496 117190 3505
rect 117134 3431 117190 3440
rect 117044 1148 117096 1154
rect 117044 1090 117096 1096
rect 116860 1012 116912 1018
rect 116860 954 116912 960
rect 116676 876 116728 882
rect 116676 818 116728 824
rect 117240 814 117268 24103
rect 521106 21992 521162 22001
rect 521106 21927 521162 21936
rect 521120 20913 521148 21927
rect 521106 20904 521162 20913
rect 521106 20839 521162 20848
rect 520738 20496 520794 20505
rect 520738 20431 520794 20440
rect 520752 19553 520780 20431
rect 520738 19544 520794 19553
rect 520738 19479 520794 19488
rect 520922 19000 520978 19009
rect 520922 18935 520978 18944
rect 520936 18193 520964 18935
rect 520922 18184 520978 18193
rect 520922 18119 520978 18128
rect 521106 9344 521162 9353
rect 521106 9279 521162 9288
rect 521120 8265 521148 9279
rect 521106 8256 521162 8265
rect 521106 8191 521162 8200
rect 520370 7984 520426 7993
rect 520370 7919 520426 7928
rect 520384 6769 520412 7919
rect 520370 6760 520426 6769
rect 520370 6695 520426 6704
rect 521106 6624 521162 6633
rect 521106 6559 521162 6568
rect 521120 5273 521148 6559
rect 520922 5264 520978 5273
rect 520922 5199 520978 5208
rect 521106 5264 521162 5273
rect 521106 5199 521162 5208
rect 520936 3777 520964 5199
rect 521014 3904 521070 3913
rect 521014 3839 521070 3848
rect 520922 3768 520978 3777
rect 520922 3703 520978 3712
rect 143644 2514 143980 2530
rect 443656 2514 443992 2530
rect 143632 2508 143980 2514
rect 143684 2502 143980 2508
rect 425796 2508 425848 2514
rect 143632 2450 143684 2456
rect 425796 2450 425848 2456
rect 443644 2508 443992 2514
rect 443696 2502 443992 2508
rect 443644 2450 443696 2456
rect 193600 2094 193936 2122
rect 243648 2094 243984 2122
rect 293604 2094 293940 2122
rect 343652 2094 343988 2122
rect 393608 2094 393944 2122
rect 163778 1592 163834 1601
rect 163778 1527 163834 1536
rect 117228 808 117280 814
rect 163792 800 163820 1527
rect 193600 1494 193628 2094
rect 229282 1728 229338 1737
rect 229282 1663 229338 1672
rect 193588 1488 193640 1494
rect 193588 1430 193640 1436
rect 229296 800 229324 1663
rect 243648 1601 243676 2094
rect 293604 1737 293632 2094
rect 293590 1728 293646 1737
rect 293590 1663 293646 1672
rect 243634 1592 243690 1601
rect 243634 1527 243690 1536
rect 294786 1456 294842 1465
rect 343652 1426 343680 2094
rect 393608 1465 393636 2094
rect 360290 1456 360346 1465
rect 294786 1391 294788 1400
rect 294840 1391 294842 1400
rect 343640 1420 343692 1426
rect 294788 1362 294840 1368
rect 360290 1391 360346 1400
rect 393594 1456 393650 1465
rect 393594 1391 393650 1400
rect 343640 1362 343692 1368
rect 294800 800 294828 1362
rect 360304 800 360332 1391
rect 425808 800 425836 2450
rect 521028 2281 521056 3839
rect 521106 2680 521162 2689
rect 521106 2615 521162 2624
rect 521014 2272 521070 2281
rect 521014 2207 521070 2216
rect 493612 2094 493948 2122
rect 493612 1426 493640 2094
rect 491300 1420 491352 1426
rect 491300 1362 491352 1368
rect 493600 1420 493652 1426
rect 493600 1362 493652 1368
rect 491312 800 491340 1362
rect 117228 750 117280 756
rect 103796 740 103848 746
rect 103796 682 103848 688
rect 110788 740 110840 746
rect 110788 682 110840 688
rect 163778 -400 163834 800
rect 229282 -400 229338 800
rect 294786 -400 294842 800
rect 360290 -400 360346 800
rect 425794 -400 425850 800
rect 491298 -400 491354 800
rect 521120 785 521148 2615
rect 521106 776 521162 785
rect 521106 711 521162 720
<< via2 >>
rect 2962 153720 3018 153776
rect 16302 159296 16358 159352
rect 16578 153856 16634 153912
rect 19890 153992 19946 154048
rect 23018 159432 23074 159488
rect 12438 152496 12494 152552
rect 8850 152360 8906 152416
rect 6090 150592 6146 150648
rect 2686 150456 2742 150512
rect 28078 156576 28134 156632
rect 29826 159568 29882 159624
rect 31482 156712 31538 156768
rect 30378 154128 30434 154184
rect 33966 157936 34022 157992
rect 40682 158208 40738 158264
rect 44086 158072 44142 158128
rect 57518 158344 57574 158400
rect 55862 156848 55918 156904
rect 54298 154264 54354 154320
rect 65982 155488 66038 155544
rect 62578 155352 62634 155408
rect 72698 156984 72754 157040
rect 68466 155216 68522 155272
rect 76010 155760 76066 155816
rect 78586 155624 78642 155680
rect 85302 155896 85358 155952
rect 85578 154400 85634 154456
rect 104622 158480 104678 158536
rect 82818 149640 82874 149696
rect 109590 148008 109646 148064
rect 115570 157120 115626 157176
rect 111062 150456 111118 150512
rect 110970 147328 111026 147384
rect 110326 146376 110382 146432
rect 110326 106256 110382 106312
rect 111338 150592 111394 150648
rect 111706 147328 111762 147384
rect 113822 144200 113878 144256
rect 116122 145152 116178 145208
rect 116030 143248 116086 143304
rect 115294 141344 115350 141400
rect 116122 139440 116178 139496
rect 116122 137536 116178 137592
rect 115202 135496 115258 135552
rect 116030 133592 116086 133648
rect 114190 132776 114246 132832
rect 113914 121352 113970 121408
rect 114006 110064 114062 110120
rect 114098 98640 114154 98696
rect 114190 87216 114246 87272
rect 116122 131688 116178 131744
rect 116582 149640 116638 149696
rect 116490 129784 116546 129840
rect 116122 125976 116178 126032
rect 116122 124108 116124 124128
rect 116124 124108 116176 124128
rect 116176 124108 116178 124128
rect 116122 124072 116178 124108
rect 115938 122168 115994 122224
rect 116122 120128 116178 120184
rect 116122 118224 116178 118280
rect 116122 116320 116178 116376
rect 116122 114452 116124 114472
rect 116124 114452 116176 114472
rect 116176 114452 116178 114472
rect 116122 114416 116178 114452
rect 115938 112512 115994 112568
rect 116122 110608 116178 110664
rect 116122 108704 116178 108760
rect 116950 102856 117006 102912
rect 121458 153720 121514 153776
rect 121642 153720 121698 153776
rect 125966 152360 126022 152416
rect 126242 152360 126298 152416
rect 128542 152496 128598 152552
rect 131026 159296 131082 159352
rect 133602 159432 133658 159488
rect 131762 153856 131818 153912
rect 133602 153040 133658 153096
rect 134338 153992 134394 154048
rect 136270 153040 136326 153096
rect 138386 159568 138442 159624
rect 137926 153992 137982 154048
rect 138110 153584 138166 153640
rect 140134 156576 140190 156632
rect 143262 156712 143318 156768
rect 142158 154128 142214 154184
rect 142434 154148 142490 154184
rect 142434 154128 142436 154148
rect 142436 154128 142488 154148
rect 142488 154128 142490 154148
rect 143078 154128 143134 154184
rect 143538 153992 143594 154048
rect 143446 153584 143502 153640
rect 145102 157936 145158 157992
rect 143538 152360 143594 152416
rect 149610 158208 149666 158264
rect 152186 158072 152242 158128
rect 161570 156848 161626 156904
rect 160650 154264 160706 154320
rect 162858 158344 162914 158400
rect 166354 155352 166410 155408
rect 169022 155488 169078 155544
rect 171230 155216 171286 155272
rect 174082 156984 174138 157040
rect 176842 155760 176898 155816
rect 178682 155624 178738 155680
rect 183742 155896 183798 155952
rect 184386 154400 184442 154456
rect 192114 153720 192170 153776
rect 198738 158480 198794 158536
rect 200118 153348 200120 153368
rect 200120 153348 200172 153368
rect 200172 153348 200174 153368
rect 200118 153312 200174 153348
rect 200854 153332 200910 153368
rect 200854 153312 200856 153332
rect 200856 153312 200908 153332
rect 200908 153312 200910 153332
rect 204718 159296 204774 159352
rect 207018 157120 207074 157176
rect 211526 153720 211582 153776
rect 226798 152360 226854 152416
rect 274546 159432 274602 159488
rect 274822 159296 274878 159352
rect 280710 153720 280766 153776
rect 292578 152360 292634 152416
rect 313370 152360 313426 152416
rect 328550 159432 328606 159488
rect 357438 152360 357494 152416
rect 407670 152360 407726 152416
rect 427726 152652 427782 152688
rect 427726 152632 427728 152652
rect 427728 152632 427780 152652
rect 427780 152632 427782 152652
rect 431222 152496 431278 152552
rect 430302 152360 430358 152416
rect 430854 152360 430910 152416
rect 432970 152632 433026 152688
rect 432418 152260 432420 152280
rect 432420 152260 432472 152280
rect 432472 152260 432474 152280
rect 432418 152224 432474 152260
rect 432326 152088 432382 152144
rect 433062 152360 433118 152416
rect 432878 152224 432934 152280
rect 432970 152124 432972 152144
rect 432972 152124 433024 152144
rect 433024 152124 433026 152144
rect 432970 152088 433026 152124
rect 448518 152496 448574 152552
rect 519726 163104 519782 163160
rect 519542 161608 519598 161664
rect 519634 160112 519690 160168
rect 519542 147872 519598 147928
rect 519818 158616 519874 158672
rect 519726 149232 519782 149288
rect 519726 148008 519782 148064
rect 519634 146512 519690 146568
rect 519450 143384 519506 143440
rect 519358 141888 519414 141944
rect 519266 140392 519322 140448
rect 520002 157120 520058 157176
rect 519910 151000 519966 151056
rect 519818 145152 519874 145208
rect 520094 153992 520150 154048
rect 520002 143792 520058 143848
rect 521106 155624 521162 155680
rect 521014 152496 521070 152552
rect 520186 149504 520242 149560
rect 520094 141072 520150 141128
rect 520094 138896 520150 138952
rect 519910 138352 519966 138408
rect 520002 137400 520058 137456
rect 519910 135768 519966 135824
rect 519726 135632 519782 135688
rect 519818 134272 519874 134328
rect 519542 132776 519598 132832
rect 519450 131552 519506 131608
rect 519358 130192 519414 130248
rect 519266 128832 519322 128888
rect 519450 128288 519506 128344
rect 117226 127880 117282 127936
rect 519358 120536 519414 120592
rect 519726 131280 519782 131336
rect 519634 129784 519690 129840
rect 519542 122032 519598 122088
rect 520922 144880 520978 144936
rect 520186 136992 520242 137048
rect 521198 146512 521254 146568
rect 521106 142432 521162 142488
rect 521014 139712 521070 139768
rect 521198 134408 521254 134464
rect 520922 132912 520978 132968
rect 520094 127472 520150 127528
rect 520186 126656 520242 126712
rect 520002 126112 520058 126168
rect 520094 125160 520150 125216
rect 519910 124752 519966 124808
rect 520002 123664 520058 123720
rect 519818 123392 519874 123448
rect 519910 122168 519966 122224
rect 519726 120672 519782 120728
rect 519634 119312 519690 119368
rect 519818 119176 519874 119232
rect 519450 117952 519506 118008
rect 519726 117544 519782 117600
rect 519542 116048 519598 116104
rect 519358 111152 519414 111208
rect 519634 114552 519690 114608
rect 519542 107072 519598 107128
rect 520186 116592 520242 116648
rect 520094 115232 520150 115288
rect 520002 113872 520058 113928
rect 521106 113056 521162 113112
rect 519910 112512 519966 112568
rect 519818 109792 519874 109848
rect 519726 108432 519782 108488
rect 521014 108432 521070 108488
rect 520922 106936 520978 106992
rect 519634 105712 519690 105768
rect 520278 105440 520334 105496
rect 117134 104760 117190 104816
rect 117042 100952 117098 101008
rect 519818 99320 519874 99376
rect 116858 99048 116914 99104
rect 519726 97824 519782 97880
rect 116766 97144 116822 97200
rect 519266 96328 519322 96384
rect 116674 95240 116730 95296
rect 116582 93336 116638 93392
rect 116122 91296 116178 91352
rect 521566 111560 521622 111616
rect 521290 110064 521346 110120
rect 521106 104352 521162 104408
rect 521198 103944 521254 104000
rect 521106 102448 521162 102504
rect 521014 100272 521070 100328
rect 520922 98912 520978 98968
rect 520278 97552 520334 97608
rect 521566 102992 521622 103048
rect 521290 101632 521346 101688
rect 521474 100952 521530 101008
rect 521198 96192 521254 96248
rect 521106 94968 521162 95024
rect 519910 94832 519966 94888
rect 519818 92112 519874 92168
rect 519726 90752 519782 90808
rect 116122 89392 116178 89448
rect 519266 89392 519322 89448
rect 521474 93472 521530 93528
rect 520186 93336 520242 93392
rect 519910 88032 519966 88088
rect 116030 87488 116086 87544
rect 521290 91840 521346 91896
rect 520922 90208 520978 90264
rect 520186 86672 520242 86728
rect 520278 85720 520334 85776
rect 115202 85584 115258 85640
rect 116582 83680 116638 83736
rect 520186 82728 520242 82784
rect 116214 81776 116270 81832
rect 519634 81096 519690 81152
rect 115938 79872 115994 79928
rect 116122 77968 116178 78024
rect 519818 79600 519874 79656
rect 519726 76608 519782 76664
rect 519634 74568 519690 74624
rect 116674 74024 116730 74080
rect 116582 72120 116638 72176
rect 113362 64504 113418 64560
rect 110326 57976 110382 58032
rect 110326 56752 110382 56808
rect 110326 53896 110382 53952
rect 110326 52536 110382 52592
rect 110326 51040 110382 51096
rect 110326 48320 110382 48376
rect 110326 47096 110382 47152
rect 110326 45056 110382 45112
rect 110878 45056 110934 45112
rect 110326 44920 110382 44976
rect 110418 41384 110474 41440
rect 110326 37304 110382 37360
rect 110326 35264 110382 35320
rect 110326 35128 110382 35184
rect 109498 3576 109554 3632
rect 109406 3440 109462 3496
rect 109498 3304 109554 3360
rect 109406 2896 109462 2952
rect 33046 2624 33102 2680
rect 42062 2624 42118 2680
rect 42706 2624 42762 2680
rect 44730 2624 44786 2680
rect 62394 2624 62450 2680
rect 63038 2624 63094 2680
rect 64050 2624 64106 2680
rect 68282 2624 68338 2680
rect 78770 2624 78826 2680
rect 87050 2624 87106 2680
rect 90086 2624 90142 2680
rect 90362 2624 90418 2680
rect 91558 2624 91614 2680
rect 91926 2624 91982 2680
rect 93030 2624 93086 2680
rect 93858 2624 93914 2680
rect 95698 2624 95754 2680
rect 97722 2624 97778 2680
rect 97906 2624 97962 2680
rect 99194 2624 99250 2680
rect 103702 2624 103758 2680
rect 104438 2624 104494 2680
rect 104990 2624 105046 2680
rect 106186 2624 106242 2680
rect 106370 2624 106426 2680
rect 29550 2488 29606 2544
rect 26054 2352 26110 2408
rect 22926 2216 22982 2272
rect 5998 1808 6054 1864
rect 19614 2080 19670 2136
rect 16210 1944 16266 2000
rect 12622 1672 12678 1728
rect 9310 1536 9366 1592
rect 55954 1400 56010 1456
rect 87050 1264 87106 1320
rect 90362 1128 90418 1184
rect 90086 992 90142 1048
rect 95698 1264 95754 1320
rect 95974 1264 96030 1320
rect 97906 1264 97962 1320
rect 98274 1264 98330 1320
rect 97722 1128 97778 1184
rect 104438 2352 104494 2408
rect 104622 2352 104678 2408
rect 104438 2216 104494 2272
rect 104622 2216 104678 2272
rect 104346 2080 104402 2136
rect 104622 2080 104678 2136
rect 99378 1128 99434 1184
rect 102598 1128 102654 1184
rect 103702 1128 103758 1184
rect 110326 33768 110382 33824
rect 110418 29688 110474 29744
rect 110602 29824 110658 29880
rect 110786 37304 110842 37360
rect 110786 29688 110842 29744
rect 110510 28736 110566 28792
rect 110326 28600 110382 28656
rect 109866 2624 109922 2680
rect 110326 28056 110382 28112
rect 110326 27648 110382 27704
rect 110050 3848 110106 3904
rect 110050 3712 110106 3768
rect 110050 3032 110106 3088
rect 110326 27104 110382 27160
rect 110602 28056 110658 28112
rect 110970 44920 111026 44976
rect 111798 44240 111854 44296
rect 111062 35264 111118 35320
rect 111062 33768 111118 33824
rect 111062 29824 111118 29880
rect 111798 28736 111854 28792
rect 111062 28600 111118 28656
rect 110970 27648 111026 27704
rect 110878 27104 110934 27160
rect 110694 4120 110750 4176
rect 110326 2896 110382 2952
rect 110326 1808 110382 1864
rect 110786 3168 110842 3224
rect 110694 2896 110750 2952
rect 109866 1264 109922 1320
rect 109498 1128 109554 1184
rect 111062 992 111118 1048
rect 116306 70216 116362 70272
rect 116122 68312 116178 68368
rect 116582 66408 116638 66464
rect 519634 73616 519690 73672
rect 519542 68992 519598 69048
rect 116214 64504 116270 64560
rect 520002 78104 520058 78160
rect 519818 73208 519874 73264
rect 521198 87216 521254 87272
rect 521106 84224 521162 84280
rect 520922 82592 520978 82648
rect 520278 78512 520334 78568
rect 521382 88712 521438 88768
rect 521290 83952 521346 84008
rect 521382 81232 521438 81288
rect 521198 79872 521254 79928
rect 521106 77152 521162 77208
rect 520186 75928 520242 75984
rect 520094 75112 520150 75168
rect 520002 72392 520058 72448
rect 519726 70488 519782 70544
rect 519910 70488 519966 70544
rect 519634 67768 519690 67824
rect 519818 66000 519874 66056
rect 519542 63688 519598 63744
rect 116122 62600 116178 62656
rect 116582 60560 116638 60616
rect 114190 53080 114246 53136
rect 116122 43288 116178 43344
rect 114098 41792 114154 41848
rect 114006 30368 114062 30424
rect 116398 26016 116454 26072
rect 116306 20304 116362 20360
rect 113914 18944 113970 19000
rect 116214 18400 116270 18456
rect 116030 16360 116086 16416
rect 115938 12552 115994 12608
rect 113822 7656 113878 7712
rect 116122 14456 116178 14512
rect 116030 2352 116086 2408
rect 116490 22208 116546 22264
rect 116306 3304 116362 3360
rect 116306 3032 116362 3088
rect 116214 2488 116270 2544
rect 116122 2216 116178 2272
rect 115938 2080 115994 2136
rect 520186 71984 520242 72040
rect 520094 69128 520150 69184
rect 520002 67496 520058 67552
rect 519910 65048 519966 65104
rect 520186 66408 520242 66464
rect 521106 64504 521162 64560
rect 520738 62872 520794 62928
rect 520278 61376 520334 61432
rect 520002 60968 520058 61024
rect 519818 59608 519874 59664
rect 520186 56888 520242 56944
rect 521106 62328 521162 62384
rect 521014 59880 521070 59936
rect 520738 58248 520794 58304
rect 520370 56888 520426 56944
rect 520278 55392 520334 55448
rect 519266 53760 519322 53816
rect 520094 52264 520150 52320
rect 520002 50768 520058 50824
rect 519266 50088 519322 50144
rect 519450 47776 519506 47832
rect 521106 58384 521162 58440
rect 521014 55528 521070 55584
rect 521106 54168 521162 54224
rect 520370 52808 520426 52864
rect 520278 51448 520334 51504
rect 520186 49272 520242 49328
rect 520094 48728 520150 48784
rect 520002 47368 520058 47424
rect 519910 46280 519966 46336
rect 519450 44648 519506 44704
rect 519818 44648 519874 44704
rect 520186 46008 520242 46064
rect 519910 43288 519966 43344
rect 520186 43152 520242 43208
rect 519818 41928 519874 41984
rect 520094 41656 520150 41712
rect 116766 39480 116822 39536
rect 116674 37576 116730 37632
rect 520186 40568 520242 40624
rect 520186 40160 520242 40216
rect 520094 39208 520150 39264
rect 519818 38664 519874 38720
rect 520186 37848 520242 37904
rect 521566 37168 521622 37224
rect 519818 36488 519874 36544
rect 521566 35944 521622 36000
rect 521106 35536 521162 35592
rect 521106 34448 521162 34504
rect 520922 34040 520978 34096
rect 116950 33768 117006 33824
rect 116858 31728 116914 31784
rect 116766 3168 116822 3224
rect 520922 33088 520978 33144
rect 520922 32544 520978 32600
rect 520922 31592 520978 31648
rect 520922 31048 520978 31104
rect 520922 30232 520978 30288
rect 117042 29824 117098 29880
rect 116950 3712 117006 3768
rect 521106 29552 521162 29608
rect 521106 28328 521162 28384
rect 117134 27920 117190 27976
rect 117226 24112 117282 24168
rect 117134 3440 117190 3496
rect 521106 21936 521162 21992
rect 521106 20848 521162 20904
rect 520738 20440 520794 20496
rect 520738 19488 520794 19544
rect 520922 18944 520978 19000
rect 520922 18128 520978 18184
rect 521106 9288 521162 9344
rect 521106 8200 521162 8256
rect 520370 7928 520426 7984
rect 520370 6704 520426 6760
rect 521106 6568 521162 6624
rect 520922 5208 520978 5264
rect 521106 5208 521162 5264
rect 521014 3848 521070 3904
rect 520922 3712 520978 3768
rect 163778 1536 163834 1592
rect 229282 1672 229338 1728
rect 293590 1672 293646 1728
rect 243634 1536 243690 1592
rect 294786 1420 294842 1456
rect 294786 1400 294788 1420
rect 294788 1400 294840 1420
rect 294840 1400 294842 1420
rect 360290 1400 360346 1456
rect 393594 1400 393650 1456
rect 521106 2624 521162 2680
rect 521014 2216 521070 2272
rect 521106 720 521162 776
<< metal3 >>
rect 519721 163162 519787 163165
rect 523200 163162 524400 163192
rect 519721 163160 524400 163162
rect 519721 163104 519726 163160
rect 519782 163104 524400 163160
rect 519721 163102 524400 163104
rect 519721 163099 519787 163102
rect 523200 163072 524400 163102
rect 519537 161666 519603 161669
rect 523200 161666 524400 161696
rect 519537 161664 524400 161666
rect 519537 161608 519542 161664
rect 519598 161608 524400 161664
rect 519537 161606 524400 161608
rect 519537 161603 519603 161606
rect 523200 161576 524400 161606
rect 519629 160170 519695 160173
rect 523200 160170 524400 160200
rect 519629 160168 524400 160170
rect 519629 160112 519634 160168
rect 519690 160112 524400 160168
rect 519629 160110 524400 160112
rect 519629 160107 519695 160110
rect 523200 160080 524400 160110
rect 29821 159626 29887 159629
rect 138381 159626 138447 159629
rect 29821 159624 138447 159626
rect 29821 159568 29826 159624
rect 29882 159568 138386 159624
rect 138442 159568 138447 159624
rect 29821 159566 138447 159568
rect 29821 159563 29887 159566
rect 138381 159563 138447 159566
rect 23013 159490 23079 159493
rect 133597 159490 133663 159493
rect 23013 159488 133663 159490
rect 23013 159432 23018 159488
rect 23074 159432 133602 159488
rect 133658 159432 133663 159488
rect 23013 159430 133663 159432
rect 23013 159427 23079 159430
rect 133597 159427 133663 159430
rect 274541 159490 274607 159493
rect 328545 159490 328611 159493
rect 274541 159488 328611 159490
rect 274541 159432 274546 159488
rect 274602 159432 328550 159488
rect 328606 159432 328611 159488
rect 274541 159430 328611 159432
rect 274541 159427 274607 159430
rect 328545 159427 328611 159430
rect 16297 159354 16363 159357
rect 131021 159354 131087 159357
rect 16297 159352 131087 159354
rect 16297 159296 16302 159352
rect 16358 159296 131026 159352
rect 131082 159296 131087 159352
rect 16297 159294 131087 159296
rect 16297 159291 16363 159294
rect 131021 159291 131087 159294
rect 204713 159354 204779 159357
rect 274817 159354 274883 159357
rect 204713 159352 274883 159354
rect 204713 159296 204718 159352
rect 204774 159296 274822 159352
rect 274878 159296 274883 159352
rect 204713 159294 274883 159296
rect 204713 159291 204779 159294
rect 274817 159291 274883 159294
rect 519813 158674 519879 158677
rect 523200 158674 524400 158704
rect 519813 158672 524400 158674
rect 519813 158616 519818 158672
rect 519874 158616 524400 158672
rect 519813 158614 524400 158616
rect 519813 158611 519879 158614
rect 523200 158584 524400 158614
rect 104617 158538 104683 158541
rect 198733 158538 198799 158541
rect 104617 158536 198799 158538
rect 104617 158480 104622 158536
rect 104678 158480 198738 158536
rect 198794 158480 198799 158536
rect 104617 158478 198799 158480
rect 104617 158475 104683 158478
rect 198733 158475 198799 158478
rect 57513 158402 57579 158405
rect 162853 158402 162919 158405
rect 57513 158400 162919 158402
rect 57513 158344 57518 158400
rect 57574 158344 162858 158400
rect 162914 158344 162919 158400
rect 57513 158342 162919 158344
rect 57513 158339 57579 158342
rect 162853 158339 162919 158342
rect 40677 158266 40743 158269
rect 149605 158266 149671 158269
rect 40677 158264 149671 158266
rect 40677 158208 40682 158264
rect 40738 158208 149610 158264
rect 149666 158208 149671 158264
rect 40677 158206 149671 158208
rect 40677 158203 40743 158206
rect 149605 158203 149671 158206
rect 44081 158130 44147 158133
rect 152181 158130 152247 158133
rect 44081 158128 152247 158130
rect 44081 158072 44086 158128
rect 44142 158072 152186 158128
rect 152242 158072 152247 158128
rect 44081 158070 152247 158072
rect 44081 158067 44147 158070
rect 152181 158067 152247 158070
rect 33961 157994 34027 157997
rect 145097 157994 145163 157997
rect 33961 157992 145163 157994
rect 33961 157936 33966 157992
rect 34022 157936 145102 157992
rect 145158 157936 145163 157992
rect 33961 157934 145163 157936
rect 33961 157931 34027 157934
rect 145097 157931 145163 157934
rect 115565 157178 115631 157181
rect 207013 157178 207079 157181
rect 115565 157176 207079 157178
rect 115565 157120 115570 157176
rect 115626 157120 207018 157176
rect 207074 157120 207079 157176
rect 115565 157118 207079 157120
rect 115565 157115 115631 157118
rect 207013 157115 207079 157118
rect 519997 157178 520063 157181
rect 523200 157178 524400 157208
rect 519997 157176 524400 157178
rect 519997 157120 520002 157176
rect 520058 157120 524400 157176
rect 519997 157118 524400 157120
rect 519997 157115 520063 157118
rect 523200 157088 524400 157118
rect 72693 157042 72759 157045
rect 174077 157042 174143 157045
rect 72693 157040 174143 157042
rect 72693 156984 72698 157040
rect 72754 156984 174082 157040
rect 174138 156984 174143 157040
rect 72693 156982 174143 156984
rect 72693 156979 72759 156982
rect 174077 156979 174143 156982
rect 55857 156906 55923 156909
rect 161565 156906 161631 156909
rect 55857 156904 161631 156906
rect 55857 156848 55862 156904
rect 55918 156848 161570 156904
rect 161626 156848 161631 156904
rect 55857 156846 161631 156848
rect 55857 156843 55923 156846
rect 161565 156843 161631 156846
rect 31477 156770 31543 156773
rect 143257 156770 143323 156773
rect 31477 156768 143323 156770
rect 31477 156712 31482 156768
rect 31538 156712 143262 156768
rect 143318 156712 143323 156768
rect 31477 156710 143323 156712
rect 31477 156707 31543 156710
rect 143257 156707 143323 156710
rect 28073 156634 28139 156637
rect 140129 156634 140195 156637
rect 28073 156632 140195 156634
rect 28073 156576 28078 156632
rect 28134 156576 140134 156632
rect 140190 156576 140195 156632
rect 28073 156574 140195 156576
rect 28073 156571 28139 156574
rect 140129 156571 140195 156574
rect 85297 155954 85363 155957
rect 183737 155954 183803 155957
rect 85297 155952 183803 155954
rect 85297 155896 85302 155952
rect 85358 155896 183742 155952
rect 183798 155896 183803 155952
rect 85297 155894 183803 155896
rect 85297 155891 85363 155894
rect 183737 155891 183803 155894
rect 76005 155818 76071 155821
rect 176837 155818 176903 155821
rect 76005 155816 176903 155818
rect 76005 155760 76010 155816
rect 76066 155760 176842 155816
rect 176898 155760 176903 155816
rect 76005 155758 176903 155760
rect 76005 155755 76071 155758
rect 176837 155755 176903 155758
rect 78581 155682 78647 155685
rect 178677 155682 178743 155685
rect 78581 155680 178743 155682
rect 78581 155624 78586 155680
rect 78642 155624 178682 155680
rect 178738 155624 178743 155680
rect 78581 155622 178743 155624
rect 78581 155619 78647 155622
rect 178677 155619 178743 155622
rect 521101 155682 521167 155685
rect 523200 155682 524400 155712
rect 521101 155680 524400 155682
rect 521101 155624 521106 155680
rect 521162 155624 524400 155680
rect 521101 155622 524400 155624
rect 521101 155619 521167 155622
rect 523200 155592 524400 155622
rect 65977 155546 66043 155549
rect 169017 155546 169083 155549
rect 65977 155544 169083 155546
rect 65977 155488 65982 155544
rect 66038 155488 169022 155544
rect 169078 155488 169083 155544
rect 65977 155486 169083 155488
rect 65977 155483 66043 155486
rect 169017 155483 169083 155486
rect 62573 155410 62639 155413
rect 166349 155410 166415 155413
rect 62573 155408 166415 155410
rect 62573 155352 62578 155408
rect 62634 155352 166354 155408
rect 166410 155352 166415 155408
rect 62573 155350 166415 155352
rect 62573 155347 62639 155350
rect 166349 155347 166415 155350
rect 68461 155274 68527 155277
rect 171225 155274 171291 155277
rect 68461 155272 171291 155274
rect 68461 155216 68466 155272
rect 68522 155216 171230 155272
rect 171286 155216 171291 155272
rect 68461 155214 171291 155216
rect 68461 155211 68527 155214
rect 171225 155211 171291 155214
rect 85573 154458 85639 154461
rect 184381 154458 184447 154461
rect 85573 154456 184447 154458
rect 85573 154400 85578 154456
rect 85634 154400 184386 154456
rect 184442 154400 184447 154456
rect 85573 154398 184447 154400
rect 85573 154395 85639 154398
rect 184381 154395 184447 154398
rect 54293 154322 54359 154325
rect 160645 154322 160711 154325
rect 54293 154320 160711 154322
rect 54293 154264 54298 154320
rect 54354 154264 160650 154320
rect 160706 154264 160711 154320
rect 54293 154262 160711 154264
rect 54293 154259 54359 154262
rect 160645 154259 160711 154262
rect 30373 154186 30439 154189
rect 142153 154186 142219 154189
rect 30373 154184 142219 154186
rect 30373 154128 30378 154184
rect 30434 154128 142158 154184
rect 142214 154128 142219 154184
rect 30373 154126 142219 154128
rect 30373 154123 30439 154126
rect 142153 154123 142219 154126
rect 142429 154186 142495 154189
rect 143073 154186 143139 154189
rect 142429 154184 143139 154186
rect 142429 154128 142434 154184
rect 142490 154128 143078 154184
rect 143134 154128 143139 154184
rect 142429 154126 143139 154128
rect 142429 154123 142495 154126
rect 143073 154123 143139 154126
rect 19885 154050 19951 154053
rect 134333 154050 134399 154053
rect 19885 154048 134399 154050
rect 19885 153992 19890 154048
rect 19946 153992 134338 154048
rect 134394 153992 134399 154048
rect 19885 153990 134399 153992
rect 19885 153987 19951 153990
rect 134333 153987 134399 153990
rect 137921 154050 137987 154053
rect 143533 154050 143599 154053
rect 137921 154048 143599 154050
rect 137921 153992 137926 154048
rect 137982 153992 143538 154048
rect 143594 153992 143599 154048
rect 137921 153990 143599 153992
rect 137921 153987 137987 153990
rect 143533 153987 143599 153990
rect 520089 154050 520155 154053
rect 523200 154050 524400 154080
rect 520089 154048 524400 154050
rect 520089 153992 520094 154048
rect 520150 153992 524400 154048
rect 520089 153990 524400 153992
rect 520089 153987 520155 153990
rect 523200 153960 524400 153990
rect 16573 153914 16639 153917
rect 131757 153914 131823 153917
rect 16573 153912 131823 153914
rect 16573 153856 16578 153912
rect 16634 153856 131762 153912
rect 131818 153856 131823 153912
rect 16573 153854 131823 153856
rect 16573 153851 16639 153854
rect 131757 153851 131823 153854
rect 2957 153778 3023 153781
rect 121453 153778 121519 153781
rect 2957 153776 121519 153778
rect 2957 153720 2962 153776
rect 3018 153720 121458 153776
rect 121514 153720 121519 153776
rect 2957 153718 121519 153720
rect 2957 153715 3023 153718
rect 121453 153715 121519 153718
rect 121637 153778 121703 153781
rect 192109 153778 192175 153781
rect 121637 153776 192175 153778
rect 121637 153720 121642 153776
rect 121698 153720 192114 153776
rect 192170 153720 192175 153776
rect 121637 153718 192175 153720
rect 121637 153715 121703 153718
rect 192109 153715 192175 153718
rect 211521 153778 211587 153781
rect 280705 153778 280771 153781
rect 211521 153776 280771 153778
rect 211521 153720 211526 153776
rect 211582 153720 280710 153776
rect 280766 153720 280771 153776
rect 211521 153718 280771 153720
rect 211521 153715 211587 153718
rect 280705 153715 280771 153718
rect 138105 153642 138171 153645
rect 143441 153642 143507 153645
rect 138105 153640 143507 153642
rect 138105 153584 138110 153640
rect 138166 153584 143446 153640
rect 143502 153584 143507 153640
rect 138105 153582 143507 153584
rect 138105 153579 138171 153582
rect 143441 153579 143507 153582
rect 200113 153370 200179 153373
rect 200849 153370 200915 153373
rect 200113 153368 200915 153370
rect 200113 153312 200118 153368
rect 200174 153312 200854 153368
rect 200910 153312 200915 153368
rect 200113 153310 200915 153312
rect 200113 153307 200179 153310
rect 200849 153307 200915 153310
rect 133597 153098 133663 153101
rect 136265 153098 136331 153101
rect 133597 153096 136331 153098
rect 133597 153040 133602 153096
rect 133658 153040 136270 153096
rect 136326 153040 136331 153096
rect 133597 153038 136331 153040
rect 133597 153035 133663 153038
rect 136265 153035 136331 153038
rect 427721 152690 427787 152693
rect 432965 152690 433031 152693
rect 427721 152688 433031 152690
rect 427721 152632 427726 152688
rect 427782 152632 432970 152688
rect 433026 152632 433031 152688
rect 427721 152630 433031 152632
rect 427721 152627 427787 152630
rect 432965 152627 433031 152630
rect 12433 152554 12499 152557
rect 128537 152554 128603 152557
rect 12433 152552 128603 152554
rect 12433 152496 12438 152552
rect 12494 152496 128542 152552
rect 128598 152496 128603 152552
rect 12433 152494 128603 152496
rect 12433 152491 12499 152494
rect 128537 152491 128603 152494
rect 431217 152554 431283 152557
rect 448513 152554 448579 152557
rect 431217 152552 448579 152554
rect 431217 152496 431222 152552
rect 431278 152496 448518 152552
rect 448574 152496 448579 152552
rect 431217 152494 448579 152496
rect 431217 152491 431283 152494
rect 448513 152491 448579 152494
rect 521009 152554 521075 152557
rect 523200 152554 524400 152584
rect 521009 152552 524400 152554
rect 521009 152496 521014 152552
rect 521070 152496 524400 152552
rect 521009 152494 524400 152496
rect 521009 152491 521075 152494
rect 523200 152464 524400 152494
rect 8845 152418 8911 152421
rect 125961 152418 126027 152421
rect 8845 152416 126027 152418
rect 8845 152360 8850 152416
rect 8906 152360 125966 152416
rect 126022 152360 126027 152416
rect 8845 152358 126027 152360
rect 8845 152355 8911 152358
rect 125961 152355 126027 152358
rect 126237 152418 126303 152421
rect 143533 152418 143599 152421
rect 126237 152416 143599 152418
rect 126237 152360 126242 152416
rect 126298 152360 143538 152416
rect 143594 152360 143599 152416
rect 126237 152358 143599 152360
rect 126237 152355 126303 152358
rect 143533 152355 143599 152358
rect 226793 152418 226859 152421
rect 292573 152418 292639 152421
rect 226793 152416 292639 152418
rect 226793 152360 226798 152416
rect 226854 152360 292578 152416
rect 292634 152360 292639 152416
rect 226793 152358 292639 152360
rect 226793 152355 226859 152358
rect 292573 152355 292639 152358
rect 313365 152418 313431 152421
rect 357433 152418 357499 152421
rect 313365 152416 357499 152418
rect 313365 152360 313370 152416
rect 313426 152360 357438 152416
rect 357494 152360 357499 152416
rect 313365 152358 357499 152360
rect 313365 152355 313431 152358
rect 357433 152355 357499 152358
rect 407665 152418 407731 152421
rect 430297 152418 430363 152421
rect 407665 152416 430363 152418
rect 407665 152360 407670 152416
rect 407726 152360 430302 152416
rect 430358 152360 430363 152416
rect 407665 152358 430363 152360
rect 407665 152355 407731 152358
rect 430297 152355 430363 152358
rect 430849 152418 430915 152421
rect 433057 152418 433123 152421
rect 430849 152416 433123 152418
rect 430849 152360 430854 152416
rect 430910 152360 433062 152416
rect 433118 152360 433123 152416
rect 430849 152358 433123 152360
rect 430849 152355 430915 152358
rect 433057 152355 433123 152358
rect 432413 152282 432479 152285
rect 432873 152282 432939 152285
rect 432413 152280 432939 152282
rect 432413 152224 432418 152280
rect 432474 152224 432878 152280
rect 432934 152224 432939 152280
rect 432413 152222 432939 152224
rect 432413 152219 432479 152222
rect 432873 152219 432939 152222
rect 432321 152146 432387 152149
rect 432965 152146 433031 152149
rect 432321 152144 433031 152146
rect 432321 152088 432326 152144
rect 432382 152088 432970 152144
rect 433026 152088 433031 152144
rect 432321 152086 433031 152088
rect 432321 152083 432387 152086
rect 432965 152083 433031 152086
rect 519905 151058 519971 151061
rect 523200 151058 524400 151088
rect 519905 151056 524400 151058
rect 519905 151000 519910 151056
rect 519966 151000 524400 151056
rect 519905 150998 524400 151000
rect 519905 150995 519971 150998
rect 523200 150968 524400 150998
rect 6085 150650 6151 150653
rect 111333 150650 111399 150653
rect 6085 150648 111399 150650
rect 6085 150592 6090 150648
rect 6146 150592 111338 150648
rect 111394 150592 111399 150648
rect 6085 150590 111399 150592
rect 6085 150587 6151 150590
rect 111333 150587 111399 150590
rect 2681 150514 2747 150517
rect 111057 150514 111123 150517
rect 2681 150512 111123 150514
rect 2681 150456 2686 150512
rect 2742 150456 111062 150512
rect 111118 150456 111123 150512
rect 2681 150454 111123 150456
rect 2681 150451 2747 150454
rect 111057 150451 111123 150454
rect 82813 149698 82879 149701
rect 116577 149698 116643 149701
rect 82813 149696 116643 149698
rect 82813 149640 82818 149696
rect 82874 149640 116582 149696
rect 116638 149640 116643 149696
rect 82813 149638 116643 149640
rect 82813 149635 82879 149638
rect 116577 149635 116643 149638
rect 520181 149562 520247 149565
rect 523200 149562 524400 149592
rect 520181 149560 524400 149562
rect 520181 149504 520186 149560
rect 520242 149504 524400 149560
rect 520181 149502 524400 149504
rect 520181 149499 520247 149502
rect 523200 149472 524400 149502
rect 519721 149290 519787 149293
rect 518788 149288 519787 149290
rect 518788 149232 519726 149288
rect 519782 149232 519787 149288
rect 518788 149230 519787 149232
rect 519721 149227 519787 149230
rect 109585 148066 109651 148069
rect 119110 148066 119170 148988
rect 109585 148064 119170 148066
rect 109585 148008 109590 148064
rect 109646 148008 119170 148064
rect 109585 148006 119170 148008
rect 519721 148066 519787 148069
rect 523200 148066 524400 148096
rect 519721 148064 524400 148066
rect 519721 148008 519726 148064
rect 519782 148008 524400 148064
rect 519721 148006 524400 148008
rect 109585 148003 109651 148006
rect 519721 148003 519787 148006
rect 523200 147976 524400 148006
rect 519537 147930 519603 147933
rect 518788 147928 519603 147930
rect 518788 147872 519542 147928
rect 519598 147872 519603 147928
rect 518788 147870 519603 147872
rect 519537 147867 519603 147870
rect 110965 147386 111031 147389
rect 111701 147386 111767 147389
rect 110965 147384 111767 147386
rect 110965 147328 110970 147384
rect 111026 147328 111706 147384
rect 111762 147328 111767 147384
rect 110965 147326 111767 147328
rect 110965 147323 111031 147326
rect 111701 147323 111767 147326
rect 110321 146434 110387 146437
rect 119110 146434 119170 147084
rect 519629 146570 519695 146573
rect 518788 146568 519695 146570
rect 518788 146512 519634 146568
rect 519690 146512 519695 146568
rect 518788 146510 519695 146512
rect 519629 146507 519695 146510
rect 521193 146570 521259 146573
rect 523200 146570 524400 146600
rect 521193 146568 524400 146570
rect 521193 146512 521198 146568
rect 521254 146512 524400 146568
rect 521193 146510 524400 146512
rect 521193 146507 521259 146510
rect 523200 146480 524400 146510
rect 110321 146432 119170 146434
rect 110321 146376 110326 146432
rect 110382 146376 119170 146432
rect 110321 146374 119170 146376
rect 110321 146371 110387 146374
rect 116117 145210 116183 145213
rect 519813 145210 519879 145213
rect 116117 145208 119140 145210
rect 116117 145152 116122 145208
rect 116178 145152 119140 145208
rect 116117 145150 119140 145152
rect 518788 145208 519879 145210
rect 518788 145152 519818 145208
rect 519874 145152 519879 145208
rect 518788 145150 519879 145152
rect 116117 145147 116183 145150
rect 519813 145147 519879 145150
rect 520917 144938 520983 144941
rect 523200 144938 524400 144968
rect 520917 144936 524400 144938
rect 520917 144880 520922 144936
rect 520978 144880 524400 144936
rect 520917 144878 524400 144880
rect 520917 144875 520983 144878
rect 523200 144848 524400 144878
rect 113817 144258 113883 144261
rect 110860 144256 113883 144258
rect 110860 144200 113822 144256
rect 113878 144200 113883 144256
rect 110860 144198 113883 144200
rect 113817 144195 113883 144198
rect 519997 143850 520063 143853
rect 518788 143848 520063 143850
rect 518788 143792 520002 143848
rect 520058 143792 520063 143848
rect 518788 143790 520063 143792
rect 519997 143787 520063 143790
rect 519445 143442 519511 143445
rect 523200 143442 524400 143472
rect 519445 143440 524400 143442
rect 519445 143384 519450 143440
rect 519506 143384 524400 143440
rect 519445 143382 524400 143384
rect 519445 143379 519511 143382
rect 523200 143352 524400 143382
rect 116025 143306 116091 143309
rect 116025 143304 119140 143306
rect 116025 143248 116030 143304
rect 116086 143248 119140 143304
rect 116025 143246 119140 143248
rect 116025 143243 116091 143246
rect 521101 142490 521167 142493
rect 518788 142488 521167 142490
rect 518788 142432 521106 142488
rect 521162 142432 521167 142488
rect 518788 142430 521167 142432
rect 521101 142427 521167 142430
rect 519353 141946 519419 141949
rect 523200 141946 524400 141976
rect 519353 141944 524400 141946
rect 519353 141888 519358 141944
rect 519414 141888 524400 141944
rect 519353 141886 524400 141888
rect 519353 141883 519419 141886
rect 523200 141856 524400 141886
rect 115289 141402 115355 141405
rect 115289 141400 119140 141402
rect 115289 141344 115294 141400
rect 115350 141344 119140 141400
rect 115289 141342 119140 141344
rect 115289 141339 115355 141342
rect 520089 141130 520155 141133
rect 518788 141128 520155 141130
rect 518788 141072 520094 141128
rect 520150 141072 520155 141128
rect 518788 141070 520155 141072
rect 520089 141067 520155 141070
rect 519261 140450 519327 140453
rect 523200 140450 524400 140480
rect 519261 140448 524400 140450
rect 519261 140392 519266 140448
rect 519322 140392 524400 140448
rect 519261 140390 524400 140392
rect 519261 140387 519327 140390
rect 523200 140360 524400 140390
rect 521009 139770 521075 139773
rect 518788 139768 521075 139770
rect 518788 139712 521014 139768
rect 521070 139712 521075 139768
rect 518788 139710 521075 139712
rect 521009 139707 521075 139710
rect 116117 139498 116183 139501
rect 116117 139496 119140 139498
rect 116117 139440 116122 139496
rect 116178 139440 119140 139496
rect 116117 139438 119140 139440
rect 116117 139435 116183 139438
rect 520089 138954 520155 138957
rect 523200 138954 524400 138984
rect 520089 138952 524400 138954
rect 520089 138896 520094 138952
rect 520150 138896 524400 138952
rect 520089 138894 524400 138896
rect 520089 138891 520155 138894
rect 523200 138864 524400 138894
rect 519905 138410 519971 138413
rect 518788 138408 519971 138410
rect 518788 138352 519910 138408
rect 519966 138352 519971 138408
rect 518788 138350 519971 138352
rect 519905 138347 519971 138350
rect 116117 137594 116183 137597
rect 116117 137592 119140 137594
rect 116117 137536 116122 137592
rect 116178 137536 119140 137592
rect 116117 137534 119140 137536
rect 116117 137531 116183 137534
rect 519997 137458 520063 137461
rect 523200 137458 524400 137488
rect 519997 137456 524400 137458
rect 519997 137400 520002 137456
rect 520058 137400 524400 137456
rect 519997 137398 524400 137400
rect 519997 137395 520063 137398
rect 523200 137368 524400 137398
rect 520181 137050 520247 137053
rect 518788 137048 520247 137050
rect 518788 136992 520186 137048
rect 520242 136992 520247 137048
rect 518788 136990 520247 136992
rect 520181 136987 520247 136990
rect 519905 135826 519971 135829
rect 523200 135826 524400 135856
rect 519905 135824 524400 135826
rect 519905 135768 519910 135824
rect 519966 135768 524400 135824
rect 519905 135766 524400 135768
rect 519905 135763 519971 135766
rect 523200 135736 524400 135766
rect 519721 135690 519787 135693
rect 518788 135688 519787 135690
rect 518788 135632 519726 135688
rect 519782 135632 519787 135688
rect 518788 135630 519787 135632
rect 519721 135627 519787 135630
rect 115197 135554 115263 135557
rect 115197 135552 119140 135554
rect 115197 135496 115202 135552
rect 115258 135496 119140 135552
rect 115197 135494 119140 135496
rect 115197 135491 115263 135494
rect 521193 134466 521259 134469
rect 518758 134464 521259 134466
rect 518758 134408 521198 134464
rect 521254 134408 521259 134464
rect 518758 134406 521259 134408
rect 518758 134300 518818 134406
rect 521193 134403 521259 134406
rect 519813 134330 519879 134333
rect 523200 134330 524400 134360
rect 519813 134328 524400 134330
rect 519813 134272 519818 134328
rect 519874 134272 524400 134328
rect 519813 134270 524400 134272
rect 519813 134267 519879 134270
rect 523200 134240 524400 134270
rect 116025 133650 116091 133653
rect 116025 133648 119140 133650
rect 116025 133592 116030 133648
rect 116086 133592 119140 133648
rect 116025 133590 119140 133592
rect 116025 133587 116091 133590
rect 520917 132970 520983 132973
rect 518788 132968 520983 132970
rect 518788 132912 520922 132968
rect 520978 132912 520983 132968
rect 518788 132910 520983 132912
rect 520917 132907 520983 132910
rect 114185 132834 114251 132837
rect 110860 132832 114251 132834
rect 110860 132776 114190 132832
rect 114246 132776 114251 132832
rect 110860 132774 114251 132776
rect 114185 132771 114251 132774
rect 519537 132834 519603 132837
rect 523200 132834 524400 132864
rect 519537 132832 524400 132834
rect 519537 132776 519542 132832
rect 519598 132776 524400 132832
rect 519537 132774 524400 132776
rect 519537 132771 519603 132774
rect 523200 132744 524400 132774
rect 116117 131746 116183 131749
rect 116117 131744 119140 131746
rect 116117 131688 116122 131744
rect 116178 131688 119140 131744
rect 116117 131686 119140 131688
rect 116117 131683 116183 131686
rect 519445 131610 519511 131613
rect 518788 131608 519511 131610
rect 518788 131552 519450 131608
rect 519506 131552 519511 131608
rect 518788 131550 519511 131552
rect 519445 131547 519511 131550
rect 519721 131338 519787 131341
rect 523200 131338 524400 131368
rect 519721 131336 524400 131338
rect 519721 131280 519726 131336
rect 519782 131280 524400 131336
rect 519721 131278 524400 131280
rect 519721 131275 519787 131278
rect 523200 131248 524400 131278
rect 519353 130250 519419 130253
rect 518788 130248 519419 130250
rect 518788 130192 519358 130248
rect 519414 130192 519419 130248
rect 518788 130190 519419 130192
rect 519353 130187 519419 130190
rect 116485 129842 116551 129845
rect 519629 129842 519695 129845
rect 523200 129842 524400 129872
rect 116485 129840 119140 129842
rect 116485 129784 116490 129840
rect 116546 129784 119140 129840
rect 116485 129782 119140 129784
rect 519629 129840 524400 129842
rect 519629 129784 519634 129840
rect 519690 129784 524400 129840
rect 519629 129782 524400 129784
rect 116485 129779 116551 129782
rect 519629 129779 519695 129782
rect 523200 129752 524400 129782
rect 519261 128890 519327 128893
rect 518788 128888 519327 128890
rect 518788 128832 519266 128888
rect 519322 128832 519327 128888
rect 518788 128830 519327 128832
rect 519261 128827 519327 128830
rect 519445 128346 519511 128349
rect 523200 128346 524400 128376
rect 519445 128344 524400 128346
rect 519445 128288 519450 128344
rect 519506 128288 524400 128344
rect 519445 128286 524400 128288
rect 519445 128283 519511 128286
rect 523200 128256 524400 128286
rect 117221 127938 117287 127941
rect 117221 127936 119140 127938
rect 117221 127880 117226 127936
rect 117282 127880 119140 127936
rect 117221 127878 119140 127880
rect 117221 127875 117287 127878
rect 520089 127530 520155 127533
rect 518788 127528 520155 127530
rect 518788 127472 520094 127528
rect 520150 127472 520155 127528
rect 518788 127470 520155 127472
rect 520089 127467 520155 127470
rect 520181 126714 520247 126717
rect 523200 126714 524400 126744
rect 520181 126712 524400 126714
rect 520181 126656 520186 126712
rect 520242 126656 524400 126712
rect 520181 126654 524400 126656
rect 520181 126651 520247 126654
rect 523200 126624 524400 126654
rect 519997 126170 520063 126173
rect 518788 126168 520063 126170
rect 518788 126112 520002 126168
rect 520058 126112 520063 126168
rect 518788 126110 520063 126112
rect 519997 126107 520063 126110
rect 116117 126034 116183 126037
rect 116117 126032 119140 126034
rect 116117 125976 116122 126032
rect 116178 125976 119140 126032
rect 116117 125974 119140 125976
rect 116117 125971 116183 125974
rect 520089 125218 520155 125221
rect 523200 125218 524400 125248
rect 520089 125216 524400 125218
rect 520089 125160 520094 125216
rect 520150 125160 524400 125216
rect 520089 125158 524400 125160
rect 520089 125155 520155 125158
rect 523200 125128 524400 125158
rect 519905 124810 519971 124813
rect 518788 124808 519971 124810
rect 518788 124752 519910 124808
rect 519966 124752 519971 124808
rect 518788 124750 519971 124752
rect 519905 124747 519971 124750
rect 116117 124130 116183 124133
rect 116117 124128 119140 124130
rect 116117 124072 116122 124128
rect 116178 124072 119140 124128
rect 116117 124070 119140 124072
rect 116117 124067 116183 124070
rect 519997 123722 520063 123725
rect 523200 123722 524400 123752
rect 519997 123720 524400 123722
rect 519997 123664 520002 123720
rect 520058 123664 524400 123720
rect 519997 123662 524400 123664
rect 519997 123659 520063 123662
rect 523200 123632 524400 123662
rect 519813 123450 519879 123453
rect 518788 123448 519879 123450
rect 518788 123392 519818 123448
rect 519874 123392 519879 123448
rect 518788 123390 519879 123392
rect 519813 123387 519879 123390
rect 115933 122226 115999 122229
rect 519905 122226 519971 122229
rect 523200 122226 524400 122256
rect 115933 122224 119140 122226
rect 115933 122168 115938 122224
rect 115994 122168 119140 122224
rect 115933 122166 119140 122168
rect 519905 122224 524400 122226
rect 519905 122168 519910 122224
rect 519966 122168 524400 122224
rect 519905 122166 524400 122168
rect 115933 122163 115999 122166
rect 519905 122163 519971 122166
rect 523200 122136 524400 122166
rect 519537 122090 519603 122093
rect 518788 122088 519603 122090
rect 518788 122032 519542 122088
rect 519598 122032 519603 122088
rect 518788 122030 519603 122032
rect 519537 122027 519603 122030
rect 113909 121410 113975 121413
rect 110860 121408 113975 121410
rect 110860 121352 113914 121408
rect 113970 121352 113975 121408
rect 110860 121350 113975 121352
rect 113909 121347 113975 121350
rect 519721 120730 519787 120733
rect 523200 120730 524400 120760
rect 518788 120728 519787 120730
rect 518788 120672 519726 120728
rect 519782 120672 519787 120728
rect 518788 120670 519787 120672
rect 519721 120667 519787 120670
rect 519862 120670 524400 120730
rect 519353 120594 519419 120597
rect 519862 120594 519922 120670
rect 523200 120640 524400 120670
rect 519353 120592 519922 120594
rect 519353 120536 519358 120592
rect 519414 120536 519922 120592
rect 519353 120534 519922 120536
rect 519353 120531 519419 120534
rect 116117 120186 116183 120189
rect 116117 120184 119140 120186
rect 116117 120128 116122 120184
rect 116178 120128 119140 120184
rect 116117 120126 119140 120128
rect 116117 120123 116183 120126
rect 519629 119370 519695 119373
rect 518788 119368 519695 119370
rect 518788 119312 519634 119368
rect 519690 119312 519695 119368
rect 518788 119310 519695 119312
rect 519629 119307 519695 119310
rect 519813 119234 519879 119237
rect 523200 119234 524400 119264
rect 519813 119232 524400 119234
rect 519813 119176 519818 119232
rect 519874 119176 524400 119232
rect 519813 119174 524400 119176
rect 519813 119171 519879 119174
rect 523200 119144 524400 119174
rect 116117 118282 116183 118285
rect 116117 118280 119140 118282
rect 116117 118224 116122 118280
rect 116178 118224 119140 118280
rect 116117 118222 119140 118224
rect 116117 118219 116183 118222
rect 519445 118010 519511 118013
rect 518788 118008 519511 118010
rect 518788 117952 519450 118008
rect 519506 117952 519511 118008
rect 518788 117950 519511 117952
rect 519445 117947 519511 117950
rect 519721 117602 519787 117605
rect 523200 117602 524400 117632
rect 519721 117600 524400 117602
rect 519721 117544 519726 117600
rect 519782 117544 524400 117600
rect 519721 117542 524400 117544
rect 519721 117539 519787 117542
rect 523200 117512 524400 117542
rect 520181 116650 520247 116653
rect 518788 116648 520247 116650
rect 518788 116592 520186 116648
rect 520242 116592 520247 116648
rect 518788 116590 520247 116592
rect 520181 116587 520247 116590
rect 116117 116378 116183 116381
rect 116117 116376 119140 116378
rect 116117 116320 116122 116376
rect 116178 116320 119140 116376
rect 116117 116318 119140 116320
rect 116117 116315 116183 116318
rect 519537 116106 519603 116109
rect 523200 116106 524400 116136
rect 519537 116104 524400 116106
rect 519537 116048 519542 116104
rect 519598 116048 524400 116104
rect 519537 116046 524400 116048
rect 519537 116043 519603 116046
rect 523200 116016 524400 116046
rect 520089 115290 520155 115293
rect 518788 115288 520155 115290
rect 518788 115232 520094 115288
rect 520150 115232 520155 115288
rect 518788 115230 520155 115232
rect 520089 115227 520155 115230
rect 519629 114610 519695 114613
rect 523200 114610 524400 114640
rect 519629 114608 524400 114610
rect 519629 114552 519634 114608
rect 519690 114552 524400 114608
rect 519629 114550 524400 114552
rect 519629 114547 519695 114550
rect 523200 114520 524400 114550
rect 116117 114474 116183 114477
rect 116117 114472 119140 114474
rect 116117 114416 116122 114472
rect 116178 114416 119140 114472
rect 116117 114414 119140 114416
rect 116117 114411 116183 114414
rect 519997 113930 520063 113933
rect 518788 113928 520063 113930
rect 518788 113872 520002 113928
rect 520058 113872 520063 113928
rect 518788 113870 520063 113872
rect 519997 113867 520063 113870
rect 521101 113114 521167 113117
rect 523200 113114 524400 113144
rect 521101 113112 524400 113114
rect 521101 113056 521106 113112
rect 521162 113056 524400 113112
rect 521101 113054 524400 113056
rect 521101 113051 521167 113054
rect 523200 113024 524400 113054
rect 115933 112570 115999 112573
rect 519905 112570 519971 112573
rect 115933 112568 119140 112570
rect 115933 112512 115938 112568
rect 115994 112512 119140 112568
rect 115933 112510 119140 112512
rect 518788 112568 519971 112570
rect 518788 112512 519910 112568
rect 519966 112512 519971 112568
rect 518788 112510 519971 112512
rect 115933 112507 115999 112510
rect 519905 112507 519971 112510
rect 521561 111618 521627 111621
rect 523200 111618 524400 111648
rect 521561 111616 524400 111618
rect 521561 111560 521566 111616
rect 521622 111560 524400 111616
rect 521561 111558 524400 111560
rect 521561 111555 521627 111558
rect 523200 111528 524400 111558
rect 519353 111210 519419 111213
rect 518788 111208 519419 111210
rect 518788 111152 519358 111208
rect 519414 111152 519419 111208
rect 518788 111150 519419 111152
rect 519353 111147 519419 111150
rect 116117 110666 116183 110669
rect 116117 110664 119140 110666
rect 116117 110608 116122 110664
rect 116178 110608 119140 110664
rect 116117 110606 119140 110608
rect 116117 110603 116183 110606
rect 114001 110122 114067 110125
rect 110860 110120 114067 110122
rect 110860 110064 114006 110120
rect 114062 110064 114067 110120
rect 110860 110062 114067 110064
rect 114001 110059 114067 110062
rect 521285 110122 521351 110125
rect 523200 110122 524400 110152
rect 521285 110120 524400 110122
rect 521285 110064 521290 110120
rect 521346 110064 524400 110120
rect 521285 110062 524400 110064
rect 521285 110059 521351 110062
rect 523200 110032 524400 110062
rect 519813 109850 519879 109853
rect 518788 109848 519879 109850
rect 518788 109792 519818 109848
rect 519874 109792 519879 109848
rect 518788 109790 519879 109792
rect 519813 109787 519879 109790
rect 116117 108762 116183 108765
rect 116117 108760 119140 108762
rect 116117 108704 116122 108760
rect 116178 108704 119140 108760
rect 116117 108702 119140 108704
rect 116117 108699 116183 108702
rect 519721 108490 519787 108493
rect 518788 108488 519787 108490
rect 518788 108432 519726 108488
rect 519782 108432 519787 108488
rect 518788 108430 519787 108432
rect 519721 108427 519787 108430
rect 521009 108490 521075 108493
rect 523200 108490 524400 108520
rect 521009 108488 524400 108490
rect 521009 108432 521014 108488
rect 521070 108432 524400 108488
rect 521009 108430 524400 108432
rect 521009 108427 521075 108430
rect 523200 108400 524400 108430
rect 519537 107130 519603 107133
rect 518788 107128 519603 107130
rect 518788 107072 519542 107128
rect 519598 107072 519603 107128
rect 518788 107070 519603 107072
rect 519537 107067 519603 107070
rect 520917 106994 520983 106997
rect 523200 106994 524400 107024
rect 520917 106992 524400 106994
rect 520917 106936 520922 106992
rect 520978 106936 524400 106992
rect 520917 106934 524400 106936
rect 520917 106931 520983 106934
rect 523200 106904 524400 106934
rect 110321 106314 110387 106317
rect 119110 106314 119170 106828
rect 110321 106312 119170 106314
rect 110321 106256 110326 106312
rect 110382 106256 119170 106312
rect 110321 106254 119170 106256
rect 110321 106251 110387 106254
rect 519629 105770 519695 105773
rect 518788 105768 519695 105770
rect 518788 105712 519634 105768
rect 519690 105712 519695 105768
rect 518788 105710 519695 105712
rect 519629 105707 519695 105710
rect 520273 105498 520339 105501
rect 523200 105498 524400 105528
rect 520273 105496 524400 105498
rect 520273 105440 520278 105496
rect 520334 105440 524400 105496
rect 520273 105438 524400 105440
rect 520273 105435 520339 105438
rect 523200 105408 524400 105438
rect 117129 104818 117195 104821
rect 117129 104816 119140 104818
rect 117129 104760 117134 104816
rect 117190 104760 119140 104816
rect 117129 104758 119140 104760
rect 117129 104755 117195 104758
rect 521101 104410 521167 104413
rect 518788 104408 521167 104410
rect 518788 104352 521106 104408
rect 521162 104352 521167 104408
rect 518788 104350 521167 104352
rect 521101 104347 521167 104350
rect 521193 104002 521259 104005
rect 523200 104002 524400 104032
rect 521193 104000 524400 104002
rect 521193 103944 521198 104000
rect 521254 103944 524400 104000
rect 521193 103942 524400 103944
rect 521193 103939 521259 103942
rect 523200 103912 524400 103942
rect 521561 103050 521627 103053
rect 518788 103048 521627 103050
rect 518788 102992 521566 103048
rect 521622 102992 521627 103048
rect 518788 102990 521627 102992
rect 521561 102987 521627 102990
rect 116945 102914 117011 102917
rect 116945 102912 119140 102914
rect 116945 102856 116950 102912
rect 117006 102856 119140 102912
rect 116945 102854 119140 102856
rect 116945 102851 117011 102854
rect 521101 102506 521167 102509
rect 523200 102506 524400 102536
rect 521101 102504 524400 102506
rect 521101 102448 521106 102504
rect 521162 102448 524400 102504
rect 521101 102446 524400 102448
rect 521101 102443 521167 102446
rect 523200 102416 524400 102446
rect 521285 101690 521351 101693
rect 518788 101688 521351 101690
rect 518788 101632 521290 101688
rect 521346 101632 521351 101688
rect 518788 101630 521351 101632
rect 521285 101627 521351 101630
rect 117037 101010 117103 101013
rect 521469 101010 521535 101013
rect 523200 101010 524400 101040
rect 117037 101008 119140 101010
rect 117037 100952 117042 101008
rect 117098 100952 119140 101008
rect 117037 100950 119140 100952
rect 521469 101008 524400 101010
rect 521469 100952 521474 101008
rect 521530 100952 524400 101008
rect 521469 100950 524400 100952
rect 117037 100947 117103 100950
rect 521469 100947 521535 100950
rect 523200 100920 524400 100950
rect 521009 100330 521075 100333
rect 518788 100328 521075 100330
rect 518788 100272 521014 100328
rect 521070 100272 521075 100328
rect 518788 100270 521075 100272
rect 521009 100267 521075 100270
rect 519813 99378 519879 99381
rect 523200 99378 524400 99408
rect 519813 99376 524400 99378
rect 519813 99320 519818 99376
rect 519874 99320 524400 99376
rect 519813 99318 524400 99320
rect 519813 99315 519879 99318
rect 523200 99288 524400 99318
rect 116853 99106 116919 99109
rect 116853 99104 119140 99106
rect 116853 99048 116858 99104
rect 116914 99048 119140 99104
rect 116853 99046 119140 99048
rect 116853 99043 116919 99046
rect 520917 98970 520983 98973
rect 518788 98968 520983 98970
rect 518788 98912 520922 98968
rect 520978 98912 520983 98968
rect 518788 98910 520983 98912
rect 520917 98907 520983 98910
rect 114093 98698 114159 98701
rect 110860 98696 114159 98698
rect 110860 98640 114098 98696
rect 114154 98640 114159 98696
rect 110860 98638 114159 98640
rect 114093 98635 114159 98638
rect 519721 97882 519787 97885
rect 523200 97882 524400 97912
rect 519721 97880 524400 97882
rect 519721 97824 519726 97880
rect 519782 97824 524400 97880
rect 519721 97822 524400 97824
rect 519721 97819 519787 97822
rect 523200 97792 524400 97822
rect 520273 97610 520339 97613
rect 518788 97608 520339 97610
rect 518788 97552 520278 97608
rect 520334 97552 520339 97608
rect 518788 97550 520339 97552
rect 520273 97547 520339 97550
rect 116761 97202 116827 97205
rect 116761 97200 119140 97202
rect 116761 97144 116766 97200
rect 116822 97144 119140 97200
rect 116761 97142 119140 97144
rect 116761 97139 116827 97142
rect 519261 96386 519327 96389
rect 523200 96386 524400 96416
rect 519261 96384 524400 96386
rect 519261 96328 519266 96384
rect 519322 96328 524400 96384
rect 519261 96326 524400 96328
rect 519261 96323 519327 96326
rect 523200 96296 524400 96326
rect 521193 96250 521259 96253
rect 518788 96248 521259 96250
rect 518788 96192 521198 96248
rect 521254 96192 521259 96248
rect 518788 96190 521259 96192
rect 521193 96187 521259 96190
rect 116669 95298 116735 95301
rect 116669 95296 119140 95298
rect 116669 95240 116674 95296
rect 116730 95240 119140 95296
rect 116669 95238 119140 95240
rect 116669 95235 116735 95238
rect 521101 95026 521167 95029
rect 518758 95024 521167 95026
rect 518758 94968 521106 95024
rect 521162 94968 521167 95024
rect 518758 94966 521167 94968
rect 518758 94860 518818 94966
rect 521101 94963 521167 94966
rect 519905 94890 519971 94893
rect 523200 94890 524400 94920
rect 519905 94888 524400 94890
rect 519905 94832 519910 94888
rect 519966 94832 524400 94888
rect 519905 94830 524400 94832
rect 519905 94827 519971 94830
rect 523200 94800 524400 94830
rect 521469 93530 521535 93533
rect 518788 93528 521535 93530
rect 518788 93472 521474 93528
rect 521530 93472 521535 93528
rect 518788 93470 521535 93472
rect 521469 93467 521535 93470
rect 116577 93394 116643 93397
rect 520181 93394 520247 93397
rect 523200 93394 524400 93424
rect 116577 93392 119140 93394
rect 116577 93336 116582 93392
rect 116638 93336 119140 93392
rect 116577 93334 119140 93336
rect 520181 93392 524400 93394
rect 520181 93336 520186 93392
rect 520242 93336 524400 93392
rect 520181 93334 524400 93336
rect 116577 93331 116643 93334
rect 520181 93331 520247 93334
rect 523200 93304 524400 93334
rect 519813 92170 519879 92173
rect 518788 92168 519879 92170
rect 518788 92112 519818 92168
rect 519874 92112 519879 92168
rect 518788 92110 519879 92112
rect 519813 92107 519879 92110
rect 521285 91898 521351 91901
rect 523200 91898 524400 91928
rect 521285 91896 524400 91898
rect 521285 91840 521290 91896
rect 521346 91840 524400 91896
rect 521285 91838 524400 91840
rect 521285 91835 521351 91838
rect 523200 91808 524400 91838
rect 116117 91354 116183 91357
rect 116117 91352 119140 91354
rect 116117 91296 116122 91352
rect 116178 91296 119140 91352
rect 116117 91294 119140 91296
rect 116117 91291 116183 91294
rect 519721 90810 519787 90813
rect 518788 90808 519787 90810
rect 518788 90752 519726 90808
rect 519782 90752 519787 90808
rect 518788 90750 519787 90752
rect 519721 90747 519787 90750
rect 520917 90266 520983 90269
rect 523200 90266 524400 90296
rect 520917 90264 524400 90266
rect 520917 90208 520922 90264
rect 520978 90208 524400 90264
rect 520917 90206 524400 90208
rect 520917 90203 520983 90206
rect 523200 90176 524400 90206
rect 116117 89450 116183 89453
rect 519261 89450 519327 89453
rect 116117 89448 119140 89450
rect 116117 89392 116122 89448
rect 116178 89392 119140 89448
rect 116117 89390 119140 89392
rect 518788 89448 519327 89450
rect 518788 89392 519266 89448
rect 519322 89392 519327 89448
rect 518788 89390 519327 89392
rect 116117 89387 116183 89390
rect 519261 89387 519327 89390
rect 521377 88770 521443 88773
rect 523200 88770 524400 88800
rect 521377 88768 524400 88770
rect 521377 88712 521382 88768
rect 521438 88712 524400 88768
rect 521377 88710 524400 88712
rect 521377 88707 521443 88710
rect 523200 88680 524400 88710
rect 519905 88090 519971 88093
rect 518788 88088 519971 88090
rect 518788 88032 519910 88088
rect 519966 88032 519971 88088
rect 518788 88030 519971 88032
rect 519905 88027 519971 88030
rect 116025 87546 116091 87549
rect 116025 87544 119140 87546
rect 116025 87488 116030 87544
rect 116086 87488 119140 87544
rect 116025 87486 119140 87488
rect 116025 87483 116091 87486
rect 114185 87274 114251 87277
rect 110860 87272 114251 87274
rect 110860 87216 114190 87272
rect 114246 87216 114251 87272
rect 110860 87214 114251 87216
rect 114185 87211 114251 87214
rect 521193 87274 521259 87277
rect 523200 87274 524400 87304
rect 521193 87272 524400 87274
rect 521193 87216 521198 87272
rect 521254 87216 524400 87272
rect 521193 87214 524400 87216
rect 521193 87211 521259 87214
rect 523200 87184 524400 87214
rect 520181 86730 520247 86733
rect 518788 86728 520247 86730
rect 518788 86672 520186 86728
rect 520242 86672 520247 86728
rect 518788 86670 520247 86672
rect 520181 86667 520247 86670
rect 520273 85778 520339 85781
rect 523200 85778 524400 85808
rect 520273 85776 524400 85778
rect 520273 85720 520278 85776
rect 520334 85720 524400 85776
rect 520273 85718 524400 85720
rect 520273 85715 520339 85718
rect 523200 85688 524400 85718
rect 115197 85642 115263 85645
rect 115197 85640 119140 85642
rect 115197 85584 115202 85640
rect 115258 85584 119140 85640
rect 115197 85582 119140 85584
rect 115197 85579 115263 85582
rect 521101 84282 521167 84285
rect 523200 84282 524400 84312
rect 521101 84280 524400 84282
rect 521101 84224 521106 84280
rect 521162 84224 524400 84280
rect 521101 84222 524400 84224
rect 521101 84219 521167 84222
rect 523200 84192 524400 84222
rect 521285 84010 521351 84013
rect 518788 84008 521351 84010
rect 518788 83952 521290 84008
rect 521346 83952 521351 84008
rect 518788 83950 521351 83952
rect 521285 83947 521351 83950
rect 116577 83738 116643 83741
rect 116577 83736 119140 83738
rect 116577 83680 116582 83736
rect 116638 83680 119140 83736
rect 116577 83678 119140 83680
rect 116577 83675 116643 83678
rect 520181 82786 520247 82789
rect 523200 82786 524400 82816
rect 520181 82784 524400 82786
rect 520181 82728 520186 82784
rect 520242 82728 524400 82784
rect 520181 82726 524400 82728
rect 520181 82723 520247 82726
rect 523200 82696 524400 82726
rect 520917 82650 520983 82653
rect 518788 82648 520983 82650
rect 518788 82592 520922 82648
rect 520978 82592 520983 82648
rect 518788 82590 520983 82592
rect 520917 82587 520983 82590
rect 116209 81834 116275 81837
rect 116209 81832 119140 81834
rect 116209 81776 116214 81832
rect 116270 81776 119140 81832
rect 116209 81774 119140 81776
rect 116209 81771 116275 81774
rect 521377 81290 521443 81293
rect 518788 81288 521443 81290
rect 518788 81232 521382 81288
rect 521438 81232 521443 81288
rect 518788 81230 521443 81232
rect 521377 81227 521443 81230
rect 519629 81154 519695 81157
rect 523200 81154 524400 81184
rect 519629 81152 524400 81154
rect 519629 81096 519634 81152
rect 519690 81096 524400 81152
rect 519629 81094 524400 81096
rect 519629 81091 519695 81094
rect 523200 81064 524400 81094
rect 115933 79930 115999 79933
rect 521193 79930 521259 79933
rect 115933 79928 119140 79930
rect 115933 79872 115938 79928
rect 115994 79872 119140 79928
rect 115933 79870 119140 79872
rect 518788 79928 521259 79930
rect 518788 79872 521198 79928
rect 521254 79872 521259 79928
rect 518788 79870 521259 79872
rect 115933 79867 115999 79870
rect 521193 79867 521259 79870
rect 519813 79658 519879 79661
rect 523200 79658 524400 79688
rect 519813 79656 524400 79658
rect 519813 79600 519818 79656
rect 519874 79600 524400 79656
rect 519813 79598 524400 79600
rect 519813 79595 519879 79598
rect 523200 79568 524400 79598
rect 520273 78570 520339 78573
rect 518788 78568 520339 78570
rect 518788 78512 520278 78568
rect 520334 78512 520339 78568
rect 518788 78510 520339 78512
rect 520273 78507 520339 78510
rect 519997 78162 520063 78165
rect 523200 78162 524400 78192
rect 519997 78160 524400 78162
rect 519997 78104 520002 78160
rect 520058 78104 524400 78160
rect 519997 78102 524400 78104
rect 519997 78099 520063 78102
rect 523200 78072 524400 78102
rect 116117 78026 116183 78029
rect 116117 78024 119140 78026
rect 116117 77968 116122 78024
rect 116178 77968 119140 78024
rect 116117 77966 119140 77968
rect 116117 77963 116183 77966
rect 521101 77210 521167 77213
rect 518788 77208 521167 77210
rect 518788 77152 521106 77208
rect 521162 77152 521167 77208
rect 518788 77150 521167 77152
rect 521101 77147 521167 77150
rect 519721 76666 519787 76669
rect 523200 76666 524400 76696
rect 519721 76664 524400 76666
rect 519721 76608 519726 76664
rect 519782 76608 524400 76664
rect 519721 76606 524400 76608
rect 519721 76603 519787 76606
rect 523200 76576 524400 76606
rect 520181 75986 520247 75989
rect 110860 75926 119140 75986
rect 518788 75984 520247 75986
rect 518788 75928 520186 75984
rect 520242 75928 520247 75984
rect 518788 75926 520247 75928
rect 520181 75923 520247 75926
rect 520089 75170 520155 75173
rect 523200 75170 524400 75200
rect 520089 75168 524400 75170
rect 520089 75112 520094 75168
rect 520150 75112 524400 75168
rect 520089 75110 524400 75112
rect 520089 75107 520155 75110
rect 523200 75080 524400 75110
rect 519629 74626 519695 74629
rect 518788 74624 519695 74626
rect 518788 74568 519634 74624
rect 519690 74568 519695 74624
rect 518788 74566 519695 74568
rect 519629 74563 519695 74566
rect 116669 74082 116735 74085
rect 116669 74080 119140 74082
rect 116669 74024 116674 74080
rect 116730 74024 119140 74080
rect 116669 74022 119140 74024
rect 116669 74019 116735 74022
rect 519629 73674 519695 73677
rect 523200 73674 524400 73704
rect 519629 73672 524400 73674
rect 519629 73616 519634 73672
rect 519690 73616 524400 73672
rect 519629 73614 524400 73616
rect 519629 73611 519695 73614
rect 523200 73584 524400 73614
rect 519813 73266 519879 73269
rect 518788 73264 519879 73266
rect 518788 73208 519818 73264
rect 519874 73208 519879 73264
rect 518788 73206 519879 73208
rect 519813 73203 519879 73206
rect 519997 72450 520063 72453
rect 518758 72448 520063 72450
rect 518758 72392 520002 72448
rect 520058 72392 520063 72448
rect 518758 72390 520063 72392
rect 116577 72178 116643 72181
rect 116577 72176 119140 72178
rect 116577 72120 116582 72176
rect 116638 72120 119140 72176
rect 116577 72118 119140 72120
rect 116577 72115 116643 72118
rect 518758 71876 518818 72390
rect 519997 72387 520063 72390
rect 520181 72042 520247 72045
rect 523200 72042 524400 72072
rect 520181 72040 524400 72042
rect 520181 71984 520186 72040
rect 520242 71984 524400 72040
rect 520181 71982 524400 71984
rect 520181 71979 520247 71982
rect 523200 71952 524400 71982
rect 519721 70546 519787 70549
rect 518788 70544 519787 70546
rect 518788 70488 519726 70544
rect 519782 70488 519787 70544
rect 518788 70486 519787 70488
rect 519721 70483 519787 70486
rect 519905 70546 519971 70549
rect 523200 70546 524400 70576
rect 519905 70544 524400 70546
rect 519905 70488 519910 70544
rect 519966 70488 524400 70544
rect 519905 70486 524400 70488
rect 519905 70483 519971 70486
rect 523200 70456 524400 70486
rect 116301 70274 116367 70277
rect 116301 70272 119140 70274
rect 116301 70216 116306 70272
rect 116362 70216 119140 70272
rect 116301 70214 119140 70216
rect 116301 70211 116367 70214
rect 520089 69186 520155 69189
rect 518788 69184 520155 69186
rect 518788 69128 520094 69184
rect 520150 69128 520155 69184
rect 518788 69126 520155 69128
rect 520089 69123 520155 69126
rect 519537 69050 519603 69053
rect 523200 69050 524400 69080
rect 519537 69048 524400 69050
rect 519537 68992 519542 69048
rect 519598 68992 524400 69048
rect 519537 68990 524400 68992
rect 519537 68987 519603 68990
rect 523200 68960 524400 68990
rect 116117 68370 116183 68373
rect 116117 68368 119140 68370
rect 116117 68312 116122 68368
rect 116178 68312 119140 68368
rect 116117 68310 119140 68312
rect 116117 68307 116183 68310
rect 519629 67826 519695 67829
rect 518788 67824 519695 67826
rect 518788 67768 519634 67824
rect 519690 67768 519695 67824
rect 518788 67766 519695 67768
rect 519629 67763 519695 67766
rect 519997 67554 520063 67557
rect 523200 67554 524400 67584
rect 519997 67552 524400 67554
rect 519997 67496 520002 67552
rect 520058 67496 524400 67552
rect 519997 67494 524400 67496
rect 519997 67491 520063 67494
rect 523200 67464 524400 67494
rect 116577 66466 116643 66469
rect 520181 66466 520247 66469
rect 116577 66464 119140 66466
rect 116577 66408 116582 66464
rect 116638 66408 119140 66464
rect 116577 66406 119140 66408
rect 518788 66464 520247 66466
rect 518788 66408 520186 66464
rect 520242 66408 520247 66464
rect 518788 66406 520247 66408
rect 116577 66403 116643 66406
rect 520181 66403 520247 66406
rect 519813 66058 519879 66061
rect 523200 66058 524400 66088
rect 519813 66056 524400 66058
rect 519813 66000 519818 66056
rect 519874 66000 524400 66056
rect 519813 65998 524400 66000
rect 519813 65995 519879 65998
rect 523200 65968 524400 65998
rect 519905 65106 519971 65109
rect 518788 65104 519971 65106
rect 518788 65048 519910 65104
rect 519966 65048 519971 65104
rect 518788 65046 519971 65048
rect 519905 65043 519971 65046
rect 113357 64562 113423 64565
rect 110860 64560 113423 64562
rect 110860 64504 113362 64560
rect 113418 64504 113423 64560
rect 110860 64502 113423 64504
rect 113357 64499 113423 64502
rect 116209 64562 116275 64565
rect 521101 64562 521167 64565
rect 523200 64562 524400 64592
rect 116209 64560 119140 64562
rect 116209 64504 116214 64560
rect 116270 64504 119140 64560
rect 116209 64502 119140 64504
rect 521101 64560 524400 64562
rect 521101 64504 521106 64560
rect 521162 64504 524400 64560
rect 521101 64502 524400 64504
rect 116209 64499 116275 64502
rect 521101 64499 521167 64502
rect 523200 64472 524400 64502
rect 519537 63746 519603 63749
rect 518788 63744 519603 63746
rect 518788 63688 519542 63744
rect 519598 63688 519603 63744
rect 518788 63686 519603 63688
rect 519537 63683 519603 63686
rect 520733 62930 520799 62933
rect 523200 62930 524400 62960
rect 520733 62928 524400 62930
rect 520733 62872 520738 62928
rect 520794 62872 524400 62928
rect 520733 62870 524400 62872
rect 520733 62867 520799 62870
rect 523200 62840 524400 62870
rect 116117 62658 116183 62661
rect 116117 62656 119140 62658
rect 116117 62600 116122 62656
rect 116178 62600 119140 62656
rect 116117 62598 119140 62600
rect 116117 62595 116183 62598
rect 521101 62386 521167 62389
rect 518788 62384 521167 62386
rect 518788 62328 521106 62384
rect 521162 62328 521167 62384
rect 518788 62326 521167 62328
rect 521101 62323 521167 62326
rect 520273 61434 520339 61437
rect 523200 61434 524400 61464
rect 520273 61432 524400 61434
rect 520273 61376 520278 61432
rect 520334 61376 524400 61432
rect 520273 61374 524400 61376
rect 520273 61371 520339 61374
rect 523200 61344 524400 61374
rect 519997 61026 520063 61029
rect 518788 61024 520063 61026
rect 518788 60968 520002 61024
rect 520058 60968 520063 61024
rect 518788 60966 520063 60968
rect 519997 60963 520063 60966
rect 116577 60618 116643 60621
rect 116577 60616 119140 60618
rect 116577 60560 116582 60616
rect 116638 60560 119140 60616
rect 116577 60558 119140 60560
rect 116577 60555 116643 60558
rect 521009 59938 521075 59941
rect 523200 59938 524400 59968
rect 521009 59936 524400 59938
rect 521009 59880 521014 59936
rect 521070 59880 524400 59936
rect 521009 59878 524400 59880
rect 521009 59875 521075 59878
rect 523200 59848 524400 59878
rect 519813 59666 519879 59669
rect 518788 59664 519879 59666
rect 518788 59608 519818 59664
rect 519874 59608 519879 59664
rect 518788 59606 519879 59608
rect 519813 59603 519879 59606
rect 110321 58034 110387 58037
rect 119110 58034 119170 58684
rect 521101 58442 521167 58445
rect 523200 58442 524400 58472
rect 521101 58440 524400 58442
rect 521101 58384 521106 58440
rect 521162 58384 524400 58440
rect 521101 58382 524400 58384
rect 521101 58379 521167 58382
rect 523200 58352 524400 58382
rect 520733 58306 520799 58309
rect 518788 58304 520799 58306
rect 518788 58248 520738 58304
rect 520794 58248 520799 58304
rect 518788 58246 520799 58248
rect 520733 58243 520799 58246
rect 110321 58032 119170 58034
rect 110321 57976 110326 58032
rect 110382 57976 119170 58032
rect 110321 57974 119170 57976
rect 110321 57971 110387 57974
rect 520181 56946 520247 56949
rect 518788 56944 520247 56946
rect 518788 56888 520186 56944
rect 520242 56888 520247 56944
rect 518788 56886 520247 56888
rect 520181 56883 520247 56886
rect 520365 56946 520431 56949
rect 523200 56946 524400 56976
rect 520365 56944 524400 56946
rect 520365 56888 520370 56944
rect 520426 56888 524400 56944
rect 520365 56886 524400 56888
rect 520365 56883 520431 56886
rect 523200 56856 524400 56886
rect 110321 56810 110387 56813
rect 110321 56808 119140 56810
rect 110321 56752 110326 56808
rect 110382 56752 119140 56808
rect 110321 56750 119140 56752
rect 110321 56747 110387 56750
rect 521009 55586 521075 55589
rect 518788 55584 521075 55586
rect 518788 55528 521014 55584
rect 521070 55528 521075 55584
rect 518788 55526 521075 55528
rect 521009 55523 521075 55526
rect 520273 55450 520339 55453
rect 523200 55450 524400 55480
rect 520273 55448 524400 55450
rect 520273 55392 520278 55448
rect 520334 55392 524400 55448
rect 520273 55390 524400 55392
rect 520273 55387 520339 55390
rect 523200 55360 524400 55390
rect 110321 53954 110387 53957
rect 119110 53954 119170 54876
rect 521101 54226 521167 54229
rect 518788 54224 521167 54226
rect 518788 54168 521106 54224
rect 521162 54168 521167 54224
rect 518788 54166 521167 54168
rect 521101 54163 521167 54166
rect 110321 53952 119170 53954
rect 110321 53896 110326 53952
rect 110382 53896 119170 53952
rect 110321 53894 119170 53896
rect 110321 53891 110387 53894
rect 519261 53818 519327 53821
rect 523200 53818 524400 53848
rect 519261 53816 524400 53818
rect 519261 53760 519266 53816
rect 519322 53760 524400 53816
rect 519261 53758 524400 53760
rect 519261 53755 519327 53758
rect 523200 53728 524400 53758
rect 114185 53138 114251 53141
rect 110860 53136 114251 53138
rect 110860 53080 114190 53136
rect 114246 53080 114251 53136
rect 110860 53078 114251 53080
rect 114185 53075 114251 53078
rect 110321 52594 110387 52597
rect 119110 52594 119170 52972
rect 520365 52866 520431 52869
rect 518788 52864 520431 52866
rect 518788 52808 520370 52864
rect 520426 52808 520431 52864
rect 518788 52806 520431 52808
rect 520365 52803 520431 52806
rect 110321 52592 119170 52594
rect 110321 52536 110326 52592
rect 110382 52536 119170 52592
rect 110321 52534 119170 52536
rect 110321 52531 110387 52534
rect 520089 52322 520155 52325
rect 523200 52322 524400 52352
rect 520089 52320 524400 52322
rect 520089 52264 520094 52320
rect 520150 52264 524400 52320
rect 520089 52262 524400 52264
rect 520089 52259 520155 52262
rect 523200 52232 524400 52262
rect 520273 51506 520339 51509
rect 518788 51504 520339 51506
rect 518788 51448 520278 51504
rect 520334 51448 520339 51504
rect 518788 51446 520339 51448
rect 520273 51443 520339 51446
rect 110321 51098 110387 51101
rect 110321 51096 119140 51098
rect 110321 51040 110326 51096
rect 110382 51040 119140 51096
rect 110321 51038 119140 51040
rect 110321 51035 110387 51038
rect 519997 50826 520063 50829
rect 523200 50826 524400 50856
rect 519997 50824 524400 50826
rect 519997 50768 520002 50824
rect 520058 50768 524400 50824
rect 519997 50766 524400 50768
rect 519997 50763 520063 50766
rect 523200 50736 524400 50766
rect 519261 50146 519327 50149
rect 518788 50144 519327 50146
rect 518788 50088 519266 50144
rect 519322 50088 519327 50144
rect 518788 50086 519327 50088
rect 519261 50083 519327 50086
rect 520181 49330 520247 49333
rect 523200 49330 524400 49360
rect 520181 49328 524400 49330
rect 520181 49272 520186 49328
rect 520242 49272 524400 49328
rect 520181 49270 524400 49272
rect 520181 49267 520247 49270
rect 523200 49240 524400 49270
rect 110321 48378 110387 48381
rect 119110 48378 119170 49164
rect 520089 48786 520155 48789
rect 518788 48784 520155 48786
rect 518788 48728 520094 48784
rect 520150 48728 520155 48784
rect 518788 48726 520155 48728
rect 520089 48723 520155 48726
rect 110321 48376 119170 48378
rect 110321 48320 110326 48376
rect 110382 48320 119170 48376
rect 110321 48318 119170 48320
rect 110321 48315 110387 48318
rect 519445 47834 519511 47837
rect 523200 47834 524400 47864
rect 519445 47832 524400 47834
rect 519445 47776 519450 47832
rect 519506 47776 524400 47832
rect 519445 47774 524400 47776
rect 519445 47771 519511 47774
rect 523200 47744 524400 47774
rect 519997 47426 520063 47429
rect 518788 47424 520063 47426
rect 518788 47368 520002 47424
rect 520058 47368 520063 47424
rect 518788 47366 520063 47368
rect 519997 47363 520063 47366
rect 110321 47154 110387 47157
rect 110321 47152 119140 47154
rect 110321 47096 110326 47152
rect 110382 47096 119140 47152
rect 110321 47094 119140 47096
rect 110321 47091 110387 47094
rect 519905 46338 519971 46341
rect 523200 46338 524400 46368
rect 519905 46336 524400 46338
rect 519905 46280 519910 46336
rect 519966 46280 524400 46336
rect 519905 46278 524400 46280
rect 519905 46275 519971 46278
rect 523200 46248 524400 46278
rect 520181 46066 520247 46069
rect 518788 46064 520247 46066
rect 518788 46008 520186 46064
rect 520242 46008 520247 46064
rect 518788 46006 520247 46008
rect 520181 46003 520247 46006
rect 110321 45114 110387 45117
rect 110873 45114 110939 45117
rect 110321 45112 110939 45114
rect 110321 45056 110326 45112
rect 110382 45056 110878 45112
rect 110934 45056 110939 45112
rect 110321 45054 110939 45056
rect 110321 45051 110387 45054
rect 110873 45051 110939 45054
rect 110321 44978 110387 44981
rect 110965 44978 111031 44981
rect 110321 44976 111031 44978
rect 110321 44920 110326 44976
rect 110382 44920 110970 44976
rect 111026 44920 111031 44976
rect 110321 44918 111031 44920
rect 110321 44915 110387 44918
rect 110965 44915 111031 44918
rect 111793 44298 111859 44301
rect 119110 44298 119170 45220
rect 519445 44706 519511 44709
rect 518788 44704 519511 44706
rect 518788 44648 519450 44704
rect 519506 44648 519511 44704
rect 518788 44646 519511 44648
rect 519445 44643 519511 44646
rect 519813 44706 519879 44709
rect 523200 44706 524400 44736
rect 519813 44704 524400 44706
rect 519813 44648 519818 44704
rect 519874 44648 524400 44704
rect 519813 44646 524400 44648
rect 519813 44643 519879 44646
rect 523200 44616 524400 44646
rect 111793 44296 119170 44298
rect 111793 44240 111798 44296
rect 111854 44240 119170 44296
rect 111793 44238 119170 44240
rect 111793 44235 111859 44238
rect 116117 43346 116183 43349
rect 519905 43346 519971 43349
rect 116117 43344 119140 43346
rect 116117 43288 116122 43344
rect 116178 43288 119140 43344
rect 116117 43286 119140 43288
rect 518788 43344 519971 43346
rect 518788 43288 519910 43344
rect 519966 43288 519971 43344
rect 518788 43286 519971 43288
rect 116117 43283 116183 43286
rect 519905 43283 519971 43286
rect 520181 43210 520247 43213
rect 523200 43210 524400 43240
rect 520181 43208 524400 43210
rect 520181 43152 520186 43208
rect 520242 43152 524400 43208
rect 520181 43150 524400 43152
rect 520181 43147 520247 43150
rect 523200 43120 524400 43150
rect 519813 41986 519879 41989
rect 518788 41984 519879 41986
rect 518788 41928 519818 41984
rect 519874 41928 519879 41984
rect 518788 41926 519879 41928
rect 519813 41923 519879 41926
rect 114093 41850 114159 41853
rect 110860 41848 114159 41850
rect 110860 41792 114098 41848
rect 114154 41792 114159 41848
rect 110860 41790 114159 41792
rect 114093 41787 114159 41790
rect 520089 41714 520155 41717
rect 523200 41714 524400 41744
rect 520089 41712 524400 41714
rect 520089 41656 520094 41712
rect 520150 41656 524400 41712
rect 520089 41654 524400 41656
rect 520089 41651 520155 41654
rect 523200 41624 524400 41654
rect 110413 41442 110479 41445
rect 110413 41440 119140 41442
rect 110413 41384 110418 41440
rect 110474 41384 119140 41440
rect 110413 41382 119140 41384
rect 110413 41379 110479 41382
rect 520181 40626 520247 40629
rect 518788 40624 520247 40626
rect 518788 40568 520186 40624
rect 520242 40568 520247 40624
rect 518788 40566 520247 40568
rect 520181 40563 520247 40566
rect 520181 40218 520247 40221
rect 523200 40218 524400 40248
rect 520181 40216 524400 40218
rect 520181 40160 520186 40216
rect 520242 40160 524400 40216
rect 520181 40158 524400 40160
rect 520181 40155 520247 40158
rect 523200 40128 524400 40158
rect 116761 39538 116827 39541
rect 116761 39536 119140 39538
rect 116761 39480 116766 39536
rect 116822 39480 119140 39536
rect 116761 39478 119140 39480
rect 116761 39475 116827 39478
rect 520089 39266 520155 39269
rect 518788 39264 520155 39266
rect 518788 39208 520094 39264
rect 520150 39208 520155 39264
rect 518788 39206 520155 39208
rect 520089 39203 520155 39206
rect 519813 38722 519879 38725
rect 523200 38722 524400 38752
rect 519813 38720 524400 38722
rect 519813 38664 519818 38720
rect 519874 38664 524400 38720
rect 519813 38662 524400 38664
rect 519813 38659 519879 38662
rect 523200 38632 524400 38662
rect 520181 37906 520247 37909
rect 518788 37904 520247 37906
rect 518788 37848 520186 37904
rect 520242 37848 520247 37904
rect 518788 37846 520247 37848
rect 520181 37843 520247 37846
rect 116669 37634 116735 37637
rect 116669 37632 119140 37634
rect 116669 37576 116674 37632
rect 116730 37576 119140 37632
rect 116669 37574 119140 37576
rect 116669 37571 116735 37574
rect 110321 37362 110387 37365
rect 110781 37362 110847 37365
rect 110321 37360 110847 37362
rect 110321 37304 110326 37360
rect 110382 37304 110786 37360
rect 110842 37304 110847 37360
rect 110321 37302 110847 37304
rect 110321 37299 110387 37302
rect 110781 37299 110847 37302
rect 521561 37226 521627 37229
rect 523200 37226 524400 37256
rect 521561 37224 524400 37226
rect 521561 37168 521566 37224
rect 521622 37168 524400 37224
rect 521561 37166 524400 37168
rect 521561 37163 521627 37166
rect 523200 37136 524400 37166
rect 519813 36546 519879 36549
rect 518788 36544 519879 36546
rect 518788 36488 519818 36544
rect 519874 36488 519879 36544
rect 518788 36486 519879 36488
rect 519813 36483 519879 36486
rect 521561 36002 521627 36005
rect 521561 36000 521670 36002
rect 521561 35944 521566 36000
rect 521622 35944 521670 36000
rect 521561 35939 521670 35944
rect 521610 35866 521670 35939
rect 518758 35806 521670 35866
rect 110321 35322 110387 35325
rect 111057 35322 111123 35325
rect 110321 35320 111123 35322
rect 110321 35264 110326 35320
rect 110382 35264 111062 35320
rect 111118 35264 111123 35320
rect 110321 35262 111123 35264
rect 110321 35259 110387 35262
rect 111057 35259 111123 35262
rect 110321 35186 110387 35189
rect 110321 35184 115950 35186
rect 110321 35128 110326 35184
rect 110382 35128 115950 35184
rect 110321 35126 115950 35128
rect 110321 35123 110387 35126
rect 115890 34642 115950 35126
rect 119110 34642 119170 35700
rect 518758 35156 518818 35806
rect 521101 35594 521167 35597
rect 523200 35594 524400 35624
rect 521101 35592 524400 35594
rect 521101 35536 521106 35592
rect 521162 35536 524400 35592
rect 521101 35534 524400 35536
rect 521101 35531 521167 35534
rect 523200 35504 524400 35534
rect 115890 34582 119170 34642
rect 521101 34506 521167 34509
rect 518758 34504 521167 34506
rect 518758 34448 521106 34504
rect 521162 34448 521167 34504
rect 518758 34446 521167 34448
rect 110321 33826 110387 33829
rect 111057 33826 111123 33829
rect 110321 33824 111123 33826
rect 110321 33768 110326 33824
rect 110382 33768 111062 33824
rect 111118 33768 111123 33824
rect 110321 33766 111123 33768
rect 110321 33763 110387 33766
rect 111057 33763 111123 33766
rect 116945 33826 117011 33829
rect 116945 33824 119140 33826
rect 116945 33768 116950 33824
rect 117006 33768 119140 33824
rect 518758 33796 518818 34446
rect 521101 34443 521167 34446
rect 520917 34098 520983 34101
rect 523200 34098 524400 34128
rect 520917 34096 524400 34098
rect 520917 34040 520922 34096
rect 520978 34040 524400 34096
rect 520917 34038 524400 34040
rect 520917 34035 520983 34038
rect 523200 34008 524400 34038
rect 116945 33766 119140 33768
rect 116945 33763 117011 33766
rect 520917 33146 520983 33149
rect 518758 33144 520983 33146
rect 518758 33088 520922 33144
rect 520978 33088 520983 33144
rect 518758 33086 520983 33088
rect 518758 32436 518818 33086
rect 520917 33083 520983 33086
rect 520917 32602 520983 32605
rect 523200 32602 524400 32632
rect 520917 32600 524400 32602
rect 520917 32544 520922 32600
rect 520978 32544 524400 32600
rect 520917 32542 524400 32544
rect 520917 32539 520983 32542
rect 523200 32512 524400 32542
rect 116853 31786 116919 31789
rect 116853 31784 119140 31786
rect 116853 31728 116858 31784
rect 116914 31728 119140 31784
rect 116853 31726 119140 31728
rect 116853 31723 116919 31726
rect 520917 31650 520983 31653
rect 518758 31648 520983 31650
rect 518758 31592 520922 31648
rect 520978 31592 520983 31648
rect 518758 31590 520983 31592
rect 518758 31076 518818 31590
rect 520917 31587 520983 31590
rect 520917 31106 520983 31109
rect 523200 31106 524400 31136
rect 520917 31104 524400 31106
rect 520917 31048 520922 31104
rect 520978 31048 524400 31104
rect 520917 31046 524400 31048
rect 520917 31043 520983 31046
rect 523200 31016 524400 31046
rect 114001 30426 114067 30429
rect 110860 30424 114067 30426
rect 110860 30368 114006 30424
rect 114062 30368 114067 30424
rect 110860 30366 114067 30368
rect 114001 30363 114067 30366
rect 520917 30290 520983 30293
rect 518758 30288 520983 30290
rect 518758 30232 520922 30288
rect 520978 30232 520983 30288
rect 518758 30230 520983 30232
rect 110597 29882 110663 29885
rect 111057 29882 111123 29885
rect 110597 29880 111123 29882
rect 110597 29824 110602 29880
rect 110658 29824 111062 29880
rect 111118 29824 111123 29880
rect 110597 29822 111123 29824
rect 110597 29819 110663 29822
rect 111057 29819 111123 29822
rect 117037 29882 117103 29885
rect 117037 29880 119140 29882
rect 117037 29824 117042 29880
rect 117098 29824 119140 29880
rect 117037 29822 119140 29824
rect 117037 29819 117103 29822
rect 110413 29746 110479 29749
rect 110781 29746 110847 29749
rect 110413 29744 110847 29746
rect 110413 29688 110418 29744
rect 110474 29688 110786 29744
rect 110842 29688 110847 29744
rect 518758 29716 518818 30230
rect 520917 30227 520983 30230
rect 110413 29686 110847 29688
rect 110413 29683 110479 29686
rect 110781 29683 110847 29686
rect 521101 29610 521167 29613
rect 523200 29610 524400 29640
rect 521101 29608 524400 29610
rect 521101 29552 521106 29608
rect 521162 29552 524400 29608
rect 521101 29550 524400 29552
rect 521101 29547 521167 29550
rect 523200 29520 524400 29550
rect 110505 28794 110571 28797
rect 111793 28794 111859 28797
rect 110505 28792 111859 28794
rect 110505 28736 110510 28792
rect 110566 28736 111798 28792
rect 111854 28736 111859 28792
rect 110505 28734 111859 28736
rect 110505 28731 110571 28734
rect 111793 28731 111859 28734
rect 110321 28658 110387 28661
rect 111057 28658 111123 28661
rect 110321 28656 111123 28658
rect 110321 28600 110326 28656
rect 110382 28600 111062 28656
rect 111118 28600 111123 28656
rect 110321 28598 111123 28600
rect 110321 28595 110387 28598
rect 111057 28595 111123 28598
rect 521101 28386 521167 28389
rect 518788 28384 521167 28386
rect 518788 28328 521106 28384
rect 521162 28328 521167 28384
rect 518788 28326 521167 28328
rect 521101 28323 521167 28326
rect 110321 28114 110387 28117
rect 110597 28114 110663 28117
rect 523200 28114 524400 28144
rect 110321 28112 110663 28114
rect 110321 28056 110326 28112
rect 110382 28056 110602 28112
rect 110658 28056 110663 28112
rect 110321 28054 110663 28056
rect 110321 28051 110387 28054
rect 110597 28051 110663 28054
rect 518850 28054 524400 28114
rect 117129 27978 117195 27981
rect 117129 27976 119140 27978
rect 117129 27920 117134 27976
rect 117190 27920 119140 27976
rect 117129 27918 119140 27920
rect 117129 27915 117195 27918
rect 110321 27706 110387 27709
rect 110965 27706 111031 27709
rect 110321 27704 111031 27706
rect 110321 27648 110326 27704
rect 110382 27648 110970 27704
rect 111026 27648 111031 27704
rect 110321 27646 111031 27648
rect 110321 27643 110387 27646
rect 110965 27643 111031 27646
rect 518850 27570 518910 28054
rect 523200 28024 524400 28054
rect 518758 27510 518910 27570
rect 110321 27162 110387 27165
rect 110873 27162 110939 27165
rect 110321 27160 110939 27162
rect 110321 27104 110326 27160
rect 110382 27104 110878 27160
rect 110934 27104 110939 27160
rect 110321 27102 110939 27104
rect 110321 27099 110387 27102
rect 110873 27099 110939 27102
rect 518758 26996 518818 27510
rect 523200 26482 524400 26512
rect 521610 26422 524400 26482
rect 521610 26210 521670 26422
rect 523200 26392 524400 26422
rect 518758 26150 521670 26210
rect 116393 26074 116459 26077
rect 116393 26072 119140 26074
rect 116393 26016 116398 26072
rect 116454 26016 119140 26072
rect 116393 26014 119140 26016
rect 116393 26011 116459 26014
rect 518758 25636 518818 26150
rect 523200 24986 524400 25016
rect 518850 24926 524400 24986
rect 518850 24850 518910 24926
rect 523200 24896 524400 24926
rect 518758 24790 518910 24850
rect 518758 24276 518818 24790
rect 117221 24170 117287 24173
rect 117221 24168 119140 24170
rect 117221 24112 117226 24168
rect 117282 24112 119140 24168
rect 117221 24110 119140 24112
rect 117221 24107 117287 24110
rect 523200 23490 524400 23520
rect 518758 23430 524400 23490
rect 518758 22916 518818 23430
rect 523200 23400 524400 23430
rect 116485 22266 116551 22269
rect 116485 22264 119140 22266
rect 116485 22208 116490 22264
rect 116546 22208 119140 22264
rect 116485 22206 119140 22208
rect 116485 22203 116551 22206
rect 521101 21994 521167 21997
rect 523200 21994 524400 22024
rect 521101 21992 524400 21994
rect 521101 21936 521106 21992
rect 521162 21936 524400 21992
rect 521101 21934 524400 21936
rect 521101 21931 521167 21934
rect 523200 21904 524400 21934
rect 518758 20906 518818 21556
rect 521101 20906 521167 20909
rect 518758 20904 521167 20906
rect 518758 20848 521106 20904
rect 521162 20848 521167 20904
rect 518758 20846 521167 20848
rect 521101 20843 521167 20846
rect 520733 20498 520799 20501
rect 523200 20498 524400 20528
rect 520733 20496 524400 20498
rect 520733 20440 520738 20496
rect 520794 20440 524400 20496
rect 520733 20438 524400 20440
rect 520733 20435 520799 20438
rect 523200 20408 524400 20438
rect 116301 20362 116367 20365
rect 116301 20360 119140 20362
rect 116301 20304 116306 20360
rect 116362 20304 119140 20360
rect 116301 20302 119140 20304
rect 116301 20299 116367 20302
rect 518758 19546 518818 20196
rect 520733 19546 520799 19549
rect 518758 19544 520799 19546
rect 518758 19488 520738 19544
rect 520794 19488 520799 19544
rect 518758 19486 520799 19488
rect 520733 19483 520799 19486
rect 113909 19002 113975 19005
rect 110860 19000 113975 19002
rect 110860 18944 113914 19000
rect 113970 18944 113975 19000
rect 110860 18942 113975 18944
rect 113909 18939 113975 18942
rect 520917 19002 520983 19005
rect 523200 19002 524400 19032
rect 520917 19000 524400 19002
rect 520917 18944 520922 19000
rect 520978 18944 524400 19000
rect 520917 18942 524400 18944
rect 520917 18939 520983 18942
rect 523200 18912 524400 18942
rect 116209 18458 116275 18461
rect 116209 18456 119140 18458
rect 116209 18400 116214 18456
rect 116270 18400 119140 18456
rect 116209 18398 119140 18400
rect 116209 18395 116275 18398
rect 518758 18186 518818 18836
rect 520917 18186 520983 18189
rect 518758 18184 520983 18186
rect 518758 18128 520922 18184
rect 520978 18128 520983 18184
rect 518758 18126 520983 18128
rect 520917 18123 520983 18126
rect 518758 16826 518818 17476
rect 523200 17370 524400 17400
rect 521150 17310 524400 17370
rect 521150 16826 521210 17310
rect 523200 17280 524400 17310
rect 518758 16766 521210 16826
rect 116025 16418 116091 16421
rect 116025 16416 119140 16418
rect 116025 16360 116030 16416
rect 116086 16360 119140 16416
rect 116025 16358 119140 16360
rect 116025 16355 116091 16358
rect 518758 15466 518818 16116
rect 523200 15874 524400 15904
rect 521104 15814 524400 15874
rect 521104 15466 521164 15814
rect 523200 15784 524400 15814
rect 518758 15406 521164 15466
rect 116117 14514 116183 14517
rect 116117 14512 119140 14514
rect 116117 14456 116122 14512
rect 116178 14456 119140 14512
rect 116117 14454 119140 14456
rect 116117 14451 116183 14454
rect 518758 14106 518818 14756
rect 523200 14378 524400 14408
rect 521104 14318 524400 14378
rect 521104 14106 521164 14318
rect 523200 14288 524400 14318
rect 518758 14046 521164 14106
rect 518758 12746 518818 13396
rect 523200 12882 524400 12912
rect 521104 12822 524400 12882
rect 521104 12746 521164 12822
rect 523200 12792 524400 12822
rect 518758 12686 521164 12746
rect 115933 12610 115999 12613
rect 115933 12608 119140 12610
rect 115933 12552 115938 12608
rect 115994 12552 119140 12608
rect 115933 12550 119140 12552
rect 115933 12547 115999 12550
rect 518758 11386 518818 12036
rect 523200 11386 524400 11416
rect 518758 11326 524400 11386
rect 523200 11296 524400 11326
rect 116526 10644 116532 10708
rect 116596 10706 116602 10708
rect 116596 10646 119140 10706
rect 116596 10644 116602 10646
rect 518758 10026 518818 10676
rect 518758 9966 518910 10026
rect 518850 9890 518910 9966
rect 523200 9890 524400 9920
rect 518850 9830 524400 9890
rect 523200 9800 524400 9830
rect 521101 9346 521167 9349
rect 518788 9344 521167 9346
rect 518788 9288 521106 9344
rect 521162 9288 521167 9344
rect 518788 9286 521167 9288
rect 521101 9283 521167 9286
rect 117262 8740 117268 8804
rect 117332 8802 117338 8804
rect 117332 8742 119140 8802
rect 117332 8740 117338 8742
rect 521101 8258 521167 8261
rect 523200 8258 524400 8288
rect 521101 8256 524400 8258
rect 521101 8200 521106 8256
rect 521162 8200 524400 8256
rect 521101 8198 524400 8200
rect 521101 8195 521167 8198
rect 523200 8168 524400 8198
rect 520365 7986 520431 7989
rect 518788 7984 520431 7986
rect 518788 7928 520370 7984
rect 520426 7928 520431 7984
rect 518788 7926 520431 7928
rect 520365 7923 520431 7926
rect 113817 7714 113883 7717
rect 110860 7712 113883 7714
rect 110860 7656 113822 7712
rect 113878 7656 113883 7712
rect 110860 7654 113883 7656
rect 113817 7651 113883 7654
rect 116158 6836 116164 6900
rect 116228 6898 116234 6900
rect 116228 6838 119140 6898
rect 116228 6836 116234 6838
rect 520365 6762 520431 6765
rect 523200 6762 524400 6792
rect 520365 6760 524400 6762
rect 520365 6704 520370 6760
rect 520426 6704 524400 6760
rect 520365 6702 524400 6704
rect 520365 6699 520431 6702
rect 523200 6672 524400 6702
rect 521101 6626 521167 6629
rect 518788 6624 521167 6626
rect 518788 6568 521106 6624
rect 521162 6568 521167 6624
rect 518788 6566 521167 6568
rect 521101 6563 521167 6566
rect 520917 5266 520983 5269
rect 518788 5264 520983 5266
rect 518788 5208 520922 5264
rect 520978 5208 520983 5264
rect 518788 5206 520983 5208
rect 520917 5203 520983 5206
rect 521101 5266 521167 5269
rect 523200 5266 524400 5296
rect 521101 5264 524400 5266
rect 521101 5208 521106 5264
rect 521162 5208 524400 5264
rect 521101 5206 524400 5208
rect 521101 5203 521167 5206
rect 523200 5176 524400 5206
rect 110689 4178 110755 4181
rect 119110 4178 119170 4964
rect 110689 4176 119170 4178
rect 110689 4120 110694 4176
rect 110750 4120 119170 4176
rect 110689 4118 119170 4120
rect 110689 4115 110755 4118
rect 63542 3982 91938 4042
rect 63542 3770 63602 3982
rect 59310 3710 63602 3770
rect 59310 3362 59370 3710
rect 42750 3302 46950 3362
rect 35850 3030 37290 3090
rect 35850 2818 35910 3030
rect 33182 2758 35910 2818
rect 33041 2682 33107 2685
rect 33182 2682 33242 2758
rect 33041 2680 33242 2682
rect 33041 2624 33046 2680
rect 33102 2624 33242 2680
rect 33041 2622 33242 2624
rect 37230 2682 37290 3030
rect 42750 2685 42810 3302
rect 46890 3226 46950 3302
rect 55170 3302 59370 3362
rect 69982 3438 91570 3498
rect 55170 3226 55230 3302
rect 46890 3166 55230 3226
rect 60690 3166 62130 3226
rect 60690 3090 60750 3166
rect 46890 3030 60750 3090
rect 42057 2682 42123 2685
rect 37230 2680 42123 2682
rect 37230 2624 42062 2680
rect 42118 2624 42123 2680
rect 37230 2622 42123 2624
rect 33041 2619 33107 2622
rect 42057 2619 42123 2622
rect 42701 2680 42810 2685
rect 42701 2624 42706 2680
rect 42762 2624 42810 2680
rect 42701 2622 42810 2624
rect 44725 2682 44791 2685
rect 46890 2682 46950 3030
rect 44725 2680 46950 2682
rect 44725 2624 44730 2680
rect 44786 2624 46950 2680
rect 44725 2622 46950 2624
rect 62070 2682 62130 3166
rect 69982 2954 70042 3438
rect 63036 2894 70042 2954
rect 73110 3302 74550 3362
rect 63036 2685 63096 2894
rect 73110 2818 73170 3302
rect 74490 2954 74550 3302
rect 82770 3302 86970 3362
rect 82770 2954 82830 3302
rect 74490 2894 82830 2954
rect 86910 2954 86970 3302
rect 86910 2894 90282 2954
rect 64094 2758 73170 2818
rect 74490 2758 90098 2818
rect 64094 2685 64154 2758
rect 62389 2682 62455 2685
rect 62070 2680 62455 2682
rect 62070 2624 62394 2680
rect 62450 2624 62455 2680
rect 62070 2622 62455 2624
rect 42701 2619 42767 2622
rect 44725 2619 44791 2622
rect 62389 2619 62455 2622
rect 63033 2680 63099 2685
rect 63033 2624 63038 2680
rect 63094 2624 63099 2680
rect 63033 2619 63099 2624
rect 64045 2680 64154 2685
rect 64045 2624 64050 2680
rect 64106 2624 64154 2680
rect 64045 2622 64154 2624
rect 68277 2682 68343 2685
rect 74490 2682 74550 2758
rect 90038 2685 90098 2758
rect 68277 2680 74550 2682
rect 68277 2624 68282 2680
rect 68338 2624 74550 2680
rect 68277 2622 74550 2624
rect 78765 2682 78831 2685
rect 87045 2682 87111 2685
rect 78765 2680 87111 2682
rect 78765 2624 78770 2680
rect 78826 2624 87050 2680
rect 87106 2624 87111 2680
rect 78765 2622 87111 2624
rect 90038 2680 90147 2685
rect 90038 2624 90086 2680
rect 90142 2624 90147 2680
rect 90038 2622 90147 2624
rect 90222 2682 90282 2894
rect 91510 2685 91570 3438
rect 91878 2685 91938 3982
rect 96570 3982 106290 4042
rect 96570 3770 96630 3982
rect 106230 3906 106290 3982
rect 110045 3906 110111 3909
rect 521009 3906 521075 3909
rect 93028 3710 96630 3770
rect 99330 3846 100770 3906
rect 93028 2685 93088 3710
rect 99330 3634 99390 3846
rect 100710 3770 100770 3846
rect 102090 3846 105738 3906
rect 106230 3904 110111 3906
rect 106230 3848 110050 3904
rect 110106 3848 110111 3904
rect 106230 3846 110111 3848
rect 518788 3904 521075 3906
rect 518788 3848 521014 3904
rect 521070 3848 521075 3904
rect 518788 3846 521075 3848
rect 102090 3770 102150 3846
rect 105678 3770 105738 3846
rect 110045 3843 110111 3846
rect 521009 3843 521075 3846
rect 110045 3770 110111 3773
rect 116945 3770 117011 3773
rect 100710 3710 102150 3770
rect 103470 3710 105554 3770
rect 105678 3710 106290 3770
rect 103470 3634 103530 3710
rect 96570 3574 99390 3634
rect 102090 3574 103530 3634
rect 96570 3226 96630 3574
rect 102090 3498 102150 3574
rect 97582 3438 102150 3498
rect 103240 3438 104496 3498
rect 97582 3226 97642 3438
rect 103240 3362 103300 3438
rect 93902 3166 96630 3226
rect 97398 3166 97642 3226
rect 102090 3302 103300 3362
rect 93902 2685 93962 3166
rect 97398 3090 97458 3166
rect 102090 3090 102150 3302
rect 95926 3030 97458 3090
rect 97766 3030 102150 3090
rect 104436 3090 104496 3438
rect 105494 3090 105554 3710
rect 106230 3362 106290 3710
rect 110045 3768 117011 3770
rect 110045 3712 110050 3768
rect 110106 3712 116950 3768
rect 117006 3712 117011 3768
rect 110045 3710 117011 3712
rect 110045 3707 110111 3710
rect 116945 3707 117011 3710
rect 520917 3770 520983 3773
rect 523200 3770 524400 3800
rect 520917 3768 524400 3770
rect 520917 3712 520922 3768
rect 520978 3712 524400 3768
rect 520917 3710 524400 3712
rect 520917 3707 520983 3710
rect 523200 3680 524400 3710
rect 109493 3634 109559 3637
rect 106782 3632 109559 3634
rect 106782 3576 109498 3632
rect 109554 3576 109559 3632
rect 106782 3574 109559 3576
rect 106782 3362 106842 3574
rect 109493 3571 109559 3574
rect 109401 3498 109467 3501
rect 117129 3498 117195 3501
rect 109401 3496 117195 3498
rect 109401 3440 109406 3496
rect 109462 3440 117134 3496
rect 117190 3440 117195 3496
rect 109401 3438 117195 3440
rect 109401 3435 109467 3438
rect 117129 3435 117195 3438
rect 106230 3302 106842 3362
rect 109493 3362 109559 3365
rect 116301 3362 116367 3365
rect 109493 3360 116367 3362
rect 109493 3304 109498 3360
rect 109554 3304 116306 3360
rect 116362 3304 116367 3360
rect 109493 3302 116367 3304
rect 109493 3299 109559 3302
rect 116301 3299 116367 3302
rect 110781 3226 110847 3229
rect 116761 3226 116827 3229
rect 110781 3224 116827 3226
rect 110781 3168 110786 3224
rect 110842 3168 116766 3224
rect 116822 3168 116827 3224
rect 110781 3166 116827 3168
rect 110781 3163 110847 3166
rect 116761 3163 116827 3166
rect 110045 3090 110111 3093
rect 104436 3030 104634 3090
rect 105494 3088 110111 3090
rect 105494 3032 110050 3088
rect 110106 3032 110111 3088
rect 105494 3030 110111 3032
rect 90357 2682 90423 2685
rect 90222 2680 90423 2682
rect 90222 2624 90362 2680
rect 90418 2624 90423 2680
rect 90222 2622 90423 2624
rect 91510 2680 91619 2685
rect 91510 2624 91558 2680
rect 91614 2624 91619 2680
rect 91510 2622 91619 2624
rect 91878 2680 91987 2685
rect 91878 2624 91926 2680
rect 91982 2624 91987 2680
rect 91878 2622 91987 2624
rect 64045 2619 64111 2622
rect 68277 2619 68343 2622
rect 78765 2619 78831 2622
rect 87045 2619 87111 2622
rect 90081 2619 90147 2622
rect 90357 2619 90423 2622
rect 91553 2619 91619 2622
rect 91921 2619 91987 2622
rect 93025 2680 93091 2685
rect 93025 2624 93030 2680
rect 93086 2624 93091 2680
rect 93025 2619 93091 2624
rect 93853 2680 93962 2685
rect 93853 2624 93858 2680
rect 93914 2624 93962 2680
rect 93853 2622 93962 2624
rect 95693 2682 95759 2685
rect 95926 2682 95986 3030
rect 97766 2685 97826 3030
rect 99054 2894 103898 2954
rect 95693 2680 95986 2682
rect 95693 2624 95698 2680
rect 95754 2624 95986 2680
rect 95693 2622 95986 2624
rect 97717 2680 97826 2685
rect 97717 2624 97722 2680
rect 97778 2624 97826 2680
rect 97717 2622 97826 2624
rect 97901 2682 97967 2685
rect 99054 2682 99114 2894
rect 103838 2818 103898 2894
rect 102090 2758 103530 2818
rect 103838 2758 104496 2818
rect 97901 2680 99114 2682
rect 97901 2624 97906 2680
rect 97962 2624 99114 2680
rect 97901 2622 99114 2624
rect 99189 2682 99255 2685
rect 102090 2682 102150 2758
rect 99189 2680 102150 2682
rect 99189 2624 99194 2680
rect 99250 2624 102150 2680
rect 99189 2622 102150 2624
rect 103470 2682 103530 2758
rect 104436 2685 104496 2758
rect 103697 2682 103763 2685
rect 103470 2680 103763 2682
rect 103470 2624 103702 2680
rect 103758 2624 103763 2680
rect 103470 2622 103763 2624
rect 93853 2619 93919 2622
rect 95693 2619 95759 2622
rect 97717 2619 97783 2622
rect 97901 2619 97967 2622
rect 99189 2619 99255 2622
rect 103697 2619 103763 2622
rect 104433 2680 104499 2685
rect 104433 2624 104438 2680
rect 104494 2624 104499 2680
rect 104433 2619 104499 2624
rect 104574 2682 104634 3030
rect 110045 3027 110111 3030
rect 116301 3090 116367 3093
rect 116301 3088 119140 3090
rect 116301 3032 116306 3088
rect 116362 3032 119140 3088
rect 116301 3030 119140 3032
rect 116301 3027 116367 3030
rect 109401 2954 109467 2957
rect 104850 2952 109467 2954
rect 104850 2896 109406 2952
rect 109462 2896 109467 2952
rect 104850 2894 109467 2896
rect 104850 2682 104910 2894
rect 109401 2891 109467 2894
rect 110321 2954 110387 2957
rect 110689 2954 110755 2957
rect 110321 2952 110755 2954
rect 110321 2896 110326 2952
rect 110382 2896 110694 2952
rect 110750 2896 110755 2952
rect 110321 2894 110755 2896
rect 110321 2891 110387 2894
rect 110689 2891 110755 2894
rect 104574 2622 104910 2682
rect 104985 2682 105051 2685
rect 106181 2682 106247 2685
rect 104985 2680 106247 2682
rect 104985 2624 104990 2680
rect 105046 2624 106186 2680
rect 106242 2624 106247 2680
rect 104985 2622 106247 2624
rect 104985 2619 105051 2622
rect 106181 2619 106247 2622
rect 106365 2682 106431 2685
rect 109861 2682 109927 2685
rect 521101 2682 521167 2685
rect 106365 2680 109927 2682
rect 106365 2624 106370 2680
rect 106426 2624 109866 2680
rect 109922 2624 109927 2680
rect 106365 2622 109927 2624
rect 518788 2680 521167 2682
rect 518788 2624 521106 2680
rect 521162 2624 521167 2680
rect 518788 2622 521167 2624
rect 106365 2619 106431 2622
rect 109861 2619 109927 2622
rect 521101 2619 521167 2622
rect 29545 2546 29611 2549
rect 116209 2546 116275 2549
rect 29545 2544 116275 2546
rect 29545 2488 29550 2544
rect 29606 2488 116214 2544
rect 116270 2488 116275 2544
rect 29545 2486 116275 2488
rect 29545 2483 29611 2486
rect 116209 2483 116275 2486
rect 26049 2410 26115 2413
rect 104433 2410 104499 2413
rect 26049 2408 104499 2410
rect 26049 2352 26054 2408
rect 26110 2352 104438 2408
rect 104494 2352 104499 2408
rect 26049 2350 104499 2352
rect 26049 2347 26115 2350
rect 104433 2347 104499 2350
rect 104617 2410 104683 2413
rect 116025 2410 116091 2413
rect 104617 2408 116091 2410
rect 104617 2352 104622 2408
rect 104678 2352 116030 2408
rect 116086 2352 116091 2408
rect 104617 2350 116091 2352
rect 104617 2347 104683 2350
rect 116025 2347 116091 2350
rect 22921 2274 22987 2277
rect 104433 2274 104499 2277
rect 22921 2272 104499 2274
rect 22921 2216 22926 2272
rect 22982 2216 104438 2272
rect 104494 2216 104499 2272
rect 22921 2214 104499 2216
rect 22921 2211 22987 2214
rect 104433 2211 104499 2214
rect 104617 2274 104683 2277
rect 116117 2274 116183 2277
rect 104617 2272 116183 2274
rect 104617 2216 104622 2272
rect 104678 2216 116122 2272
rect 116178 2216 116183 2272
rect 104617 2214 116183 2216
rect 104617 2211 104683 2214
rect 116117 2211 116183 2214
rect 521009 2274 521075 2277
rect 523200 2274 524400 2304
rect 521009 2272 524400 2274
rect 521009 2216 521014 2272
rect 521070 2216 524400 2272
rect 521009 2214 524400 2216
rect 521009 2211 521075 2214
rect 523200 2184 524400 2214
rect 19609 2138 19675 2141
rect 104341 2138 104407 2141
rect 19609 2136 104407 2138
rect 19609 2080 19614 2136
rect 19670 2080 104346 2136
rect 104402 2080 104407 2136
rect 19609 2078 104407 2080
rect 19609 2075 19675 2078
rect 104341 2075 104407 2078
rect 104617 2138 104683 2141
rect 115933 2138 115999 2141
rect 104617 2136 115999 2138
rect 104617 2080 104622 2136
rect 104678 2080 115938 2136
rect 115994 2080 115999 2136
rect 104617 2078 115999 2080
rect 104617 2075 104683 2078
rect 115933 2075 115999 2078
rect 16205 2002 16271 2005
rect 116526 2002 116532 2004
rect 16205 2000 116532 2002
rect 16205 1944 16210 2000
rect 16266 1944 116532 2000
rect 16205 1942 116532 1944
rect 16205 1939 16271 1942
rect 116526 1940 116532 1942
rect 116596 1940 116602 2004
rect 5993 1866 6059 1869
rect 110321 1866 110387 1869
rect 5993 1864 110387 1866
rect 5993 1808 5998 1864
rect 6054 1808 110326 1864
rect 110382 1808 110387 1864
rect 5993 1806 110387 1808
rect 5993 1803 6059 1806
rect 110321 1803 110387 1806
rect 12617 1730 12683 1733
rect 117262 1730 117268 1732
rect 12617 1728 117268 1730
rect 12617 1672 12622 1728
rect 12678 1672 117268 1728
rect 12617 1670 117268 1672
rect 12617 1667 12683 1670
rect 117262 1668 117268 1670
rect 117332 1668 117338 1732
rect 229277 1730 229343 1733
rect 293585 1730 293651 1733
rect 229277 1728 293651 1730
rect 229277 1672 229282 1728
rect 229338 1672 293590 1728
rect 293646 1672 293651 1728
rect 229277 1670 293651 1672
rect 229277 1667 229343 1670
rect 293585 1667 293651 1670
rect 9305 1594 9371 1597
rect 116158 1594 116164 1596
rect 9305 1592 116164 1594
rect 9305 1536 9310 1592
rect 9366 1536 116164 1592
rect 9305 1534 116164 1536
rect 9305 1531 9371 1534
rect 116158 1532 116164 1534
rect 116228 1532 116234 1596
rect 163773 1594 163839 1597
rect 243629 1594 243695 1597
rect 163773 1592 243695 1594
rect 163773 1536 163778 1592
rect 163834 1536 243634 1592
rect 243690 1536 243695 1592
rect 163773 1534 243695 1536
rect 163773 1531 163839 1534
rect 243629 1531 243695 1534
rect 55949 1458 56015 1461
rect 294781 1458 294847 1461
rect 55949 1456 294847 1458
rect 55949 1400 55954 1456
rect 56010 1400 294786 1456
rect 294842 1400 294847 1456
rect 55949 1398 294847 1400
rect 55949 1395 56015 1398
rect 294781 1395 294847 1398
rect 360285 1458 360351 1461
rect 393589 1458 393655 1461
rect 360285 1456 393655 1458
rect 360285 1400 360290 1456
rect 360346 1400 393594 1456
rect 393650 1400 393655 1456
rect 360285 1398 393655 1400
rect 360285 1395 360351 1398
rect 393589 1395 393655 1398
rect 87045 1322 87111 1325
rect 95693 1322 95759 1325
rect 87045 1320 95759 1322
rect 87045 1264 87050 1320
rect 87106 1264 95698 1320
rect 95754 1264 95759 1320
rect 87045 1262 95759 1264
rect 87045 1259 87111 1262
rect 95693 1259 95759 1262
rect 95969 1322 96035 1325
rect 97901 1322 97967 1325
rect 95969 1320 97967 1322
rect 95969 1264 95974 1320
rect 96030 1264 97906 1320
rect 97962 1264 97967 1320
rect 95969 1262 97967 1264
rect 95969 1259 96035 1262
rect 97901 1259 97967 1262
rect 98269 1322 98335 1325
rect 109861 1322 109927 1325
rect 98269 1320 109927 1322
rect 98269 1264 98274 1320
rect 98330 1264 109866 1320
rect 109922 1264 109927 1320
rect 98269 1262 109927 1264
rect 98269 1259 98335 1262
rect 109861 1259 109927 1262
rect 90357 1186 90423 1189
rect 97717 1186 97783 1189
rect 90357 1184 97783 1186
rect 90357 1128 90362 1184
rect 90418 1128 97722 1184
rect 97778 1128 97783 1184
rect 90357 1126 97783 1128
rect 90357 1123 90423 1126
rect 97717 1123 97783 1126
rect 99373 1186 99439 1189
rect 102593 1186 102659 1189
rect 99373 1184 102659 1186
rect 99373 1128 99378 1184
rect 99434 1128 102598 1184
rect 102654 1128 102659 1184
rect 99373 1126 102659 1128
rect 99373 1123 99439 1126
rect 102593 1123 102659 1126
rect 103697 1186 103763 1189
rect 109493 1186 109559 1189
rect 103697 1184 109559 1186
rect 103697 1128 103702 1184
rect 103758 1128 109498 1184
rect 109554 1128 109559 1184
rect 103697 1126 109559 1128
rect 103697 1123 103763 1126
rect 109493 1123 109559 1126
rect 90081 1050 90147 1053
rect 111057 1050 111123 1053
rect 90081 1048 111123 1050
rect 90081 992 90086 1048
rect 90142 992 111062 1048
rect 111118 992 111123 1048
rect 90081 990 111123 992
rect 90081 987 90147 990
rect 111057 987 111123 990
rect 521101 778 521167 781
rect 523200 778 524400 808
rect 521101 776 524400 778
rect 521101 720 521106 776
rect 521162 720 524400 776
rect 521101 718 524400 720
rect 521101 715 521167 718
rect 523200 688 524400 718
<< via3 >>
rect 116532 10644 116596 10708
rect 117268 8740 117332 8804
rect 116164 6836 116228 6900
rect 116532 1940 116596 2004
rect 117268 1668 117332 1732
rect 116164 1532 116228 1596
<< metal4 >>
rect 1664 144454 1984 144496
rect 1664 144218 1706 144454
rect 1942 144218 1984 144454
rect 1664 144134 1984 144218
rect 1664 143898 1706 144134
rect 1942 143898 1984 144134
rect 1664 143856 1984 143898
rect 109956 144454 110276 144496
rect 109956 144218 109998 144454
rect 110234 144218 110276 144454
rect 109956 144134 110276 144218
rect 109956 143898 109998 144134
rect 110234 143898 110276 144134
rect 109956 143856 110276 143898
rect 119664 144454 119984 144496
rect 119664 144218 119706 144454
rect 119942 144218 119984 144454
rect 119664 144134 119984 144218
rect 119664 143898 119706 144134
rect 119942 143898 119984 144134
rect 119664 143856 119984 143898
rect 517940 144454 518260 144496
rect 517940 144218 517982 144454
rect 518218 144218 518260 144454
rect 517940 144134 518260 144218
rect 517940 143898 517982 144134
rect 518218 143898 518260 144134
rect 517940 143856 518260 143898
rect 1096 131454 1332 131496
rect 1096 131134 1332 131218
rect 1096 130856 1332 130898
rect 110616 131454 110936 131496
rect 110616 131218 110658 131454
rect 110894 131218 110936 131454
rect 110616 131134 110936 131218
rect 110616 130898 110658 131134
rect 110894 130898 110936 131134
rect 110616 130856 110936 130898
rect 119004 131454 119324 131496
rect 119004 131218 119046 131454
rect 119282 131218 119324 131454
rect 119004 131134 119324 131218
rect 119004 130898 119046 131134
rect 119282 130898 119324 131134
rect 119004 130856 119324 130898
rect 518600 131454 518920 131496
rect 518600 131218 518642 131454
rect 518878 131218 518920 131454
rect 518600 131134 518920 131218
rect 518600 130898 518642 131134
rect 518878 130898 518920 131134
rect 518600 130856 518920 130898
rect 1664 118454 1984 118496
rect 1664 118218 1706 118454
rect 1942 118218 1984 118454
rect 1664 118134 1984 118218
rect 1664 117898 1706 118134
rect 1942 117898 1984 118134
rect 1664 117856 1984 117898
rect 109956 118454 110276 118496
rect 109956 118218 109998 118454
rect 110234 118218 110276 118454
rect 109956 118134 110276 118218
rect 109956 117898 109998 118134
rect 110234 117898 110276 118134
rect 109956 117856 110276 117898
rect 119664 118454 119984 118496
rect 119664 118218 119706 118454
rect 119942 118218 119984 118454
rect 119664 118134 119984 118218
rect 119664 117898 119706 118134
rect 119942 117898 119984 118134
rect 119664 117856 119984 117898
rect 517940 118454 518260 118496
rect 517940 118218 517982 118454
rect 518218 118218 518260 118454
rect 517940 118134 518260 118218
rect 517940 117898 517982 118134
rect 518218 117898 518260 118134
rect 517940 117856 518260 117898
rect 1096 105454 1332 105496
rect 1096 105134 1332 105218
rect 1096 104856 1332 104898
rect 110616 105454 110936 105496
rect 110616 105218 110658 105454
rect 110894 105218 110936 105454
rect 110616 105134 110936 105218
rect 110616 104898 110658 105134
rect 110894 104898 110936 105134
rect 110616 104856 110936 104898
rect 119004 105454 119324 105496
rect 119004 105218 119046 105454
rect 119282 105218 119324 105454
rect 119004 105134 119324 105218
rect 119004 104898 119046 105134
rect 119282 104898 119324 105134
rect 119004 104856 119324 104898
rect 518600 105454 518920 105496
rect 518600 105218 518642 105454
rect 518878 105218 518920 105454
rect 518600 105134 518920 105218
rect 518600 104898 518642 105134
rect 518878 104898 518920 105134
rect 518600 104856 518920 104898
rect 1664 92454 1984 92496
rect 1664 92218 1706 92454
rect 1942 92218 1984 92454
rect 1664 92134 1984 92218
rect 1664 91898 1706 92134
rect 1942 91898 1984 92134
rect 1664 91856 1984 91898
rect 109956 92454 110276 92496
rect 109956 92218 109998 92454
rect 110234 92218 110276 92454
rect 109956 92134 110276 92218
rect 109956 91898 109998 92134
rect 110234 91898 110276 92134
rect 109956 91856 110276 91898
rect 119664 92454 119984 92496
rect 119664 92218 119706 92454
rect 119942 92218 119984 92454
rect 119664 92134 119984 92218
rect 119664 91898 119706 92134
rect 119942 91898 119984 92134
rect 119664 91856 119984 91898
rect 517940 92454 518260 92496
rect 517940 92218 517982 92454
rect 518218 92218 518260 92454
rect 517940 92134 518260 92218
rect 517940 91898 517982 92134
rect 518218 91898 518260 92134
rect 517940 91856 518260 91898
rect 1096 79454 1332 79496
rect 1096 79134 1332 79218
rect 1096 78856 1332 78898
rect 110616 79454 110936 79496
rect 110616 79218 110658 79454
rect 110894 79218 110936 79454
rect 110616 79134 110936 79218
rect 110616 78898 110658 79134
rect 110894 78898 110936 79134
rect 110616 78856 110936 78898
rect 119004 79454 119324 79496
rect 119004 79218 119046 79454
rect 119282 79218 119324 79454
rect 119004 79134 119324 79218
rect 119004 78898 119046 79134
rect 119282 78898 119324 79134
rect 119004 78856 119324 78898
rect 518600 79454 518920 79496
rect 518600 79218 518642 79454
rect 518878 79218 518920 79454
rect 518600 79134 518920 79218
rect 518600 78898 518642 79134
rect 518878 78898 518920 79134
rect 518600 78856 518920 78898
rect 1664 66454 1984 66496
rect 1664 66218 1706 66454
rect 1942 66218 1984 66454
rect 1664 66134 1984 66218
rect 1664 65898 1706 66134
rect 1942 65898 1984 66134
rect 1664 65856 1984 65898
rect 109956 66454 110276 66496
rect 109956 66218 109998 66454
rect 110234 66218 110276 66454
rect 109956 66134 110276 66218
rect 109956 65898 109998 66134
rect 110234 65898 110276 66134
rect 109956 65856 110276 65898
rect 119664 66454 119984 66496
rect 119664 66218 119706 66454
rect 119942 66218 119984 66454
rect 119664 66134 119984 66218
rect 119664 65898 119706 66134
rect 119942 65898 119984 66134
rect 119664 65856 119984 65898
rect 517940 66454 518260 66496
rect 517940 66218 517982 66454
rect 518218 66218 518260 66454
rect 517940 66134 518260 66218
rect 517940 65898 517982 66134
rect 518218 65898 518260 66134
rect 517940 65856 518260 65898
rect 1096 53454 1332 53496
rect 1096 53134 1332 53218
rect 1096 52856 1332 52898
rect 110616 53454 110936 53496
rect 110616 53218 110658 53454
rect 110894 53218 110936 53454
rect 110616 53134 110936 53218
rect 110616 52898 110658 53134
rect 110894 52898 110936 53134
rect 110616 52856 110936 52898
rect 119004 53454 119324 53496
rect 119004 53218 119046 53454
rect 119282 53218 119324 53454
rect 119004 53134 119324 53218
rect 119004 52898 119046 53134
rect 119282 52898 119324 53134
rect 119004 52856 119324 52898
rect 518600 53454 518920 53496
rect 518600 53218 518642 53454
rect 518878 53218 518920 53454
rect 518600 53134 518920 53218
rect 518600 52898 518642 53134
rect 518878 52898 518920 53134
rect 518600 52856 518920 52898
rect 1664 40454 1984 40496
rect 1664 40218 1706 40454
rect 1942 40218 1984 40454
rect 1664 40134 1984 40218
rect 1664 39898 1706 40134
rect 1942 39898 1984 40134
rect 1664 39856 1984 39898
rect 109956 40454 110276 40496
rect 109956 40218 109998 40454
rect 110234 40218 110276 40454
rect 109956 40134 110276 40218
rect 109956 39898 109998 40134
rect 110234 39898 110276 40134
rect 109956 39856 110276 39898
rect 119664 40454 119984 40496
rect 119664 40218 119706 40454
rect 119942 40218 119984 40454
rect 119664 40134 119984 40218
rect 119664 39898 119706 40134
rect 119942 39898 119984 40134
rect 119664 39856 119984 39898
rect 517940 40454 518260 40496
rect 517940 40218 517982 40454
rect 518218 40218 518260 40454
rect 517940 40134 518260 40218
rect 517940 39898 517982 40134
rect 518218 39898 518260 40134
rect 517940 39856 518260 39898
rect 1096 27454 1332 27496
rect 1096 27134 1332 27218
rect 1096 26856 1332 26898
rect 110616 27454 110936 27496
rect 110616 27218 110658 27454
rect 110894 27218 110936 27454
rect 110616 27134 110936 27218
rect 110616 26898 110658 27134
rect 110894 26898 110936 27134
rect 110616 26856 110936 26898
rect 119004 27454 119324 27496
rect 119004 27218 119046 27454
rect 119282 27218 119324 27454
rect 119004 27134 119324 27218
rect 119004 26898 119046 27134
rect 119282 26898 119324 27134
rect 119004 26856 119324 26898
rect 518600 27454 518920 27496
rect 518600 27218 518642 27454
rect 518878 27218 518920 27454
rect 518600 27134 518920 27218
rect 518600 26898 518642 27134
rect 518878 26898 518920 27134
rect 518600 26856 518920 26898
rect 1664 14454 1984 14496
rect 1664 14218 1706 14454
rect 1942 14218 1984 14454
rect 1664 14134 1984 14218
rect 1664 13898 1706 14134
rect 1942 13898 1984 14134
rect 1664 13856 1984 13898
rect 109956 14454 110276 14496
rect 109956 14218 109998 14454
rect 110234 14218 110276 14454
rect 109956 14134 110276 14218
rect 109956 13898 109998 14134
rect 110234 13898 110276 14134
rect 109956 13856 110276 13898
rect 119664 14454 119984 14496
rect 119664 14218 119706 14454
rect 119942 14218 119984 14454
rect 119664 14134 119984 14218
rect 119664 13898 119706 14134
rect 119942 13898 119984 14134
rect 119664 13856 119984 13898
rect 517940 14454 518260 14496
rect 517940 14218 517982 14454
rect 518218 14218 518260 14454
rect 517940 14134 518260 14218
rect 517940 13898 517982 14134
rect 518218 13898 518260 14134
rect 517940 13856 518260 13898
rect 116531 10708 116597 10709
rect 116531 10644 116532 10708
rect 116596 10644 116597 10708
rect 116531 10643 116597 10644
rect 116163 6900 116229 6901
rect 116163 6836 116164 6900
rect 116228 6836 116229 6900
rect 116163 6835 116229 6836
rect 116166 1597 116226 6835
rect 116534 2005 116594 10643
rect 117267 8804 117333 8805
rect 117267 8740 117268 8804
rect 117332 8740 117333 8804
rect 117267 8739 117333 8740
rect 116531 2004 116597 2005
rect 116531 1940 116532 2004
rect 116596 1940 116597 2004
rect 116531 1939 116597 1940
rect 117270 1733 117330 8739
rect 117267 1732 117333 1733
rect 117267 1668 117268 1732
rect 117332 1668 117333 1732
rect 117267 1667 117333 1668
rect 116163 1596 116229 1597
rect 116163 1532 116164 1596
rect 116228 1532 116229 1596
rect 116163 1531 116229 1532
<< via4 >>
rect 1706 144218 1942 144454
rect 1706 143898 1942 144134
rect 109998 144218 110234 144454
rect 109998 143898 110234 144134
rect 119706 144218 119942 144454
rect 119706 143898 119942 144134
rect 517982 144218 518218 144454
rect 517982 143898 518218 144134
rect 1096 131218 1332 131454
rect 1096 130898 1332 131134
rect 110658 131218 110894 131454
rect 110658 130898 110894 131134
rect 119046 131218 119282 131454
rect 119046 130898 119282 131134
rect 518642 131218 518878 131454
rect 518642 130898 518878 131134
rect 1706 118218 1942 118454
rect 1706 117898 1942 118134
rect 109998 118218 110234 118454
rect 109998 117898 110234 118134
rect 119706 118218 119942 118454
rect 119706 117898 119942 118134
rect 517982 118218 518218 118454
rect 517982 117898 518218 118134
rect 1096 105218 1332 105454
rect 1096 104898 1332 105134
rect 110658 105218 110894 105454
rect 110658 104898 110894 105134
rect 119046 105218 119282 105454
rect 119046 104898 119282 105134
rect 518642 105218 518878 105454
rect 518642 104898 518878 105134
rect 1706 92218 1942 92454
rect 1706 91898 1942 92134
rect 109998 92218 110234 92454
rect 109998 91898 110234 92134
rect 119706 92218 119942 92454
rect 119706 91898 119942 92134
rect 517982 92218 518218 92454
rect 517982 91898 518218 92134
rect 1096 79218 1332 79454
rect 1096 78898 1332 79134
rect 110658 79218 110894 79454
rect 110658 78898 110894 79134
rect 119046 79218 119282 79454
rect 119046 78898 119282 79134
rect 518642 79218 518878 79454
rect 518642 78898 518878 79134
rect 1706 66218 1942 66454
rect 1706 65898 1942 66134
rect 109998 66218 110234 66454
rect 109998 65898 110234 66134
rect 119706 66218 119942 66454
rect 119706 65898 119942 66134
rect 517982 66218 518218 66454
rect 517982 65898 518218 66134
rect 1096 53218 1332 53454
rect 1096 52898 1332 53134
rect 110658 53218 110894 53454
rect 110658 52898 110894 53134
rect 119046 53218 119282 53454
rect 119046 52898 119282 53134
rect 518642 53218 518878 53454
rect 518642 52898 518878 53134
rect 1706 40218 1942 40454
rect 1706 39898 1942 40134
rect 109998 40218 110234 40454
rect 109998 39898 110234 40134
rect 119706 40218 119942 40454
rect 119706 39898 119942 40134
rect 517982 40218 518218 40454
rect 517982 39898 518218 40134
rect 1096 27218 1332 27454
rect 1096 26898 1332 27134
rect 110658 27218 110894 27454
rect 110658 26898 110894 27134
rect 119046 27218 119282 27454
rect 119046 26898 119282 27134
rect 518642 27218 518878 27454
rect 518642 26898 518878 27134
rect 1706 14218 1942 14454
rect 1706 13898 1942 14134
rect 109998 14218 110234 14454
rect 109998 13898 110234 14134
rect 119706 14218 119942 14454
rect 119706 13898 119942 14134
rect 517982 14218 518218 14454
rect 517982 13898 518218 14134
<< metal5 >>
rect 1104 156856 522836 157496
rect 1104 144454 2200 144496
rect 1104 144218 1706 144454
rect 1942 144218 2200 144454
rect 1104 144134 2200 144218
rect 1104 143898 1706 144134
rect 1942 143898 2200 144134
rect 1104 143856 2200 143898
rect 109800 144454 120200 144496
rect 109800 144218 109998 144454
rect 110234 144218 119706 144454
rect 119942 144218 120200 144454
rect 109800 144134 120200 144218
rect 109800 143898 109998 144134
rect 110234 143898 119706 144134
rect 119942 143898 120200 144134
rect 109800 143856 120200 143898
rect 517800 144454 522836 144496
rect 517800 144218 517982 144454
rect 518218 144218 522836 144454
rect 517800 144134 522836 144218
rect 517800 143898 517982 144134
rect 518218 143898 522836 144134
rect 517800 143856 522836 143898
rect 1072 131454 2200 131496
rect 1072 131218 1096 131454
rect 1332 131218 2200 131454
rect 1072 131134 2200 131218
rect 1072 130898 1096 131134
rect 1332 130898 2200 131134
rect 1072 130856 2200 130898
rect 109800 131454 120200 131496
rect 109800 131218 110658 131454
rect 110894 131218 119046 131454
rect 119282 131218 120200 131454
rect 109800 131134 120200 131218
rect 109800 130898 110658 131134
rect 110894 130898 119046 131134
rect 119282 130898 120200 131134
rect 109800 130856 120200 130898
rect 517800 131454 522836 131496
rect 517800 131218 518642 131454
rect 518878 131218 522836 131454
rect 517800 131134 522836 131218
rect 517800 130898 518642 131134
rect 518878 130898 522836 131134
rect 517800 130856 522836 130898
rect 1104 118454 2200 118496
rect 1104 118218 1706 118454
rect 1942 118218 2200 118454
rect 1104 118134 2200 118218
rect 1104 117898 1706 118134
rect 1942 117898 2200 118134
rect 1104 117856 2200 117898
rect 109800 118454 120200 118496
rect 109800 118218 109998 118454
rect 110234 118218 119706 118454
rect 119942 118218 120200 118454
rect 109800 118134 120200 118218
rect 109800 117898 109998 118134
rect 110234 117898 119706 118134
rect 119942 117898 120200 118134
rect 109800 117856 120200 117898
rect 517800 118454 522836 118496
rect 517800 118218 517982 118454
rect 518218 118218 522836 118454
rect 517800 118134 522836 118218
rect 517800 117898 517982 118134
rect 518218 117898 522836 118134
rect 517800 117856 522836 117898
rect 1072 105454 2200 105496
rect 1072 105218 1096 105454
rect 1332 105218 2200 105454
rect 1072 105134 2200 105218
rect 1072 104898 1096 105134
rect 1332 104898 2200 105134
rect 1072 104856 2200 104898
rect 109800 105454 120200 105496
rect 109800 105218 110658 105454
rect 110894 105218 119046 105454
rect 119282 105218 120200 105454
rect 109800 105134 120200 105218
rect 109800 104898 110658 105134
rect 110894 104898 119046 105134
rect 119282 104898 120200 105134
rect 109800 104856 120200 104898
rect 517800 105454 522836 105496
rect 517800 105218 518642 105454
rect 518878 105218 522836 105454
rect 517800 105134 522836 105218
rect 517800 104898 518642 105134
rect 518878 104898 522836 105134
rect 517800 104856 522836 104898
rect 1104 92454 2200 92496
rect 1104 92218 1706 92454
rect 1942 92218 2200 92454
rect 1104 92134 2200 92218
rect 1104 91898 1706 92134
rect 1942 91898 2200 92134
rect 1104 91856 2200 91898
rect 109800 92454 120200 92496
rect 109800 92218 109998 92454
rect 110234 92218 119706 92454
rect 119942 92218 120200 92454
rect 109800 92134 120200 92218
rect 109800 91898 109998 92134
rect 110234 91898 119706 92134
rect 119942 91898 120200 92134
rect 109800 91856 120200 91898
rect 517800 92454 522836 92496
rect 517800 92218 517982 92454
rect 518218 92218 522836 92454
rect 517800 92134 522836 92218
rect 517800 91898 517982 92134
rect 518218 91898 522836 92134
rect 517800 91856 522836 91898
rect 1072 79454 2200 79496
rect 1072 79218 1096 79454
rect 1332 79218 2200 79454
rect 1072 79134 2200 79218
rect 1072 78898 1096 79134
rect 1332 78898 2200 79134
rect 1072 78856 2200 78898
rect 109800 79454 120200 79496
rect 109800 79218 110658 79454
rect 110894 79218 119046 79454
rect 119282 79218 120200 79454
rect 109800 79134 120200 79218
rect 109800 78898 110658 79134
rect 110894 78898 119046 79134
rect 119282 78898 120200 79134
rect 109800 78856 120200 78898
rect 517800 79454 522836 79496
rect 517800 79218 518642 79454
rect 518878 79218 522836 79454
rect 517800 79134 522836 79218
rect 517800 78898 518642 79134
rect 518878 78898 522836 79134
rect 517800 78856 522836 78898
rect 1104 66454 2200 66496
rect 1104 66218 1706 66454
rect 1942 66218 2200 66454
rect 1104 66134 2200 66218
rect 1104 65898 1706 66134
rect 1942 65898 2200 66134
rect 1104 65856 2200 65898
rect 109800 66454 120200 66496
rect 109800 66218 109998 66454
rect 110234 66218 119706 66454
rect 119942 66218 120200 66454
rect 109800 66134 120200 66218
rect 109800 65898 109998 66134
rect 110234 65898 119706 66134
rect 119942 65898 120200 66134
rect 109800 65856 120200 65898
rect 517800 66454 522836 66496
rect 517800 66218 517982 66454
rect 518218 66218 522836 66454
rect 517800 66134 522836 66218
rect 517800 65898 517982 66134
rect 518218 65898 522836 66134
rect 517800 65856 522836 65898
rect 1072 53454 2200 53496
rect 1072 53218 1096 53454
rect 1332 53218 2200 53454
rect 1072 53134 2200 53218
rect 1072 52898 1096 53134
rect 1332 52898 2200 53134
rect 1072 52856 2200 52898
rect 109800 53454 120200 53496
rect 109800 53218 110658 53454
rect 110894 53218 119046 53454
rect 119282 53218 120200 53454
rect 109800 53134 120200 53218
rect 109800 52898 110658 53134
rect 110894 52898 119046 53134
rect 119282 52898 120200 53134
rect 109800 52856 120200 52898
rect 517800 53454 522836 53496
rect 517800 53218 518642 53454
rect 518878 53218 522836 53454
rect 517800 53134 522836 53218
rect 517800 52898 518642 53134
rect 518878 52898 522836 53134
rect 517800 52856 522836 52898
rect 1104 40454 2200 40496
rect 1104 40218 1706 40454
rect 1942 40218 2200 40454
rect 1104 40134 2200 40218
rect 1104 39898 1706 40134
rect 1942 39898 2200 40134
rect 1104 39856 2200 39898
rect 109800 40454 120200 40496
rect 109800 40218 109998 40454
rect 110234 40218 119706 40454
rect 119942 40218 120200 40454
rect 109800 40134 120200 40218
rect 109800 39898 109998 40134
rect 110234 39898 119706 40134
rect 119942 39898 120200 40134
rect 109800 39856 120200 39898
rect 517800 40454 522836 40496
rect 517800 40218 517982 40454
rect 518218 40218 522836 40454
rect 517800 40134 522836 40218
rect 517800 39898 517982 40134
rect 518218 39898 522836 40134
rect 517800 39856 522836 39898
rect 1072 27454 2200 27496
rect 1072 27218 1096 27454
rect 1332 27218 2200 27454
rect 1072 27134 2200 27218
rect 1072 26898 1096 27134
rect 1332 26898 2200 27134
rect 1072 26856 2200 26898
rect 109800 27454 120200 27496
rect 109800 27218 110658 27454
rect 110894 27218 119046 27454
rect 119282 27218 120200 27454
rect 109800 27134 120200 27218
rect 109800 26898 110658 27134
rect 110894 26898 119046 27134
rect 119282 26898 120200 27134
rect 109800 26856 120200 26898
rect 517800 27454 522836 27496
rect 517800 27218 518642 27454
rect 518878 27218 522836 27454
rect 517800 27134 522836 27218
rect 517800 26898 518642 27134
rect 518878 26898 522836 27134
rect 517800 26856 522836 26898
rect 1104 14454 2200 14496
rect 1104 14218 1706 14454
rect 1942 14218 2200 14454
rect 1104 14134 2200 14218
rect 1104 13898 1706 14134
rect 1942 13898 2200 14134
rect 1104 13856 2200 13898
rect 109800 14454 120200 14496
rect 109800 14218 109998 14454
rect 110234 14218 119706 14454
rect 119942 14218 120200 14454
rect 109800 14134 120200 14218
rect 109800 13898 109998 14134
rect 110234 13898 119706 14134
rect 119942 13898 120200 14134
rect 109800 13856 120200 13898
rect 517800 14454 522836 14496
rect 517800 14218 517982 14454
rect 518218 14218 522836 14454
rect 517800 14134 522836 14218
rect 517800 13898 517982 14134
rect 518218 13898 522836 14134
rect 517800 13856 522836 13898
use mgmt_core  core
timestamp 1638213420
transform 1 0 119000 0 1 2000
box 0 0 400000 148000
use DFFRAM  DFFRAM
timestamp 1638213420
transform 1 0 1000 0 1 2000
box 4 0 110000 148000
<< labels >>
rlabel metal5 s 1104 26856 2200 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 26856 120200 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 26856 522836 27496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 52856 2200 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 52856 120200 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 52856 522836 53496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 78856 2200 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 78856 120200 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 78856 522836 79496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 104856 2200 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 104856 120200 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 104856 522836 105496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 130856 2200 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 109800 130856 120200 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 517800 130856 522836 131496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 156856 522836 157496 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 13856 2200 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 13856 120200 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 13856 522836 14496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 39856 2200 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 39856 120200 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 39856 522836 40496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 65856 2200 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 65856 120200 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 65856 522836 66496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 91856 2200 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 91856 120200 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 91856 522836 92496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 117856 2200 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 117856 120200 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 117856 522836 118496 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 143856 2200 144496 6 VPWR
port 1 nsew power input
rlabel metal5 s 109800 143856 120200 144496 6 VPWR
port 1 nsew power input
rlabel metal5 s 517800 143856 522836 144496 6 VPWR
port 1 nsew power input
rlabel metal2 s 294786 -400 294842 800 6 core_clk
port 2 nsew signal input
rlabel metal2 s 98274 -400 98330 800 6 core_rstn
port 3 nsew signal input
rlabel metal3 s 523200 64472 524400 64592 6 debug_in
port 4 nsew signal input
rlabel metal3 s 523200 65968 524400 66088 6 debug_mode
port 5 nsew signal tristate
rlabel metal3 s 523200 67464 524400 67584 6 debug_oeb
port 6 nsew signal tristate
rlabel metal3 s 523200 68960 524400 69080 6 debug_out
port 7 nsew signal tristate
rlabel metal3 s 523200 144848 524400 144968 6 flash_clk
port 8 nsew signal tristate
rlabel metal3 s 523200 143352 524400 143472 6 flash_csb
port 9 nsew signal tristate
rlabel metal3 s 523200 146480 524400 146600 6 flash_io0_di
port 10 nsew signal input
rlabel metal3 s 523200 147976 524400 148096 6 flash_io0_do
port 11 nsew signal tristate
rlabel metal3 s 523200 149472 524400 149592 6 flash_io0_oeb
port 12 nsew signal tristate
rlabel metal3 s 523200 150968 524400 151088 6 flash_io1_di
port 13 nsew signal input
rlabel metal3 s 523200 152464 524400 152584 6 flash_io1_do
port 14 nsew signal tristate
rlabel metal3 s 523200 153960 524400 154080 6 flash_io1_oeb
port 15 nsew signal tristate
rlabel metal3 s 523200 155592 524400 155712 6 flash_io2_di
port 16 nsew signal input
rlabel metal3 s 523200 157088 524400 157208 6 flash_io2_do
port 17 nsew signal tristate
rlabel metal3 s 523200 158584 524400 158704 6 flash_io2_oeb
port 18 nsew signal tristate
rlabel metal3 s 523200 160080 524400 160200 6 flash_io3_di
port 19 nsew signal input
rlabel metal3 s 523200 161576 524400 161696 6 flash_io3_do
port 20 nsew signal tristate
rlabel metal3 s 523200 163072 524400 163192 6 flash_io3_oeb
port 21 nsew signal tristate
rlabel metal2 s 32770 -400 32826 800 6 gpio_in_pad
port 22 nsew signal input
rlabel metal2 s 163778 -400 163834 800 6 gpio_inenb_pad
port 23 nsew signal tristate
rlabel metal2 s 229282 -400 229338 800 6 gpio_mode0_pad
port 24 nsew signal tristate
rlabel metal2 s 360290 -400 360346 800 6 gpio_mode1_pad
port 25 nsew signal tristate
rlabel metal2 s 425794 -400 425850 800 6 gpio_out_pad
port 26 nsew signal tristate
rlabel metal2 s 491298 -400 491354 800 6 gpio_outenb_pad
port 27 nsew signal tristate
rlabel metal3 s 523200 91808 524400 91928 6 hk_ack_i
port 28 nsew signal input
rlabel metal3 s 523200 94800 524400 94920 6 hk_dat_i[0]
port 29 nsew signal input
rlabel metal3 s 523200 110032 524400 110152 6 hk_dat_i[10]
port 30 nsew signal input
rlabel metal3 s 523200 111528 524400 111648 6 hk_dat_i[11]
port 31 nsew signal input
rlabel metal3 s 523200 113024 524400 113144 6 hk_dat_i[12]
port 32 nsew signal input
rlabel metal3 s 523200 114520 524400 114640 6 hk_dat_i[13]
port 33 nsew signal input
rlabel metal3 s 523200 116016 524400 116136 6 hk_dat_i[14]
port 34 nsew signal input
rlabel metal3 s 523200 117512 524400 117632 6 hk_dat_i[15]
port 35 nsew signal input
rlabel metal3 s 523200 119144 524400 119264 6 hk_dat_i[16]
port 36 nsew signal input
rlabel metal3 s 523200 120640 524400 120760 6 hk_dat_i[17]
port 37 nsew signal input
rlabel metal3 s 523200 122136 524400 122256 6 hk_dat_i[18]
port 38 nsew signal input
rlabel metal3 s 523200 123632 524400 123752 6 hk_dat_i[19]
port 39 nsew signal input
rlabel metal3 s 523200 96296 524400 96416 6 hk_dat_i[1]
port 40 nsew signal input
rlabel metal3 s 523200 125128 524400 125248 6 hk_dat_i[20]
port 41 nsew signal input
rlabel metal3 s 523200 126624 524400 126744 6 hk_dat_i[21]
port 42 nsew signal input
rlabel metal3 s 523200 128256 524400 128376 6 hk_dat_i[22]
port 43 nsew signal input
rlabel metal3 s 523200 129752 524400 129872 6 hk_dat_i[23]
port 44 nsew signal input
rlabel metal3 s 523200 131248 524400 131368 6 hk_dat_i[24]
port 45 nsew signal input
rlabel metal3 s 523200 132744 524400 132864 6 hk_dat_i[25]
port 46 nsew signal input
rlabel metal3 s 523200 134240 524400 134360 6 hk_dat_i[26]
port 47 nsew signal input
rlabel metal3 s 523200 135736 524400 135856 6 hk_dat_i[27]
port 48 nsew signal input
rlabel metal3 s 523200 137368 524400 137488 6 hk_dat_i[28]
port 49 nsew signal input
rlabel metal3 s 523200 138864 524400 138984 6 hk_dat_i[29]
port 50 nsew signal input
rlabel metal3 s 523200 97792 524400 97912 6 hk_dat_i[2]
port 51 nsew signal input
rlabel metal3 s 523200 140360 524400 140480 6 hk_dat_i[30]
port 52 nsew signal input
rlabel metal3 s 523200 141856 524400 141976 6 hk_dat_i[31]
port 53 nsew signal input
rlabel metal3 s 523200 99288 524400 99408 6 hk_dat_i[3]
port 54 nsew signal input
rlabel metal3 s 523200 100920 524400 101040 6 hk_dat_i[4]
port 55 nsew signal input
rlabel metal3 s 523200 102416 524400 102536 6 hk_dat_i[5]
port 56 nsew signal input
rlabel metal3 s 523200 103912 524400 104032 6 hk_dat_i[6]
port 57 nsew signal input
rlabel metal3 s 523200 105408 524400 105528 6 hk_dat_i[7]
port 58 nsew signal input
rlabel metal3 s 523200 106904 524400 107024 6 hk_dat_i[8]
port 59 nsew signal input
rlabel metal3 s 523200 108400 524400 108520 6 hk_dat_i[9]
port 60 nsew signal input
rlabel metal3 s 523200 93304 524400 93424 6 hk_stb_o
port 61 nsew signal tristate
rlabel metal2 s 521842 163200 521898 164400 6 irq[0]
port 62 nsew signal input
rlabel metal2 s 522670 163200 522726 164400 6 irq[1]
port 63 nsew signal input
rlabel metal2 s 523498 163200 523554 164400 6 irq[2]
port 64 nsew signal input
rlabel metal3 s 523200 75080 524400 75200 6 irq[3]
port 65 nsew signal input
rlabel metal3 s 523200 73584 524400 73704 6 irq[4]
port 66 nsew signal input
rlabel metal3 s 523200 71952 524400 72072 6 irq[5]
port 67 nsew signal input
rlabel metal2 s 386 163200 442 164400 6 la_iena[0]
port 68 nsew signal tristate
rlabel metal2 s 336830 163200 336886 164400 6 la_iena[100]
port 69 nsew signal tristate
rlabel metal2 s 340142 163200 340198 164400 6 la_iena[101]
port 70 nsew signal tristate
rlabel metal2 s 343546 163200 343602 164400 6 la_iena[102]
port 71 nsew signal tristate
rlabel metal2 s 346858 163200 346914 164400 6 la_iena[103]
port 72 nsew signal tristate
rlabel metal2 s 350262 163200 350318 164400 6 la_iena[104]
port 73 nsew signal tristate
rlabel metal2 s 353666 163200 353722 164400 6 la_iena[105]
port 74 nsew signal tristate
rlabel metal2 s 356978 163200 357034 164400 6 la_iena[106]
port 75 nsew signal tristate
rlabel metal2 s 360382 163200 360438 164400 6 la_iena[107]
port 76 nsew signal tristate
rlabel metal2 s 363694 163200 363750 164400 6 la_iena[108]
port 77 nsew signal tristate
rlabel metal2 s 367098 163200 367154 164400 6 la_iena[109]
port 78 nsew signal tristate
rlabel metal2 s 33966 163200 34022 164400 6 la_iena[10]
port 79 nsew signal tristate
rlabel metal2 s 370410 163200 370466 164400 6 la_iena[110]
port 80 nsew signal tristate
rlabel metal2 s 373814 163200 373870 164400 6 la_iena[111]
port 81 nsew signal tristate
rlabel metal2 s 377218 163200 377274 164400 6 la_iena[112]
port 82 nsew signal tristate
rlabel metal2 s 380530 163200 380586 164400 6 la_iena[113]
port 83 nsew signal tristate
rlabel metal2 s 383934 163200 383990 164400 6 la_iena[114]
port 84 nsew signal tristate
rlabel metal2 s 387246 163200 387302 164400 6 la_iena[115]
port 85 nsew signal tristate
rlabel metal2 s 390650 163200 390706 164400 6 la_iena[116]
port 86 nsew signal tristate
rlabel metal2 s 393962 163200 394018 164400 6 la_iena[117]
port 87 nsew signal tristate
rlabel metal2 s 397366 163200 397422 164400 6 la_iena[118]
port 88 nsew signal tristate
rlabel metal2 s 400770 163200 400826 164400 6 la_iena[119]
port 89 nsew signal tristate
rlabel metal2 s 37370 163200 37426 164400 6 la_iena[11]
port 90 nsew signal tristate
rlabel metal2 s 404082 163200 404138 164400 6 la_iena[120]
port 91 nsew signal tristate
rlabel metal2 s 407486 163200 407542 164400 6 la_iena[121]
port 92 nsew signal tristate
rlabel metal2 s 410798 163200 410854 164400 6 la_iena[122]
port 93 nsew signal tristate
rlabel metal2 s 414202 163200 414258 164400 6 la_iena[123]
port 94 nsew signal tristate
rlabel metal2 s 417514 163200 417570 164400 6 la_iena[124]
port 95 nsew signal tristate
rlabel metal2 s 420918 163200 420974 164400 6 la_iena[125]
port 96 nsew signal tristate
rlabel metal2 s 424322 163200 424378 164400 6 la_iena[126]
port 97 nsew signal tristate
rlabel metal2 s 427634 163200 427690 164400 6 la_iena[127]
port 98 nsew signal tristate
rlabel metal2 s 40682 163200 40738 164400 6 la_iena[12]
port 99 nsew signal tristate
rlabel metal2 s 44086 163200 44142 164400 6 la_iena[13]
port 100 nsew signal tristate
rlabel metal2 s 47490 163200 47546 164400 6 la_iena[14]
port 101 nsew signal tristate
rlabel metal2 s 50802 163200 50858 164400 6 la_iena[15]
port 102 nsew signal tristate
rlabel metal2 s 54206 163200 54262 164400 6 la_iena[16]
port 103 nsew signal tristate
rlabel metal2 s 57518 163200 57574 164400 6 la_iena[17]
port 104 nsew signal tristate
rlabel metal2 s 60922 163200 60978 164400 6 la_iena[18]
port 105 nsew signal tristate
rlabel metal2 s 64234 163200 64290 164400 6 la_iena[19]
port 106 nsew signal tristate
rlabel metal2 s 3698 163200 3754 164400 6 la_iena[1]
port 107 nsew signal tristate
rlabel metal2 s 67638 163200 67694 164400 6 la_iena[20]
port 108 nsew signal tristate
rlabel metal2 s 71042 163200 71098 164400 6 la_iena[21]
port 109 nsew signal tristate
rlabel metal2 s 74354 163200 74410 164400 6 la_iena[22]
port 110 nsew signal tristate
rlabel metal2 s 77758 163200 77814 164400 6 la_iena[23]
port 111 nsew signal tristate
rlabel metal2 s 81070 163200 81126 164400 6 la_iena[24]
port 112 nsew signal tristate
rlabel metal2 s 84474 163200 84530 164400 6 la_iena[25]
port 113 nsew signal tristate
rlabel metal2 s 87786 163200 87842 164400 6 la_iena[26]
port 114 nsew signal tristate
rlabel metal2 s 91190 163200 91246 164400 6 la_iena[27]
port 115 nsew signal tristate
rlabel metal2 s 94594 163200 94650 164400 6 la_iena[28]
port 116 nsew signal tristate
rlabel metal2 s 97906 163200 97962 164400 6 la_iena[29]
port 117 nsew signal tristate
rlabel metal2 s 7102 163200 7158 164400 6 la_iena[2]
port 118 nsew signal tristate
rlabel metal2 s 101310 163200 101366 164400 6 la_iena[30]
port 119 nsew signal tristate
rlabel metal2 s 104622 163200 104678 164400 6 la_iena[31]
port 120 nsew signal tristate
rlabel metal2 s 108026 163200 108082 164400 6 la_iena[32]
port 121 nsew signal tristate
rlabel metal2 s 111338 163200 111394 164400 6 la_iena[33]
port 122 nsew signal tristate
rlabel metal2 s 114742 163200 114798 164400 6 la_iena[34]
port 123 nsew signal tristate
rlabel metal2 s 118146 163200 118202 164400 6 la_iena[35]
port 124 nsew signal tristate
rlabel metal2 s 121458 163200 121514 164400 6 la_iena[36]
port 125 nsew signal tristate
rlabel metal2 s 124862 163200 124918 164400 6 la_iena[37]
port 126 nsew signal tristate
rlabel metal2 s 128174 163200 128230 164400 6 la_iena[38]
port 127 nsew signal tristate
rlabel metal2 s 131578 163200 131634 164400 6 la_iena[39]
port 128 nsew signal tristate
rlabel metal2 s 10414 163200 10470 164400 6 la_iena[3]
port 129 nsew signal tristate
rlabel metal2 s 134890 163200 134946 164400 6 la_iena[40]
port 130 nsew signal tristate
rlabel metal2 s 138294 163200 138350 164400 6 la_iena[41]
port 131 nsew signal tristate
rlabel metal2 s 141698 163200 141754 164400 6 la_iena[42]
port 132 nsew signal tristate
rlabel metal2 s 145010 163200 145066 164400 6 la_iena[43]
port 133 nsew signal tristate
rlabel metal2 s 148414 163200 148470 164400 6 la_iena[44]
port 134 nsew signal tristate
rlabel metal2 s 151726 163200 151782 164400 6 la_iena[45]
port 135 nsew signal tristate
rlabel metal2 s 155130 163200 155186 164400 6 la_iena[46]
port 136 nsew signal tristate
rlabel metal2 s 158442 163200 158498 164400 6 la_iena[47]
port 137 nsew signal tristate
rlabel metal2 s 161846 163200 161902 164400 6 la_iena[48]
port 138 nsew signal tristate
rlabel metal2 s 165250 163200 165306 164400 6 la_iena[49]
port 139 nsew signal tristate
rlabel metal2 s 13818 163200 13874 164400 6 la_iena[4]
port 140 nsew signal tristate
rlabel metal2 s 168562 163200 168618 164400 6 la_iena[50]
port 141 nsew signal tristate
rlabel metal2 s 171966 163200 172022 164400 6 la_iena[51]
port 142 nsew signal tristate
rlabel metal2 s 175278 163200 175334 164400 6 la_iena[52]
port 143 nsew signal tristate
rlabel metal2 s 178682 163200 178738 164400 6 la_iena[53]
port 144 nsew signal tristate
rlabel metal2 s 181994 163200 182050 164400 6 la_iena[54]
port 145 nsew signal tristate
rlabel metal2 s 185398 163200 185454 164400 6 la_iena[55]
port 146 nsew signal tristate
rlabel metal2 s 188802 163200 188858 164400 6 la_iena[56]
port 147 nsew signal tristate
rlabel metal2 s 192114 163200 192170 164400 6 la_iena[57]
port 148 nsew signal tristate
rlabel metal2 s 195518 163200 195574 164400 6 la_iena[58]
port 149 nsew signal tristate
rlabel metal2 s 198830 163200 198886 164400 6 la_iena[59]
port 150 nsew signal tristate
rlabel metal2 s 17130 163200 17186 164400 6 la_iena[5]
port 151 nsew signal tristate
rlabel metal2 s 202234 163200 202290 164400 6 la_iena[60]
port 152 nsew signal tristate
rlabel metal2 s 205546 163200 205602 164400 6 la_iena[61]
port 153 nsew signal tristate
rlabel metal2 s 208950 163200 209006 164400 6 la_iena[62]
port 154 nsew signal tristate
rlabel metal2 s 212354 163200 212410 164400 6 la_iena[63]
port 155 nsew signal tristate
rlabel metal2 s 215666 163200 215722 164400 6 la_iena[64]
port 156 nsew signal tristate
rlabel metal2 s 219070 163200 219126 164400 6 la_iena[65]
port 157 nsew signal tristate
rlabel metal2 s 222382 163200 222438 164400 6 la_iena[66]
port 158 nsew signal tristate
rlabel metal2 s 225786 163200 225842 164400 6 la_iena[67]
port 159 nsew signal tristate
rlabel metal2 s 229098 163200 229154 164400 6 la_iena[68]
port 160 nsew signal tristate
rlabel metal2 s 232502 163200 232558 164400 6 la_iena[69]
port 161 nsew signal tristate
rlabel metal2 s 20534 163200 20590 164400 6 la_iena[6]
port 162 nsew signal tristate
rlabel metal2 s 235906 163200 235962 164400 6 la_iena[70]
port 163 nsew signal tristate
rlabel metal2 s 239218 163200 239274 164400 6 la_iena[71]
port 164 nsew signal tristate
rlabel metal2 s 242622 163200 242678 164400 6 la_iena[72]
port 165 nsew signal tristate
rlabel metal2 s 245934 163200 245990 164400 6 la_iena[73]
port 166 nsew signal tristate
rlabel metal2 s 249338 163200 249394 164400 6 la_iena[74]
port 167 nsew signal tristate
rlabel metal2 s 252650 163200 252706 164400 6 la_iena[75]
port 168 nsew signal tristate
rlabel metal2 s 256054 163200 256110 164400 6 la_iena[76]
port 169 nsew signal tristate
rlabel metal2 s 259458 163200 259514 164400 6 la_iena[77]
port 170 nsew signal tristate
rlabel metal2 s 262770 163200 262826 164400 6 la_iena[78]
port 171 nsew signal tristate
rlabel metal2 s 266174 163200 266230 164400 6 la_iena[79]
port 172 nsew signal tristate
rlabel metal2 s 23938 163200 23994 164400 6 la_iena[7]
port 173 nsew signal tristate
rlabel metal2 s 269486 163200 269542 164400 6 la_iena[80]
port 174 nsew signal tristate
rlabel metal2 s 272890 163200 272946 164400 6 la_iena[81]
port 175 nsew signal tristate
rlabel metal2 s 276202 163200 276258 164400 6 la_iena[82]
port 176 nsew signal tristate
rlabel metal2 s 279606 163200 279662 164400 6 la_iena[83]
port 177 nsew signal tristate
rlabel metal2 s 283010 163200 283066 164400 6 la_iena[84]
port 178 nsew signal tristate
rlabel metal2 s 286322 163200 286378 164400 6 la_iena[85]
port 179 nsew signal tristate
rlabel metal2 s 289726 163200 289782 164400 6 la_iena[86]
port 180 nsew signal tristate
rlabel metal2 s 293038 163200 293094 164400 6 la_iena[87]
port 181 nsew signal tristate
rlabel metal2 s 296442 163200 296498 164400 6 la_iena[88]
port 182 nsew signal tristate
rlabel metal2 s 299754 163200 299810 164400 6 la_iena[89]
port 183 nsew signal tristate
rlabel metal2 s 27250 163200 27306 164400 6 la_iena[8]
port 184 nsew signal tristate
rlabel metal2 s 303158 163200 303214 164400 6 la_iena[90]
port 185 nsew signal tristate
rlabel metal2 s 306562 163200 306618 164400 6 la_iena[91]
port 186 nsew signal tristate
rlabel metal2 s 309874 163200 309930 164400 6 la_iena[92]
port 187 nsew signal tristate
rlabel metal2 s 313278 163200 313334 164400 6 la_iena[93]
port 188 nsew signal tristate
rlabel metal2 s 316590 163200 316646 164400 6 la_iena[94]
port 189 nsew signal tristate
rlabel metal2 s 319994 163200 320050 164400 6 la_iena[95]
port 190 nsew signal tristate
rlabel metal2 s 323306 163200 323362 164400 6 la_iena[96]
port 191 nsew signal tristate
rlabel metal2 s 326710 163200 326766 164400 6 la_iena[97]
port 192 nsew signal tristate
rlabel metal2 s 330114 163200 330170 164400 6 la_iena[98]
port 193 nsew signal tristate
rlabel metal2 s 333426 163200 333482 164400 6 la_iena[99]
port 194 nsew signal tristate
rlabel metal2 s 30654 163200 30710 164400 6 la_iena[9]
port 195 nsew signal tristate
rlabel metal2 s 1214 163200 1270 164400 6 la_input[0]
port 196 nsew signal input
rlabel metal2 s 337658 163200 337714 164400 6 la_input[100]
port 197 nsew signal input
rlabel metal2 s 340970 163200 341026 164400 6 la_input[101]
port 198 nsew signal input
rlabel metal2 s 344374 163200 344430 164400 6 la_input[102]
port 199 nsew signal input
rlabel metal2 s 347778 163200 347834 164400 6 la_input[103]
port 200 nsew signal input
rlabel metal2 s 351090 163200 351146 164400 6 la_input[104]
port 201 nsew signal input
rlabel metal2 s 354494 163200 354550 164400 6 la_input[105]
port 202 nsew signal input
rlabel metal2 s 357806 163200 357862 164400 6 la_input[106]
port 203 nsew signal input
rlabel metal2 s 361210 163200 361266 164400 6 la_input[107]
port 204 nsew signal input
rlabel metal2 s 364522 163200 364578 164400 6 la_input[108]
port 205 nsew signal input
rlabel metal2 s 367926 163200 367982 164400 6 la_input[109]
port 206 nsew signal input
rlabel metal2 s 34794 163200 34850 164400 6 la_input[10]
port 207 nsew signal input
rlabel metal2 s 371330 163200 371386 164400 6 la_input[110]
port 208 nsew signal input
rlabel metal2 s 374642 163200 374698 164400 6 la_input[111]
port 209 nsew signal input
rlabel metal2 s 378046 163200 378102 164400 6 la_input[112]
port 210 nsew signal input
rlabel metal2 s 381358 163200 381414 164400 6 la_input[113]
port 211 nsew signal input
rlabel metal2 s 384762 163200 384818 164400 6 la_input[114]
port 212 nsew signal input
rlabel metal2 s 388074 163200 388130 164400 6 la_input[115]
port 213 nsew signal input
rlabel metal2 s 391478 163200 391534 164400 6 la_input[116]
port 214 nsew signal input
rlabel metal2 s 394882 163200 394938 164400 6 la_input[117]
port 215 nsew signal input
rlabel metal2 s 398194 163200 398250 164400 6 la_input[118]
port 216 nsew signal input
rlabel metal2 s 401598 163200 401654 164400 6 la_input[119]
port 217 nsew signal input
rlabel metal2 s 38198 163200 38254 164400 6 la_input[11]
port 218 nsew signal input
rlabel metal2 s 404910 163200 404966 164400 6 la_input[120]
port 219 nsew signal input
rlabel metal2 s 408314 163200 408370 164400 6 la_input[121]
port 220 nsew signal input
rlabel metal2 s 411626 163200 411682 164400 6 la_input[122]
port 221 nsew signal input
rlabel metal2 s 415030 163200 415086 164400 6 la_input[123]
port 222 nsew signal input
rlabel metal2 s 418434 163200 418490 164400 6 la_input[124]
port 223 nsew signal input
rlabel metal2 s 421746 163200 421802 164400 6 la_input[125]
port 224 nsew signal input
rlabel metal2 s 425150 163200 425206 164400 6 la_input[126]
port 225 nsew signal input
rlabel metal2 s 428462 163200 428518 164400 6 la_input[127]
port 226 nsew signal input
rlabel metal2 s 41602 163200 41658 164400 6 la_input[12]
port 227 nsew signal input
rlabel metal2 s 44914 163200 44970 164400 6 la_input[13]
port 228 nsew signal input
rlabel metal2 s 48318 163200 48374 164400 6 la_input[14]
port 229 nsew signal input
rlabel metal2 s 51630 163200 51686 164400 6 la_input[15]
port 230 nsew signal input
rlabel metal2 s 55034 163200 55090 164400 6 la_input[16]
port 231 nsew signal input
rlabel metal2 s 58346 163200 58402 164400 6 la_input[17]
port 232 nsew signal input
rlabel metal2 s 61750 163200 61806 164400 6 la_input[18]
port 233 nsew signal input
rlabel metal2 s 65154 163200 65210 164400 6 la_input[19]
port 234 nsew signal input
rlabel metal2 s 4526 163200 4582 164400 6 la_input[1]
port 235 nsew signal input
rlabel metal2 s 68466 163200 68522 164400 6 la_input[20]
port 236 nsew signal input
rlabel metal2 s 71870 163200 71926 164400 6 la_input[21]
port 237 nsew signal input
rlabel metal2 s 75182 163200 75238 164400 6 la_input[22]
port 238 nsew signal input
rlabel metal2 s 78586 163200 78642 164400 6 la_input[23]
port 239 nsew signal input
rlabel metal2 s 81898 163200 81954 164400 6 la_input[24]
port 240 nsew signal input
rlabel metal2 s 85302 163200 85358 164400 6 la_input[25]
port 241 nsew signal input
rlabel metal2 s 88706 163200 88762 164400 6 la_input[26]
port 242 nsew signal input
rlabel metal2 s 92018 163200 92074 164400 6 la_input[27]
port 243 nsew signal input
rlabel metal2 s 95422 163200 95478 164400 6 la_input[28]
port 244 nsew signal input
rlabel metal2 s 98734 163200 98790 164400 6 la_input[29]
port 245 nsew signal input
rlabel metal2 s 7930 163200 7986 164400 6 la_input[2]
port 246 nsew signal input
rlabel metal2 s 102138 163200 102194 164400 6 la_input[30]
port 247 nsew signal input
rlabel metal2 s 105450 163200 105506 164400 6 la_input[31]
port 248 nsew signal input
rlabel metal2 s 108854 163200 108910 164400 6 la_input[32]
port 249 nsew signal input
rlabel metal2 s 112258 163200 112314 164400 6 la_input[33]
port 250 nsew signal input
rlabel metal2 s 115570 163200 115626 164400 6 la_input[34]
port 251 nsew signal input
rlabel metal2 s 118974 163200 119030 164400 6 la_input[35]
port 252 nsew signal input
rlabel metal2 s 122286 163200 122342 164400 6 la_input[36]
port 253 nsew signal input
rlabel metal2 s 125690 163200 125746 164400 6 la_input[37]
port 254 nsew signal input
rlabel metal2 s 129002 163200 129058 164400 6 la_input[38]
port 255 nsew signal input
rlabel metal2 s 132406 163200 132462 164400 6 la_input[39]
port 256 nsew signal input
rlabel metal2 s 11242 163200 11298 164400 6 la_input[3]
port 257 nsew signal input
rlabel metal2 s 135810 163200 135866 164400 6 la_input[40]
port 258 nsew signal input
rlabel metal2 s 139122 163200 139178 164400 6 la_input[41]
port 259 nsew signal input
rlabel metal2 s 142526 163200 142582 164400 6 la_input[42]
port 260 nsew signal input
rlabel metal2 s 145838 163200 145894 164400 6 la_input[43]
port 261 nsew signal input
rlabel metal2 s 149242 163200 149298 164400 6 la_input[44]
port 262 nsew signal input
rlabel metal2 s 152554 163200 152610 164400 6 la_input[45]
port 263 nsew signal input
rlabel metal2 s 155958 163200 156014 164400 6 la_input[46]
port 264 nsew signal input
rlabel metal2 s 159362 163200 159418 164400 6 la_input[47]
port 265 nsew signal input
rlabel metal2 s 162674 163200 162730 164400 6 la_input[48]
port 266 nsew signal input
rlabel metal2 s 166078 163200 166134 164400 6 la_input[49]
port 267 nsew signal input
rlabel metal2 s 14646 163200 14702 164400 6 la_input[4]
port 268 nsew signal input
rlabel metal2 s 169390 163200 169446 164400 6 la_input[50]
port 269 nsew signal input
rlabel metal2 s 172794 163200 172850 164400 6 la_input[51]
port 270 nsew signal input
rlabel metal2 s 176106 163200 176162 164400 6 la_input[52]
port 271 nsew signal input
rlabel metal2 s 179510 163200 179566 164400 6 la_input[53]
port 272 nsew signal input
rlabel metal2 s 182914 163200 182970 164400 6 la_input[54]
port 273 nsew signal input
rlabel metal2 s 186226 163200 186282 164400 6 la_input[55]
port 274 nsew signal input
rlabel metal2 s 189630 163200 189686 164400 6 la_input[56]
port 275 nsew signal input
rlabel metal2 s 192942 163200 192998 164400 6 la_input[57]
port 276 nsew signal input
rlabel metal2 s 196346 163200 196402 164400 6 la_input[58]
port 277 nsew signal input
rlabel metal2 s 199658 163200 199714 164400 6 la_input[59]
port 278 nsew signal input
rlabel metal2 s 18050 163200 18106 164400 6 la_input[5]
port 279 nsew signal input
rlabel metal2 s 203062 163200 203118 164400 6 la_input[60]
port 280 nsew signal input
rlabel metal2 s 206466 163200 206522 164400 6 la_input[61]
port 281 nsew signal input
rlabel metal2 s 209778 163200 209834 164400 6 la_input[62]
port 282 nsew signal input
rlabel metal2 s 213182 163200 213238 164400 6 la_input[63]
port 283 nsew signal input
rlabel metal2 s 216494 163200 216550 164400 6 la_input[64]
port 284 nsew signal input
rlabel metal2 s 219898 163200 219954 164400 6 la_input[65]
port 285 nsew signal input
rlabel metal2 s 223210 163200 223266 164400 6 la_input[66]
port 286 nsew signal input
rlabel metal2 s 226614 163200 226670 164400 6 la_input[67]
port 287 nsew signal input
rlabel metal2 s 230018 163200 230074 164400 6 la_input[68]
port 288 nsew signal input
rlabel metal2 s 233330 163200 233386 164400 6 la_input[69]
port 289 nsew signal input
rlabel metal2 s 21362 163200 21418 164400 6 la_input[6]
port 290 nsew signal input
rlabel metal2 s 236734 163200 236790 164400 6 la_input[70]
port 291 nsew signal input
rlabel metal2 s 240046 163200 240102 164400 6 la_input[71]
port 292 nsew signal input
rlabel metal2 s 243450 163200 243506 164400 6 la_input[72]
port 293 nsew signal input
rlabel metal2 s 246762 163200 246818 164400 6 la_input[73]
port 294 nsew signal input
rlabel metal2 s 250166 163200 250222 164400 6 la_input[74]
port 295 nsew signal input
rlabel metal2 s 253570 163200 253626 164400 6 la_input[75]
port 296 nsew signal input
rlabel metal2 s 256882 163200 256938 164400 6 la_input[76]
port 297 nsew signal input
rlabel metal2 s 260286 163200 260342 164400 6 la_input[77]
port 298 nsew signal input
rlabel metal2 s 263598 163200 263654 164400 6 la_input[78]
port 299 nsew signal input
rlabel metal2 s 267002 163200 267058 164400 6 la_input[79]
port 300 nsew signal input
rlabel metal2 s 24766 163200 24822 164400 6 la_input[7]
port 301 nsew signal input
rlabel metal2 s 270314 163200 270370 164400 6 la_input[80]
port 302 nsew signal input
rlabel metal2 s 273718 163200 273774 164400 6 la_input[81]
port 303 nsew signal input
rlabel metal2 s 277122 163200 277178 164400 6 la_input[82]
port 304 nsew signal input
rlabel metal2 s 280434 163200 280490 164400 6 la_input[83]
port 305 nsew signal input
rlabel metal2 s 283838 163200 283894 164400 6 la_input[84]
port 306 nsew signal input
rlabel metal2 s 287150 163200 287206 164400 6 la_input[85]
port 307 nsew signal input
rlabel metal2 s 290554 163200 290610 164400 6 la_input[86]
port 308 nsew signal input
rlabel metal2 s 293866 163200 293922 164400 6 la_input[87]
port 309 nsew signal input
rlabel metal2 s 297270 163200 297326 164400 6 la_input[88]
port 310 nsew signal input
rlabel metal2 s 300674 163200 300730 164400 6 la_input[89]
port 311 nsew signal input
rlabel metal2 s 28078 163200 28134 164400 6 la_input[8]
port 312 nsew signal input
rlabel metal2 s 303986 163200 304042 164400 6 la_input[90]
port 313 nsew signal input
rlabel metal2 s 307390 163200 307446 164400 6 la_input[91]
port 314 nsew signal input
rlabel metal2 s 310702 163200 310758 164400 6 la_input[92]
port 315 nsew signal input
rlabel metal2 s 314106 163200 314162 164400 6 la_input[93]
port 316 nsew signal input
rlabel metal2 s 317418 163200 317474 164400 6 la_input[94]
port 317 nsew signal input
rlabel metal2 s 320822 163200 320878 164400 6 la_input[95]
port 318 nsew signal input
rlabel metal2 s 324226 163200 324282 164400 6 la_input[96]
port 319 nsew signal input
rlabel metal2 s 327538 163200 327594 164400 6 la_input[97]
port 320 nsew signal input
rlabel metal2 s 330942 163200 330998 164400 6 la_input[98]
port 321 nsew signal input
rlabel metal2 s 334254 163200 334310 164400 6 la_input[99]
port 322 nsew signal input
rlabel metal2 s 31482 163200 31538 164400 6 la_input[9]
port 323 nsew signal input
rlabel metal2 s 2042 163200 2098 164400 6 la_oenb[0]
port 324 nsew signal tristate
rlabel metal2 s 338486 163200 338542 164400 6 la_oenb[100]
port 325 nsew signal tristate
rlabel metal2 s 341890 163200 341946 164400 6 la_oenb[101]
port 326 nsew signal tristate
rlabel metal2 s 345202 163200 345258 164400 6 la_oenb[102]
port 327 nsew signal tristate
rlabel metal2 s 348606 163200 348662 164400 6 la_oenb[103]
port 328 nsew signal tristate
rlabel metal2 s 351918 163200 351974 164400 6 la_oenb[104]
port 329 nsew signal tristate
rlabel metal2 s 355322 163200 355378 164400 6 la_oenb[105]
port 330 nsew signal tristate
rlabel metal2 s 358634 163200 358690 164400 6 la_oenb[106]
port 331 nsew signal tristate
rlabel metal2 s 362038 163200 362094 164400 6 la_oenb[107]
port 332 nsew signal tristate
rlabel metal2 s 365442 163200 365498 164400 6 la_oenb[108]
port 333 nsew signal tristate
rlabel metal2 s 368754 163200 368810 164400 6 la_oenb[109]
port 334 nsew signal tristate
rlabel metal2 s 35714 163200 35770 164400 6 la_oenb[10]
port 335 nsew signal tristate
rlabel metal2 s 372158 163200 372214 164400 6 la_oenb[110]
port 336 nsew signal tristate
rlabel metal2 s 375470 163200 375526 164400 6 la_oenb[111]
port 337 nsew signal tristate
rlabel metal2 s 378874 163200 378930 164400 6 la_oenb[112]
port 338 nsew signal tristate
rlabel metal2 s 382186 163200 382242 164400 6 la_oenb[113]
port 339 nsew signal tristate
rlabel metal2 s 385590 163200 385646 164400 6 la_oenb[114]
port 340 nsew signal tristate
rlabel metal2 s 388994 163200 389050 164400 6 la_oenb[115]
port 341 nsew signal tristate
rlabel metal2 s 392306 163200 392362 164400 6 la_oenb[116]
port 342 nsew signal tristate
rlabel metal2 s 395710 163200 395766 164400 6 la_oenb[117]
port 343 nsew signal tristate
rlabel metal2 s 399022 163200 399078 164400 6 la_oenb[118]
port 344 nsew signal tristate
rlabel metal2 s 402426 163200 402482 164400 6 la_oenb[119]
port 345 nsew signal tristate
rlabel metal2 s 39026 163200 39082 164400 6 la_oenb[11]
port 346 nsew signal tristate
rlabel metal2 s 405738 163200 405794 164400 6 la_oenb[120]
port 347 nsew signal tristate
rlabel metal2 s 409142 163200 409198 164400 6 la_oenb[121]
port 348 nsew signal tristate
rlabel metal2 s 412546 163200 412602 164400 6 la_oenb[122]
port 349 nsew signal tristate
rlabel metal2 s 415858 163200 415914 164400 6 la_oenb[123]
port 350 nsew signal tristate
rlabel metal2 s 419262 163200 419318 164400 6 la_oenb[124]
port 351 nsew signal tristate
rlabel metal2 s 422574 163200 422630 164400 6 la_oenb[125]
port 352 nsew signal tristate
rlabel metal2 s 425978 163200 426034 164400 6 la_oenb[126]
port 353 nsew signal tristate
rlabel metal2 s 429290 163200 429346 164400 6 la_oenb[127]
port 354 nsew signal tristate
rlabel metal2 s 42430 163200 42486 164400 6 la_oenb[12]
port 355 nsew signal tristate
rlabel metal2 s 45742 163200 45798 164400 6 la_oenb[13]
port 356 nsew signal tristate
rlabel metal2 s 49146 163200 49202 164400 6 la_oenb[14]
port 357 nsew signal tristate
rlabel metal2 s 52458 163200 52514 164400 6 la_oenb[15]
port 358 nsew signal tristate
rlabel metal2 s 55862 163200 55918 164400 6 la_oenb[16]
port 359 nsew signal tristate
rlabel metal2 s 59266 163200 59322 164400 6 la_oenb[17]
port 360 nsew signal tristate
rlabel metal2 s 62578 163200 62634 164400 6 la_oenb[18]
port 361 nsew signal tristate
rlabel metal2 s 65982 163200 66038 164400 6 la_oenb[19]
port 362 nsew signal tristate
rlabel metal2 s 5354 163200 5410 164400 6 la_oenb[1]
port 363 nsew signal tristate
rlabel metal2 s 69294 163200 69350 164400 6 la_oenb[20]
port 364 nsew signal tristate
rlabel metal2 s 72698 163200 72754 164400 6 la_oenb[21]
port 365 nsew signal tristate
rlabel metal2 s 76010 163200 76066 164400 6 la_oenb[22]
port 366 nsew signal tristate
rlabel metal2 s 79414 163200 79470 164400 6 la_oenb[23]
port 367 nsew signal tristate
rlabel metal2 s 82818 163200 82874 164400 6 la_oenb[24]
port 368 nsew signal tristate
rlabel metal2 s 86130 163200 86186 164400 6 la_oenb[25]
port 369 nsew signal tristate
rlabel metal2 s 89534 163200 89590 164400 6 la_oenb[26]
port 370 nsew signal tristate
rlabel metal2 s 92846 163200 92902 164400 6 la_oenb[27]
port 371 nsew signal tristate
rlabel metal2 s 96250 163200 96306 164400 6 la_oenb[28]
port 372 nsew signal tristate
rlabel metal2 s 99562 163200 99618 164400 6 la_oenb[29]
port 373 nsew signal tristate
rlabel metal2 s 8758 163200 8814 164400 6 la_oenb[2]
port 374 nsew signal tristate
rlabel metal2 s 102966 163200 103022 164400 6 la_oenb[30]
port 375 nsew signal tristate
rlabel metal2 s 106370 163200 106426 164400 6 la_oenb[31]
port 376 nsew signal tristate
rlabel metal2 s 109682 163200 109738 164400 6 la_oenb[32]
port 377 nsew signal tristate
rlabel metal2 s 113086 163200 113142 164400 6 la_oenb[33]
port 378 nsew signal tristate
rlabel metal2 s 116398 163200 116454 164400 6 la_oenb[34]
port 379 nsew signal tristate
rlabel metal2 s 119802 163200 119858 164400 6 la_oenb[35]
port 380 nsew signal tristate
rlabel metal2 s 123114 163200 123170 164400 6 la_oenb[36]
port 381 nsew signal tristate
rlabel metal2 s 126518 163200 126574 164400 6 la_oenb[37]
port 382 nsew signal tristate
rlabel metal2 s 129922 163200 129978 164400 6 la_oenb[38]
port 383 nsew signal tristate
rlabel metal2 s 133234 163200 133290 164400 6 la_oenb[39]
port 384 nsew signal tristate
rlabel metal2 s 12162 163200 12218 164400 6 la_oenb[3]
port 385 nsew signal tristate
rlabel metal2 s 136638 163200 136694 164400 6 la_oenb[40]
port 386 nsew signal tristate
rlabel metal2 s 139950 163200 140006 164400 6 la_oenb[41]
port 387 nsew signal tristate
rlabel metal2 s 143354 163200 143410 164400 6 la_oenb[42]
port 388 nsew signal tristate
rlabel metal2 s 146666 163200 146722 164400 6 la_oenb[43]
port 389 nsew signal tristate
rlabel metal2 s 150070 163200 150126 164400 6 la_oenb[44]
port 390 nsew signal tristate
rlabel metal2 s 153474 163200 153530 164400 6 la_oenb[45]
port 391 nsew signal tristate
rlabel metal2 s 156786 163200 156842 164400 6 la_oenb[46]
port 392 nsew signal tristate
rlabel metal2 s 160190 163200 160246 164400 6 la_oenb[47]
port 393 nsew signal tristate
rlabel metal2 s 163502 163200 163558 164400 6 la_oenb[48]
port 394 nsew signal tristate
rlabel metal2 s 166906 163200 166962 164400 6 la_oenb[49]
port 395 nsew signal tristate
rlabel metal2 s 15474 163200 15530 164400 6 la_oenb[4]
port 396 nsew signal tristate
rlabel metal2 s 170218 163200 170274 164400 6 la_oenb[50]
port 397 nsew signal tristate
rlabel metal2 s 173622 163200 173678 164400 6 la_oenb[51]
port 398 nsew signal tristate
rlabel metal2 s 177026 163200 177082 164400 6 la_oenb[52]
port 399 nsew signal tristate
rlabel metal2 s 180338 163200 180394 164400 6 la_oenb[53]
port 400 nsew signal tristate
rlabel metal2 s 183742 163200 183798 164400 6 la_oenb[54]
port 401 nsew signal tristate
rlabel metal2 s 187054 163200 187110 164400 6 la_oenb[55]
port 402 nsew signal tristate
rlabel metal2 s 190458 163200 190514 164400 6 la_oenb[56]
port 403 nsew signal tristate
rlabel metal2 s 193770 163200 193826 164400 6 la_oenb[57]
port 404 nsew signal tristate
rlabel metal2 s 197174 163200 197230 164400 6 la_oenb[58]
port 405 nsew signal tristate
rlabel metal2 s 200578 163200 200634 164400 6 la_oenb[59]
port 406 nsew signal tristate
rlabel metal2 s 18878 163200 18934 164400 6 la_oenb[5]
port 407 nsew signal tristate
rlabel metal2 s 203890 163200 203946 164400 6 la_oenb[60]
port 408 nsew signal tristate
rlabel metal2 s 207294 163200 207350 164400 6 la_oenb[61]
port 409 nsew signal tristate
rlabel metal2 s 210606 163200 210662 164400 6 la_oenb[62]
port 410 nsew signal tristate
rlabel metal2 s 214010 163200 214066 164400 6 la_oenb[63]
port 411 nsew signal tristate
rlabel metal2 s 217322 163200 217378 164400 6 la_oenb[64]
port 412 nsew signal tristate
rlabel metal2 s 220726 163200 220782 164400 6 la_oenb[65]
port 413 nsew signal tristate
rlabel metal2 s 224130 163200 224186 164400 6 la_oenb[66]
port 414 nsew signal tristate
rlabel metal2 s 227442 163200 227498 164400 6 la_oenb[67]
port 415 nsew signal tristate
rlabel metal2 s 230846 163200 230902 164400 6 la_oenb[68]
port 416 nsew signal tristate
rlabel metal2 s 234158 163200 234214 164400 6 la_oenb[69]
port 417 nsew signal tristate
rlabel metal2 s 22190 163200 22246 164400 6 la_oenb[6]
port 418 nsew signal tristate
rlabel metal2 s 237562 163200 237618 164400 6 la_oenb[70]
port 419 nsew signal tristate
rlabel metal2 s 240874 163200 240930 164400 6 la_oenb[71]
port 420 nsew signal tristate
rlabel metal2 s 244278 163200 244334 164400 6 la_oenb[72]
port 421 nsew signal tristate
rlabel metal2 s 247682 163200 247738 164400 6 la_oenb[73]
port 422 nsew signal tristate
rlabel metal2 s 250994 163200 251050 164400 6 la_oenb[74]
port 423 nsew signal tristate
rlabel metal2 s 254398 163200 254454 164400 6 la_oenb[75]
port 424 nsew signal tristate
rlabel metal2 s 257710 163200 257766 164400 6 la_oenb[76]
port 425 nsew signal tristate
rlabel metal2 s 261114 163200 261170 164400 6 la_oenb[77]
port 426 nsew signal tristate
rlabel metal2 s 264426 163200 264482 164400 6 la_oenb[78]
port 427 nsew signal tristate
rlabel metal2 s 267830 163200 267886 164400 6 la_oenb[79]
port 428 nsew signal tristate
rlabel metal2 s 25594 163200 25650 164400 6 la_oenb[7]
port 429 nsew signal tristate
rlabel metal2 s 271234 163200 271290 164400 6 la_oenb[80]
port 430 nsew signal tristate
rlabel metal2 s 274546 163200 274602 164400 6 la_oenb[81]
port 431 nsew signal tristate
rlabel metal2 s 277950 163200 278006 164400 6 la_oenb[82]
port 432 nsew signal tristate
rlabel metal2 s 281262 163200 281318 164400 6 la_oenb[83]
port 433 nsew signal tristate
rlabel metal2 s 284666 163200 284722 164400 6 la_oenb[84]
port 434 nsew signal tristate
rlabel metal2 s 287978 163200 288034 164400 6 la_oenb[85]
port 435 nsew signal tristate
rlabel metal2 s 291382 163200 291438 164400 6 la_oenb[86]
port 436 nsew signal tristate
rlabel metal2 s 294786 163200 294842 164400 6 la_oenb[87]
port 437 nsew signal tristate
rlabel metal2 s 298098 163200 298154 164400 6 la_oenb[88]
port 438 nsew signal tristate
rlabel metal2 s 301502 163200 301558 164400 6 la_oenb[89]
port 439 nsew signal tristate
rlabel metal2 s 28906 163200 28962 164400 6 la_oenb[8]
port 440 nsew signal tristate
rlabel metal2 s 304814 163200 304870 164400 6 la_oenb[90]
port 441 nsew signal tristate
rlabel metal2 s 308218 163200 308274 164400 6 la_oenb[91]
port 442 nsew signal tristate
rlabel metal2 s 311530 163200 311586 164400 6 la_oenb[92]
port 443 nsew signal tristate
rlabel metal2 s 314934 163200 314990 164400 6 la_oenb[93]
port 444 nsew signal tristate
rlabel metal2 s 318338 163200 318394 164400 6 la_oenb[94]
port 445 nsew signal tristate
rlabel metal2 s 321650 163200 321706 164400 6 la_oenb[95]
port 446 nsew signal tristate
rlabel metal2 s 325054 163200 325110 164400 6 la_oenb[96]
port 447 nsew signal tristate
rlabel metal2 s 328366 163200 328422 164400 6 la_oenb[97]
port 448 nsew signal tristate
rlabel metal2 s 331770 163200 331826 164400 6 la_oenb[98]
port 449 nsew signal tristate
rlabel metal2 s 335082 163200 335138 164400 6 la_oenb[99]
port 450 nsew signal tristate
rlabel metal2 s 32310 163200 32366 164400 6 la_oenb[9]
port 451 nsew signal tristate
rlabel metal2 s 2870 163200 2926 164400 6 la_output[0]
port 452 nsew signal tristate
rlabel metal2 s 339314 163200 339370 164400 6 la_output[100]
port 453 nsew signal tristate
rlabel metal2 s 342718 163200 342774 164400 6 la_output[101]
port 454 nsew signal tristate
rlabel metal2 s 346030 163200 346086 164400 6 la_output[102]
port 455 nsew signal tristate
rlabel metal2 s 349434 163200 349490 164400 6 la_output[103]
port 456 nsew signal tristate
rlabel metal2 s 352746 163200 352802 164400 6 la_output[104]
port 457 nsew signal tristate
rlabel metal2 s 356150 163200 356206 164400 6 la_output[105]
port 458 nsew signal tristate
rlabel metal2 s 359554 163200 359610 164400 6 la_output[106]
port 459 nsew signal tristate
rlabel metal2 s 362866 163200 362922 164400 6 la_output[107]
port 460 nsew signal tristate
rlabel metal2 s 366270 163200 366326 164400 6 la_output[108]
port 461 nsew signal tristate
rlabel metal2 s 369582 163200 369638 164400 6 la_output[109]
port 462 nsew signal tristate
rlabel metal2 s 36542 163200 36598 164400 6 la_output[10]
port 463 nsew signal tristate
rlabel metal2 s 372986 163200 373042 164400 6 la_output[110]
port 464 nsew signal tristate
rlabel metal2 s 376298 163200 376354 164400 6 la_output[111]
port 465 nsew signal tristate
rlabel metal2 s 379702 163200 379758 164400 6 la_output[112]
port 466 nsew signal tristate
rlabel metal2 s 383106 163200 383162 164400 6 la_output[113]
port 467 nsew signal tristate
rlabel metal2 s 386418 163200 386474 164400 6 la_output[114]
port 468 nsew signal tristate
rlabel metal2 s 389822 163200 389878 164400 6 la_output[115]
port 469 nsew signal tristate
rlabel metal2 s 393134 163200 393190 164400 6 la_output[116]
port 470 nsew signal tristate
rlabel metal2 s 396538 163200 396594 164400 6 la_output[117]
port 471 nsew signal tristate
rlabel metal2 s 399850 163200 399906 164400 6 la_output[118]
port 472 nsew signal tristate
rlabel metal2 s 403254 163200 403310 164400 6 la_output[119]
port 473 nsew signal tristate
rlabel metal2 s 39854 163200 39910 164400 6 la_output[11]
port 474 nsew signal tristate
rlabel metal2 s 406658 163200 406714 164400 6 la_output[120]
port 475 nsew signal tristate
rlabel metal2 s 409970 163200 410026 164400 6 la_output[121]
port 476 nsew signal tristate
rlabel metal2 s 413374 163200 413430 164400 6 la_output[122]
port 477 nsew signal tristate
rlabel metal2 s 416686 163200 416742 164400 6 la_output[123]
port 478 nsew signal tristate
rlabel metal2 s 420090 163200 420146 164400 6 la_output[124]
port 479 nsew signal tristate
rlabel metal2 s 423402 163200 423458 164400 6 la_output[125]
port 480 nsew signal tristate
rlabel metal2 s 426806 163200 426862 164400 6 la_output[126]
port 481 nsew signal tristate
rlabel metal2 s 430210 163200 430266 164400 6 la_output[127]
port 482 nsew signal tristate
rlabel metal2 s 43258 163200 43314 164400 6 la_output[12]
port 483 nsew signal tristate
rlabel metal2 s 46570 163200 46626 164400 6 la_output[13]
port 484 nsew signal tristate
rlabel metal2 s 49974 163200 50030 164400 6 la_output[14]
port 485 nsew signal tristate
rlabel metal2 s 53378 163200 53434 164400 6 la_output[15]
port 486 nsew signal tristate
rlabel metal2 s 56690 163200 56746 164400 6 la_output[16]
port 487 nsew signal tristate
rlabel metal2 s 60094 163200 60150 164400 6 la_output[17]
port 488 nsew signal tristate
rlabel metal2 s 63406 163200 63462 164400 6 la_output[18]
port 489 nsew signal tristate
rlabel metal2 s 66810 163200 66866 164400 6 la_output[19]
port 490 nsew signal tristate
rlabel metal2 s 6274 163200 6330 164400 6 la_output[1]
port 491 nsew signal tristate
rlabel metal2 s 70122 163200 70178 164400 6 la_output[20]
port 492 nsew signal tristate
rlabel metal2 s 73526 163200 73582 164400 6 la_output[21]
port 493 nsew signal tristate
rlabel metal2 s 76930 163200 76986 164400 6 la_output[22]
port 494 nsew signal tristate
rlabel metal2 s 80242 163200 80298 164400 6 la_output[23]
port 495 nsew signal tristate
rlabel metal2 s 83646 163200 83702 164400 6 la_output[24]
port 496 nsew signal tristate
rlabel metal2 s 86958 163200 87014 164400 6 la_output[25]
port 497 nsew signal tristate
rlabel metal2 s 90362 163200 90418 164400 6 la_output[26]
port 498 nsew signal tristate
rlabel metal2 s 93674 163200 93730 164400 6 la_output[27]
port 499 nsew signal tristate
rlabel metal2 s 97078 163200 97134 164400 6 la_output[28]
port 500 nsew signal tristate
rlabel metal2 s 100482 163200 100538 164400 6 la_output[29]
port 501 nsew signal tristate
rlabel metal2 s 9586 163200 9642 164400 6 la_output[2]
port 502 nsew signal tristate
rlabel metal2 s 103794 163200 103850 164400 6 la_output[30]
port 503 nsew signal tristate
rlabel metal2 s 107198 163200 107254 164400 6 la_output[31]
port 504 nsew signal tristate
rlabel metal2 s 110510 163200 110566 164400 6 la_output[32]
port 505 nsew signal tristate
rlabel metal2 s 113914 163200 113970 164400 6 la_output[33]
port 506 nsew signal tristate
rlabel metal2 s 117226 163200 117282 164400 6 la_output[34]
port 507 nsew signal tristate
rlabel metal2 s 120630 163200 120686 164400 6 la_output[35]
port 508 nsew signal tristate
rlabel metal2 s 124034 163200 124090 164400 6 la_output[36]
port 509 nsew signal tristate
rlabel metal2 s 127346 163200 127402 164400 6 la_output[37]
port 510 nsew signal tristate
rlabel metal2 s 130750 163200 130806 164400 6 la_output[38]
port 511 nsew signal tristate
rlabel metal2 s 134062 163200 134118 164400 6 la_output[39]
port 512 nsew signal tristate
rlabel metal2 s 12990 163200 13046 164400 6 la_output[3]
port 513 nsew signal tristate
rlabel metal2 s 137466 163200 137522 164400 6 la_output[40]
port 514 nsew signal tristate
rlabel metal2 s 140778 163200 140834 164400 6 la_output[41]
port 515 nsew signal tristate
rlabel metal2 s 144182 163200 144238 164400 6 la_output[42]
port 516 nsew signal tristate
rlabel metal2 s 147586 163200 147642 164400 6 la_output[43]
port 517 nsew signal tristate
rlabel metal2 s 150898 163200 150954 164400 6 la_output[44]
port 518 nsew signal tristate
rlabel metal2 s 154302 163200 154358 164400 6 la_output[45]
port 519 nsew signal tristate
rlabel metal2 s 157614 163200 157670 164400 6 la_output[46]
port 520 nsew signal tristate
rlabel metal2 s 161018 163200 161074 164400 6 la_output[47]
port 521 nsew signal tristate
rlabel metal2 s 164330 163200 164386 164400 6 la_output[48]
port 522 nsew signal tristate
rlabel metal2 s 167734 163200 167790 164400 6 la_output[49]
port 523 nsew signal tristate
rlabel metal2 s 16302 163200 16358 164400 6 la_output[4]
port 524 nsew signal tristate
rlabel metal2 s 171138 163200 171194 164400 6 la_output[50]
port 525 nsew signal tristate
rlabel metal2 s 174450 163200 174506 164400 6 la_output[51]
port 526 nsew signal tristate
rlabel metal2 s 177854 163200 177910 164400 6 la_output[52]
port 527 nsew signal tristate
rlabel metal2 s 181166 163200 181222 164400 6 la_output[53]
port 528 nsew signal tristate
rlabel metal2 s 184570 163200 184626 164400 6 la_output[54]
port 529 nsew signal tristate
rlabel metal2 s 187882 163200 187938 164400 6 la_output[55]
port 530 nsew signal tristate
rlabel metal2 s 191286 163200 191342 164400 6 la_output[56]
port 531 nsew signal tristate
rlabel metal2 s 194690 163200 194746 164400 6 la_output[57]
port 532 nsew signal tristate
rlabel metal2 s 198002 163200 198058 164400 6 la_output[58]
port 533 nsew signal tristate
rlabel metal2 s 201406 163200 201462 164400 6 la_output[59]
port 534 nsew signal tristate
rlabel metal2 s 19706 163200 19762 164400 6 la_output[5]
port 535 nsew signal tristate
rlabel metal2 s 204718 163200 204774 164400 6 la_output[60]
port 536 nsew signal tristate
rlabel metal2 s 208122 163200 208178 164400 6 la_output[61]
port 537 nsew signal tristate
rlabel metal2 s 211434 163200 211490 164400 6 la_output[62]
port 538 nsew signal tristate
rlabel metal2 s 214838 163200 214894 164400 6 la_output[63]
port 539 nsew signal tristate
rlabel metal2 s 218242 163200 218298 164400 6 la_output[64]
port 540 nsew signal tristate
rlabel metal2 s 221554 163200 221610 164400 6 la_output[65]
port 541 nsew signal tristate
rlabel metal2 s 224958 163200 225014 164400 6 la_output[66]
port 542 nsew signal tristate
rlabel metal2 s 228270 163200 228326 164400 6 la_output[67]
port 543 nsew signal tristate
rlabel metal2 s 231674 163200 231730 164400 6 la_output[68]
port 544 nsew signal tristate
rlabel metal2 s 234986 163200 235042 164400 6 la_output[69]
port 545 nsew signal tristate
rlabel metal2 s 23018 163200 23074 164400 6 la_output[6]
port 546 nsew signal tristate
rlabel metal2 s 238390 163200 238446 164400 6 la_output[70]
port 547 nsew signal tristate
rlabel metal2 s 241794 163200 241850 164400 6 la_output[71]
port 548 nsew signal tristate
rlabel metal2 s 245106 163200 245162 164400 6 la_output[72]
port 549 nsew signal tristate
rlabel metal2 s 248510 163200 248566 164400 6 la_output[73]
port 550 nsew signal tristate
rlabel metal2 s 251822 163200 251878 164400 6 la_output[74]
port 551 nsew signal tristate
rlabel metal2 s 255226 163200 255282 164400 6 la_output[75]
port 552 nsew signal tristate
rlabel metal2 s 258538 163200 258594 164400 6 la_output[76]
port 553 nsew signal tristate
rlabel metal2 s 261942 163200 261998 164400 6 la_output[77]
port 554 nsew signal tristate
rlabel metal2 s 265346 163200 265402 164400 6 la_output[78]
port 555 nsew signal tristate
rlabel metal2 s 268658 163200 268714 164400 6 la_output[79]
port 556 nsew signal tristate
rlabel metal2 s 26422 163200 26478 164400 6 la_output[7]
port 557 nsew signal tristate
rlabel metal2 s 272062 163200 272118 164400 6 la_output[80]
port 558 nsew signal tristate
rlabel metal2 s 275374 163200 275430 164400 6 la_output[81]
port 559 nsew signal tristate
rlabel metal2 s 278778 163200 278834 164400 6 la_output[82]
port 560 nsew signal tristate
rlabel metal2 s 282090 163200 282146 164400 6 la_output[83]
port 561 nsew signal tristate
rlabel metal2 s 285494 163200 285550 164400 6 la_output[84]
port 562 nsew signal tristate
rlabel metal2 s 288898 163200 288954 164400 6 la_output[85]
port 563 nsew signal tristate
rlabel metal2 s 292210 163200 292266 164400 6 la_output[86]
port 564 nsew signal tristate
rlabel metal2 s 295614 163200 295670 164400 6 la_output[87]
port 565 nsew signal tristate
rlabel metal2 s 298926 163200 298982 164400 6 la_output[88]
port 566 nsew signal tristate
rlabel metal2 s 302330 163200 302386 164400 6 la_output[89]
port 567 nsew signal tristate
rlabel metal2 s 29826 163200 29882 164400 6 la_output[8]
port 568 nsew signal tristate
rlabel metal2 s 305642 163200 305698 164400 6 la_output[90]
port 569 nsew signal tristate
rlabel metal2 s 309046 163200 309102 164400 6 la_output[91]
port 570 nsew signal tristate
rlabel metal2 s 312450 163200 312506 164400 6 la_output[92]
port 571 nsew signal tristate
rlabel metal2 s 315762 163200 315818 164400 6 la_output[93]
port 572 nsew signal tristate
rlabel metal2 s 319166 163200 319222 164400 6 la_output[94]
port 573 nsew signal tristate
rlabel metal2 s 322478 163200 322534 164400 6 la_output[95]
port 574 nsew signal tristate
rlabel metal2 s 325882 163200 325938 164400 6 la_output[96]
port 575 nsew signal tristate
rlabel metal2 s 329194 163200 329250 164400 6 la_output[97]
port 576 nsew signal tristate
rlabel metal2 s 332598 163200 332654 164400 6 la_output[98]
port 577 nsew signal tristate
rlabel metal2 s 336002 163200 336058 164400 6 la_output[99]
port 578 nsew signal tristate
rlabel metal2 s 33138 163200 33194 164400 6 la_output[9]
port 579 nsew signal tristate
rlabel metal2 s 431038 163200 431094 164400 6 mprj_ack_i
port 580 nsew signal input
rlabel metal2 s 435178 163200 435234 164400 6 mprj_adr_o[0]
port 581 nsew signal tristate
rlabel metal2 s 463790 163200 463846 164400 6 mprj_adr_o[10]
port 582 nsew signal tristate
rlabel metal2 s 466366 163200 466422 164400 6 mprj_adr_o[11]
port 583 nsew signal tristate
rlabel metal2 s 468850 163200 468906 164400 6 mprj_adr_o[12]
port 584 nsew signal tristate
rlabel metal2 s 471426 163200 471482 164400 6 mprj_adr_o[13]
port 585 nsew signal tristate
rlabel metal2 s 473910 163200 473966 164400 6 mprj_adr_o[14]
port 586 nsew signal tristate
rlabel metal2 s 476394 163200 476450 164400 6 mprj_adr_o[15]
port 587 nsew signal tristate
rlabel metal2 s 478970 163200 479026 164400 6 mprj_adr_o[16]
port 588 nsew signal tristate
rlabel metal2 s 481454 163200 481510 164400 6 mprj_adr_o[17]
port 589 nsew signal tristate
rlabel metal2 s 484030 163200 484086 164400 6 mprj_adr_o[18]
port 590 nsew signal tristate
rlabel metal2 s 486514 163200 486570 164400 6 mprj_adr_o[19]
port 591 nsew signal tristate
rlabel metal2 s 438582 163200 438638 164400 6 mprj_adr_o[1]
port 592 nsew signal tristate
rlabel metal2 s 489090 163200 489146 164400 6 mprj_adr_o[20]
port 593 nsew signal tristate
rlabel metal2 s 491574 163200 491630 164400 6 mprj_adr_o[21]
port 594 nsew signal tristate
rlabel metal2 s 494058 163200 494114 164400 6 mprj_adr_o[22]
port 595 nsew signal tristate
rlabel metal2 s 496634 163200 496690 164400 6 mprj_adr_o[23]
port 596 nsew signal tristate
rlabel metal2 s 499118 163200 499174 164400 6 mprj_adr_o[24]
port 597 nsew signal tristate
rlabel metal2 s 501694 163200 501750 164400 6 mprj_adr_o[25]
port 598 nsew signal tristate
rlabel metal2 s 504178 163200 504234 164400 6 mprj_adr_o[26]
port 599 nsew signal tristate
rlabel metal2 s 506754 163200 506810 164400 6 mprj_adr_o[27]
port 600 nsew signal tristate
rlabel metal2 s 509238 163200 509294 164400 6 mprj_adr_o[28]
port 601 nsew signal tristate
rlabel metal2 s 511722 163200 511778 164400 6 mprj_adr_o[29]
port 602 nsew signal tristate
rlabel metal2 s 441986 163200 442042 164400 6 mprj_adr_o[2]
port 603 nsew signal tristate
rlabel metal2 s 514298 163200 514354 164400 6 mprj_adr_o[30]
port 604 nsew signal tristate
rlabel metal2 s 516782 163200 516838 164400 6 mprj_adr_o[31]
port 605 nsew signal tristate
rlabel metal2 s 445298 163200 445354 164400 6 mprj_adr_o[3]
port 606 nsew signal tristate
rlabel metal2 s 448702 163200 448758 164400 6 mprj_adr_o[4]
port 607 nsew signal tristate
rlabel metal2 s 451186 163200 451242 164400 6 mprj_adr_o[5]
port 608 nsew signal tristate
rlabel metal2 s 453762 163200 453818 164400 6 mprj_adr_o[6]
port 609 nsew signal tristate
rlabel metal2 s 456246 163200 456302 164400 6 mprj_adr_o[7]
port 610 nsew signal tristate
rlabel metal2 s 458730 163200 458786 164400 6 mprj_adr_o[8]
port 611 nsew signal tristate
rlabel metal2 s 461306 163200 461362 164400 6 mprj_adr_o[9]
port 612 nsew signal tristate
rlabel metal2 s 431866 163200 431922 164400 6 mprj_cyc_o
port 613 nsew signal tristate
rlabel metal2 s 436098 163200 436154 164400 6 mprj_dat_i[0]
port 614 nsew signal input
rlabel metal2 s 464618 163200 464674 164400 6 mprj_dat_i[10]
port 615 nsew signal input
rlabel metal2 s 467194 163200 467250 164400 6 mprj_dat_i[11]
port 616 nsew signal input
rlabel metal2 s 469678 163200 469734 164400 6 mprj_dat_i[12]
port 617 nsew signal input
rlabel metal2 s 472254 163200 472310 164400 6 mprj_dat_i[13]
port 618 nsew signal input
rlabel metal2 s 474738 163200 474794 164400 6 mprj_dat_i[14]
port 619 nsew signal input
rlabel metal2 s 477314 163200 477370 164400 6 mprj_dat_i[15]
port 620 nsew signal input
rlabel metal2 s 479798 163200 479854 164400 6 mprj_dat_i[16]
port 621 nsew signal input
rlabel metal2 s 482282 163200 482338 164400 6 mprj_dat_i[17]
port 622 nsew signal input
rlabel metal2 s 484858 163200 484914 164400 6 mprj_dat_i[18]
port 623 nsew signal input
rlabel metal2 s 487342 163200 487398 164400 6 mprj_dat_i[19]
port 624 nsew signal input
rlabel metal2 s 439410 163200 439466 164400 6 mprj_dat_i[1]
port 625 nsew signal input
rlabel metal2 s 489918 163200 489974 164400 6 mprj_dat_i[20]
port 626 nsew signal input
rlabel metal2 s 492402 163200 492458 164400 6 mprj_dat_i[21]
port 627 nsew signal input
rlabel metal2 s 494978 163200 495034 164400 6 mprj_dat_i[22]
port 628 nsew signal input
rlabel metal2 s 497462 163200 497518 164400 6 mprj_dat_i[23]
port 629 nsew signal input
rlabel metal2 s 499946 163200 500002 164400 6 mprj_dat_i[24]
port 630 nsew signal input
rlabel metal2 s 502522 163200 502578 164400 6 mprj_dat_i[25]
port 631 nsew signal input
rlabel metal2 s 505006 163200 505062 164400 6 mprj_dat_i[26]
port 632 nsew signal input
rlabel metal2 s 507582 163200 507638 164400 6 mprj_dat_i[27]
port 633 nsew signal input
rlabel metal2 s 510066 163200 510122 164400 6 mprj_dat_i[28]
port 634 nsew signal input
rlabel metal2 s 512642 163200 512698 164400 6 mprj_dat_i[29]
port 635 nsew signal input
rlabel metal2 s 442814 163200 442870 164400 6 mprj_dat_i[2]
port 636 nsew signal input
rlabel metal2 s 515126 163200 515182 164400 6 mprj_dat_i[30]
port 637 nsew signal input
rlabel metal2 s 517610 163200 517666 164400 6 mprj_dat_i[31]
port 638 nsew signal input
rlabel metal2 s 446126 163200 446182 164400 6 mprj_dat_i[3]
port 639 nsew signal input
rlabel metal2 s 449530 163200 449586 164400 6 mprj_dat_i[4]
port 640 nsew signal input
rlabel metal2 s 452014 163200 452070 164400 6 mprj_dat_i[5]
port 641 nsew signal input
rlabel metal2 s 454590 163200 454646 164400 6 mprj_dat_i[6]
port 642 nsew signal input
rlabel metal2 s 457074 163200 457130 164400 6 mprj_dat_i[7]
port 643 nsew signal input
rlabel metal2 s 459650 163200 459706 164400 6 mprj_dat_i[8]
port 644 nsew signal input
rlabel metal2 s 462134 163200 462190 164400 6 mprj_dat_i[9]
port 645 nsew signal input
rlabel metal2 s 436926 163200 436982 164400 6 mprj_dat_o[0]
port 646 nsew signal tristate
rlabel metal2 s 465538 163200 465594 164400 6 mprj_dat_o[10]
port 647 nsew signal tristate
rlabel metal2 s 468022 163200 468078 164400 6 mprj_dat_o[11]
port 648 nsew signal tristate
rlabel metal2 s 470506 163200 470562 164400 6 mprj_dat_o[12]
port 649 nsew signal tristate
rlabel metal2 s 473082 163200 473138 164400 6 mprj_dat_o[13]
port 650 nsew signal tristate
rlabel metal2 s 475566 163200 475622 164400 6 mprj_dat_o[14]
port 651 nsew signal tristate
rlabel metal2 s 478142 163200 478198 164400 6 mprj_dat_o[15]
port 652 nsew signal tristate
rlabel metal2 s 480626 163200 480682 164400 6 mprj_dat_o[16]
port 653 nsew signal tristate
rlabel metal2 s 483202 163200 483258 164400 6 mprj_dat_o[17]
port 654 nsew signal tristate
rlabel metal2 s 485686 163200 485742 164400 6 mprj_dat_o[18]
port 655 nsew signal tristate
rlabel metal2 s 488170 163200 488226 164400 6 mprj_dat_o[19]
port 656 nsew signal tristate
rlabel metal2 s 440238 163200 440294 164400 6 mprj_dat_o[1]
port 657 nsew signal tristate
rlabel metal2 s 490746 163200 490802 164400 6 mprj_dat_o[20]
port 658 nsew signal tristate
rlabel metal2 s 493230 163200 493286 164400 6 mprj_dat_o[21]
port 659 nsew signal tristate
rlabel metal2 s 495806 163200 495862 164400 6 mprj_dat_o[22]
port 660 nsew signal tristate
rlabel metal2 s 498290 163200 498346 164400 6 mprj_dat_o[23]
port 661 nsew signal tristate
rlabel metal2 s 500866 163200 500922 164400 6 mprj_dat_o[24]
port 662 nsew signal tristate
rlabel metal2 s 503350 163200 503406 164400 6 mprj_dat_o[25]
port 663 nsew signal tristate
rlabel metal2 s 505834 163200 505890 164400 6 mprj_dat_o[26]
port 664 nsew signal tristate
rlabel metal2 s 508410 163200 508466 164400 6 mprj_dat_o[27]
port 665 nsew signal tristate
rlabel metal2 s 510894 163200 510950 164400 6 mprj_dat_o[28]
port 666 nsew signal tristate
rlabel metal2 s 513470 163200 513526 164400 6 mprj_dat_o[29]
port 667 nsew signal tristate
rlabel metal2 s 443642 163200 443698 164400 6 mprj_dat_o[2]
port 668 nsew signal tristate
rlabel metal2 s 515954 163200 516010 164400 6 mprj_dat_o[30]
port 669 nsew signal tristate
rlabel metal2 s 518530 163200 518586 164400 6 mprj_dat_o[31]
port 670 nsew signal tristate
rlabel metal2 s 446954 163200 447010 164400 6 mprj_dat_o[3]
port 671 nsew signal tristate
rlabel metal2 s 450358 163200 450414 164400 6 mprj_dat_o[4]
port 672 nsew signal tristate
rlabel metal2 s 452842 163200 452898 164400 6 mprj_dat_o[5]
port 673 nsew signal tristate
rlabel metal2 s 455418 163200 455474 164400 6 mprj_dat_o[6]
port 674 nsew signal tristate
rlabel metal2 s 457902 163200 457958 164400 6 mprj_dat_o[7]
port 675 nsew signal tristate
rlabel metal2 s 460478 163200 460534 164400 6 mprj_dat_o[8]
port 676 nsew signal tristate
rlabel metal2 s 462962 163200 463018 164400 6 mprj_dat_o[9]
port 677 nsew signal tristate
rlabel metal2 s 437754 163200 437810 164400 6 mprj_sel_o[0]
port 678 nsew signal tristate
rlabel metal2 s 441066 163200 441122 164400 6 mprj_sel_o[1]
port 679 nsew signal tristate
rlabel metal2 s 444470 163200 444526 164400 6 mprj_sel_o[2]
port 680 nsew signal tristate
rlabel metal2 s 447874 163200 447930 164400 6 mprj_sel_o[3]
port 681 nsew signal tristate
rlabel metal2 s 432694 163200 432750 164400 6 mprj_stb_o
port 682 nsew signal tristate
rlabel metal2 s 433522 163200 433578 164400 6 mprj_wb_iena
port 683 nsew signal tristate
rlabel metal2 s 434350 163200 434406 164400 6 mprj_we_o
port 684 nsew signal tristate
rlabel metal3 s 523200 90176 524400 90296 6 qspi_enabled
port 685 nsew signal tristate
rlabel metal3 s 523200 84192 524400 84312 6 ser_rx
port 686 nsew signal input
rlabel metal3 s 523200 85688 524400 85808 6 ser_tx
port 687 nsew signal tristate
rlabel metal3 s 523200 81064 524400 81184 6 spi_csb
port 688 nsew signal tristate
rlabel metal3 s 523200 87184 524400 87304 6 spi_enabled
port 689 nsew signal tristate
rlabel metal3 s 523200 79568 524400 79688 6 spi_sck
port 690 nsew signal tristate
rlabel metal3 s 523200 82696 524400 82816 6 spi_sdi
port 691 nsew signal input
rlabel metal3 s 523200 78072 524400 78192 6 spi_sdo
port 692 nsew signal tristate
rlabel metal3 s 523200 76576 524400 76696 6 spi_sdoenb
port 693 nsew signal tristate
rlabel metal3 s 523200 2184 524400 2304 6 sram_ro_addr[0]
port 694 nsew signal input
rlabel metal3 s 523200 3680 524400 3800 6 sram_ro_addr[1]
port 695 nsew signal input
rlabel metal3 s 523200 5176 524400 5296 6 sram_ro_addr[2]
port 696 nsew signal input
rlabel metal3 s 523200 6672 524400 6792 6 sram_ro_addr[3]
port 697 nsew signal input
rlabel metal3 s 523200 8168 524400 8288 6 sram_ro_addr[4]
port 698 nsew signal input
rlabel metal3 s 523200 9800 524400 9920 6 sram_ro_addr[5]
port 699 nsew signal input
rlabel metal3 s 523200 11296 524400 11416 6 sram_ro_addr[6]
port 700 nsew signal input
rlabel metal3 s 523200 12792 524400 12912 6 sram_ro_addr[7]
port 701 nsew signal input
rlabel metal3 s 523200 14288 524400 14408 6 sram_ro_clk
port 702 nsew signal input
rlabel metal3 s 523200 688 524400 808 6 sram_ro_csb
port 703 nsew signal input
rlabel metal3 s 523200 15784 524400 15904 6 sram_ro_data[0]
port 704 nsew signal tristate
rlabel metal3 s 523200 31016 524400 31136 6 sram_ro_data[10]
port 705 nsew signal tristate
rlabel metal3 s 523200 32512 524400 32632 6 sram_ro_data[11]
port 706 nsew signal tristate
rlabel metal3 s 523200 34008 524400 34128 6 sram_ro_data[12]
port 707 nsew signal tristate
rlabel metal3 s 523200 35504 524400 35624 6 sram_ro_data[13]
port 708 nsew signal tristate
rlabel metal3 s 523200 37136 524400 37256 6 sram_ro_data[14]
port 709 nsew signal tristate
rlabel metal3 s 523200 38632 524400 38752 6 sram_ro_data[15]
port 710 nsew signal tristate
rlabel metal3 s 523200 40128 524400 40248 6 sram_ro_data[16]
port 711 nsew signal tristate
rlabel metal3 s 523200 41624 524400 41744 6 sram_ro_data[17]
port 712 nsew signal tristate
rlabel metal3 s 523200 43120 524400 43240 6 sram_ro_data[18]
port 713 nsew signal tristate
rlabel metal3 s 523200 44616 524400 44736 6 sram_ro_data[19]
port 714 nsew signal tristate
rlabel metal3 s 523200 17280 524400 17400 6 sram_ro_data[1]
port 715 nsew signal tristate
rlabel metal3 s 523200 46248 524400 46368 6 sram_ro_data[20]
port 716 nsew signal tristate
rlabel metal3 s 523200 47744 524400 47864 6 sram_ro_data[21]
port 717 nsew signal tristate
rlabel metal3 s 523200 49240 524400 49360 6 sram_ro_data[22]
port 718 nsew signal tristate
rlabel metal3 s 523200 50736 524400 50856 6 sram_ro_data[23]
port 719 nsew signal tristate
rlabel metal3 s 523200 52232 524400 52352 6 sram_ro_data[24]
port 720 nsew signal tristate
rlabel metal3 s 523200 53728 524400 53848 6 sram_ro_data[25]
port 721 nsew signal tristate
rlabel metal3 s 523200 55360 524400 55480 6 sram_ro_data[26]
port 722 nsew signal tristate
rlabel metal3 s 523200 56856 524400 56976 6 sram_ro_data[27]
port 723 nsew signal tristate
rlabel metal3 s 523200 58352 524400 58472 6 sram_ro_data[28]
port 724 nsew signal tristate
rlabel metal3 s 523200 59848 524400 59968 6 sram_ro_data[29]
port 725 nsew signal tristate
rlabel metal3 s 523200 18912 524400 19032 6 sram_ro_data[2]
port 726 nsew signal tristate
rlabel metal3 s 523200 61344 524400 61464 6 sram_ro_data[30]
port 727 nsew signal tristate
rlabel metal3 s 523200 62840 524400 62960 6 sram_ro_data[31]
port 728 nsew signal tristate
rlabel metal3 s 523200 20408 524400 20528 6 sram_ro_data[3]
port 729 nsew signal tristate
rlabel metal3 s 523200 21904 524400 22024 6 sram_ro_data[4]
port 730 nsew signal tristate
rlabel metal3 s 523200 23400 524400 23520 6 sram_ro_data[5]
port 731 nsew signal tristate
rlabel metal3 s 523200 24896 524400 25016 6 sram_ro_data[6]
port 732 nsew signal tristate
rlabel metal3 s 523200 26392 524400 26512 6 sram_ro_data[7]
port 733 nsew signal tristate
rlabel metal3 s 523200 28024 524400 28144 6 sram_ro_data[8]
port 734 nsew signal tristate
rlabel metal3 s 523200 29520 524400 29640 6 sram_ro_data[9]
port 735 nsew signal tristate
rlabel metal3 s 523200 70456 524400 70576 6 trap
port 736 nsew signal tristate
rlabel metal3 s 523200 88680 524400 88800 6 uart_enabled
port 737 nsew signal tristate
rlabel metal2 s 519358 163200 519414 164400 6 user_irq_ena[0]
port 738 nsew signal tristate
rlabel metal2 s 520186 163200 520242 164400 6 user_irq_ena[1]
port 739 nsew signal tristate
rlabel metal2 s 521014 163200 521070 164400 6 user_irq_ena[2]
port 740 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 524000 164000
<< end >>
