magic
tech sky130A
magscale 1 2
timestamp 1638405022
<< obsli1 >>
rect 2869 4159 516900 147809
<< obsm1 >>
rect 382 688 523558 160132
<< metal2 >>
rect 386 163200 442 164400
rect 1214 163200 1270 164400
rect 2042 163200 2098 164400
rect 2870 163200 2926 164400
rect 3698 163200 3754 164400
rect 4526 163200 4582 164400
rect 5354 163200 5410 164400
rect 6182 163200 6238 164400
rect 7102 163200 7158 164400
rect 7930 163200 7986 164400
rect 8758 163200 8814 164400
rect 9586 163200 9642 164400
rect 10414 163200 10470 164400
rect 11242 163200 11298 164400
rect 12070 163200 12126 164400
rect 12898 163200 12954 164400
rect 13818 163200 13874 164400
rect 14646 163200 14702 164400
rect 15474 163200 15530 164400
rect 16302 163200 16358 164400
rect 17130 163200 17186 164400
rect 17958 163200 18014 164400
rect 18786 163200 18842 164400
rect 19614 163200 19670 164400
rect 20534 163200 20590 164400
rect 21362 163200 21418 164400
rect 22190 163200 22246 164400
rect 23018 163200 23074 164400
rect 23846 163200 23902 164400
rect 24674 163200 24730 164400
rect 25502 163200 25558 164400
rect 26330 163200 26386 164400
rect 27250 163200 27306 164400
rect 28078 163200 28134 164400
rect 28906 163200 28962 164400
rect 29734 163200 29790 164400
rect 30562 163200 30618 164400
rect 31390 163200 31446 164400
rect 32218 163200 32274 164400
rect 33138 163200 33194 164400
rect 33966 163200 34022 164400
rect 34794 163200 34850 164400
rect 35622 163200 35678 164400
rect 36450 163200 36506 164400
rect 37278 163200 37334 164400
rect 38106 163200 38162 164400
rect 38934 163200 38990 164400
rect 39854 163200 39910 164400
rect 40682 163200 40738 164400
rect 41510 163200 41566 164400
rect 42338 163200 42394 164400
rect 43166 163200 43222 164400
rect 43994 163200 44050 164400
rect 44822 163200 44878 164400
rect 45650 163200 45706 164400
rect 46570 163200 46626 164400
rect 47398 163200 47454 164400
rect 48226 163200 48282 164400
rect 49054 163200 49110 164400
rect 49882 163200 49938 164400
rect 50710 163200 50766 164400
rect 51538 163200 51594 164400
rect 52366 163200 52422 164400
rect 53286 163200 53342 164400
rect 54114 163200 54170 164400
rect 54942 163200 54998 164400
rect 55770 163200 55826 164400
rect 56598 163200 56654 164400
rect 57426 163200 57482 164400
rect 58254 163200 58310 164400
rect 59082 163200 59138 164400
rect 60002 163200 60058 164400
rect 60830 163200 60886 164400
rect 61658 163200 61714 164400
rect 62486 163200 62542 164400
rect 63314 163200 63370 164400
rect 64142 163200 64198 164400
rect 64970 163200 65026 164400
rect 65890 163200 65946 164400
rect 66718 163200 66774 164400
rect 67546 163200 67602 164400
rect 68374 163200 68430 164400
rect 69202 163200 69258 164400
rect 70030 163200 70086 164400
rect 70858 163200 70914 164400
rect 71686 163200 71742 164400
rect 72606 163200 72662 164400
rect 73434 163200 73490 164400
rect 74262 163200 74318 164400
rect 75090 163200 75146 164400
rect 75918 163200 75974 164400
rect 76746 163200 76802 164400
rect 77574 163200 77630 164400
rect 78402 163200 78458 164400
rect 79322 163200 79378 164400
rect 80150 163200 80206 164400
rect 80978 163200 81034 164400
rect 81806 163200 81862 164400
rect 82634 163200 82690 164400
rect 83462 163200 83518 164400
rect 84290 163200 84346 164400
rect 85118 163200 85174 164400
rect 86038 163200 86094 164400
rect 86866 163200 86922 164400
rect 87694 163200 87750 164400
rect 88522 163200 88578 164400
rect 89350 163200 89406 164400
rect 90178 163200 90234 164400
rect 91006 163200 91062 164400
rect 91834 163200 91890 164400
rect 92754 163200 92810 164400
rect 93582 163200 93638 164400
rect 94410 163200 94466 164400
rect 95238 163200 95294 164400
rect 96066 163200 96122 164400
rect 96894 163200 96950 164400
rect 97722 163200 97778 164400
rect 98642 163200 98698 164400
rect 99470 163200 99526 164400
rect 100298 163200 100354 164400
rect 101126 163200 101182 164400
rect 101954 163200 102010 164400
rect 102782 163200 102838 164400
rect 103610 163200 103666 164400
rect 104438 163200 104494 164400
rect 105358 163200 105414 164400
rect 106186 163200 106242 164400
rect 107014 163200 107070 164400
rect 107842 163200 107898 164400
rect 108670 163200 108726 164400
rect 109498 163200 109554 164400
rect 110326 163200 110382 164400
rect 111154 163200 111210 164400
rect 112074 163200 112130 164400
rect 112902 163200 112958 164400
rect 113730 163200 113786 164400
rect 114558 163200 114614 164400
rect 115386 163200 115442 164400
rect 116214 163200 116270 164400
rect 117042 163200 117098 164400
rect 117870 163200 117926 164400
rect 118790 163200 118846 164400
rect 119618 163200 119674 164400
rect 120446 163200 120502 164400
rect 121274 163200 121330 164400
rect 122102 163200 122158 164400
rect 122930 163200 122986 164400
rect 123758 163200 123814 164400
rect 124586 163200 124642 164400
rect 125506 163200 125562 164400
rect 126334 163200 126390 164400
rect 127162 163200 127218 164400
rect 127990 163200 128046 164400
rect 128818 163200 128874 164400
rect 129646 163200 129702 164400
rect 130474 163200 130530 164400
rect 131394 163200 131450 164400
rect 132222 163200 132278 164400
rect 133050 163200 133106 164400
rect 133878 163200 133934 164400
rect 134706 163200 134762 164400
rect 135534 163200 135590 164400
rect 136362 163200 136418 164400
rect 137190 163200 137246 164400
rect 138110 163200 138166 164400
rect 138938 163200 138994 164400
rect 139766 163200 139822 164400
rect 140594 163200 140650 164400
rect 141422 163200 141478 164400
rect 142250 163200 142306 164400
rect 143078 163200 143134 164400
rect 143906 163200 143962 164400
rect 144826 163200 144882 164400
rect 145654 163200 145710 164400
rect 146482 163200 146538 164400
rect 147310 163200 147366 164400
rect 148138 163200 148194 164400
rect 148966 163200 149022 164400
rect 149794 163200 149850 164400
rect 150622 163200 150678 164400
rect 151542 163200 151598 164400
rect 152370 163200 152426 164400
rect 153198 163200 153254 164400
rect 154026 163200 154082 164400
rect 154854 163200 154910 164400
rect 155682 163200 155738 164400
rect 156510 163200 156566 164400
rect 157338 163200 157394 164400
rect 158258 163200 158314 164400
rect 159086 163200 159142 164400
rect 159914 163200 159970 164400
rect 160742 163200 160798 164400
rect 161570 163200 161626 164400
rect 162398 163200 162454 164400
rect 163226 163200 163282 164400
rect 164146 163200 164202 164400
rect 164974 163200 165030 164400
rect 165802 163200 165858 164400
rect 166630 163200 166686 164400
rect 167458 163200 167514 164400
rect 168286 163200 168342 164400
rect 169114 163200 169170 164400
rect 169942 163200 169998 164400
rect 170862 163200 170918 164400
rect 171690 163200 171746 164400
rect 172518 163200 172574 164400
rect 173346 163200 173402 164400
rect 174174 163200 174230 164400
rect 175002 163200 175058 164400
rect 175830 163200 175886 164400
rect 176658 163200 176714 164400
rect 177578 163200 177634 164400
rect 178406 163200 178462 164400
rect 179234 163200 179290 164400
rect 180062 163200 180118 164400
rect 180890 163200 180946 164400
rect 181718 163200 181774 164400
rect 182546 163200 182602 164400
rect 183374 163200 183430 164400
rect 184294 163200 184350 164400
rect 185122 163200 185178 164400
rect 185950 163200 186006 164400
rect 186778 163200 186834 164400
rect 187606 163200 187662 164400
rect 188434 163200 188490 164400
rect 189262 163200 189318 164400
rect 190090 163200 190146 164400
rect 191010 163200 191066 164400
rect 191838 163200 191894 164400
rect 192666 163200 192722 164400
rect 193494 163200 193550 164400
rect 194322 163200 194378 164400
rect 195150 163200 195206 164400
rect 195978 163200 196034 164400
rect 196898 163200 196954 164400
rect 197726 163200 197782 164400
rect 198554 163200 198610 164400
rect 199382 163200 199438 164400
rect 200210 163200 200266 164400
rect 201038 163200 201094 164400
rect 201866 163200 201922 164400
rect 202694 163200 202750 164400
rect 203614 163200 203670 164400
rect 204442 163200 204498 164400
rect 205270 163200 205326 164400
rect 206098 163200 206154 164400
rect 206926 163200 206982 164400
rect 207754 163200 207810 164400
rect 208582 163200 208638 164400
rect 209410 163200 209466 164400
rect 210330 163200 210386 164400
rect 211158 163200 211214 164400
rect 211986 163200 212042 164400
rect 212814 163200 212870 164400
rect 213642 163200 213698 164400
rect 214470 163200 214526 164400
rect 215298 163200 215354 164400
rect 216126 163200 216182 164400
rect 217046 163200 217102 164400
rect 217874 163200 217930 164400
rect 218702 163200 218758 164400
rect 219530 163200 219586 164400
rect 220358 163200 220414 164400
rect 221186 163200 221242 164400
rect 222014 163200 222070 164400
rect 222842 163200 222898 164400
rect 223762 163200 223818 164400
rect 224590 163200 224646 164400
rect 225418 163200 225474 164400
rect 226246 163200 226302 164400
rect 227074 163200 227130 164400
rect 227902 163200 227958 164400
rect 228730 163200 228786 164400
rect 229650 163200 229706 164400
rect 230478 163200 230534 164400
rect 231306 163200 231362 164400
rect 232134 163200 232190 164400
rect 232962 163200 233018 164400
rect 233790 163200 233846 164400
rect 234618 163200 234674 164400
rect 235446 163200 235502 164400
rect 236366 163200 236422 164400
rect 237194 163200 237250 164400
rect 238022 163200 238078 164400
rect 238850 163200 238906 164400
rect 239678 163200 239734 164400
rect 240506 163200 240562 164400
rect 241334 163200 241390 164400
rect 242162 163200 242218 164400
rect 243082 163200 243138 164400
rect 243910 163200 243966 164400
rect 244738 163200 244794 164400
rect 245566 163200 245622 164400
rect 246394 163200 246450 164400
rect 247222 163200 247278 164400
rect 248050 163200 248106 164400
rect 248878 163200 248934 164400
rect 249798 163200 249854 164400
rect 250626 163200 250682 164400
rect 251454 163200 251510 164400
rect 252282 163200 252338 164400
rect 253110 163200 253166 164400
rect 253938 163200 253994 164400
rect 254766 163200 254822 164400
rect 255594 163200 255650 164400
rect 256514 163200 256570 164400
rect 257342 163200 257398 164400
rect 258170 163200 258226 164400
rect 258998 163200 259054 164400
rect 259826 163200 259882 164400
rect 260654 163200 260710 164400
rect 261482 163200 261538 164400
rect 262402 163200 262458 164400
rect 263230 163200 263286 164400
rect 264058 163200 264114 164400
rect 264886 163200 264942 164400
rect 265714 163200 265770 164400
rect 266542 163200 266598 164400
rect 267370 163200 267426 164400
rect 268198 163200 268254 164400
rect 269118 163200 269174 164400
rect 269946 163200 270002 164400
rect 270774 163200 270830 164400
rect 271602 163200 271658 164400
rect 272430 163200 272486 164400
rect 273258 163200 273314 164400
rect 274086 163200 274142 164400
rect 274914 163200 274970 164400
rect 275834 163200 275890 164400
rect 276662 163200 276718 164400
rect 277490 163200 277546 164400
rect 278318 163200 278374 164400
rect 279146 163200 279202 164400
rect 279974 163200 280030 164400
rect 280802 163200 280858 164400
rect 281630 163200 281686 164400
rect 282550 163200 282606 164400
rect 283378 163200 283434 164400
rect 284206 163200 284262 164400
rect 285034 163200 285090 164400
rect 285862 163200 285918 164400
rect 286690 163200 286746 164400
rect 287518 163200 287574 164400
rect 288346 163200 288402 164400
rect 289266 163200 289322 164400
rect 290094 163200 290150 164400
rect 290922 163200 290978 164400
rect 291750 163200 291806 164400
rect 292578 163200 292634 164400
rect 293406 163200 293462 164400
rect 294234 163200 294290 164400
rect 295154 163200 295210 164400
rect 295982 163200 296038 164400
rect 296810 163200 296866 164400
rect 297638 163200 297694 164400
rect 298466 163200 298522 164400
rect 299294 163200 299350 164400
rect 300122 163200 300178 164400
rect 300950 163200 301006 164400
rect 301870 163200 301926 164400
rect 302698 163200 302754 164400
rect 303526 163200 303582 164400
rect 304354 163200 304410 164400
rect 305182 163200 305238 164400
rect 306010 163200 306066 164400
rect 306838 163200 306894 164400
rect 307666 163200 307722 164400
rect 308586 163200 308642 164400
rect 309414 163200 309470 164400
rect 310242 163200 310298 164400
rect 311070 163200 311126 164400
rect 311898 163200 311954 164400
rect 312726 163200 312782 164400
rect 313554 163200 313610 164400
rect 314382 163200 314438 164400
rect 315302 163200 315358 164400
rect 316130 163200 316186 164400
rect 316958 163200 317014 164400
rect 317786 163200 317842 164400
rect 318614 163200 318670 164400
rect 319442 163200 319498 164400
rect 320270 163200 320326 164400
rect 321098 163200 321154 164400
rect 322018 163200 322074 164400
rect 322846 163200 322902 164400
rect 323674 163200 323730 164400
rect 324502 163200 324558 164400
rect 325330 163200 325386 164400
rect 326158 163200 326214 164400
rect 326986 163200 327042 164400
rect 327906 163200 327962 164400
rect 328734 163200 328790 164400
rect 329562 163200 329618 164400
rect 330390 163200 330446 164400
rect 331218 163200 331274 164400
rect 332046 163200 332102 164400
rect 332874 163200 332930 164400
rect 333702 163200 333758 164400
rect 334622 163200 334678 164400
rect 335450 163200 335506 164400
rect 336278 163200 336334 164400
rect 337106 163200 337162 164400
rect 337934 163200 337990 164400
rect 338762 163200 338818 164400
rect 339590 163200 339646 164400
rect 340418 163200 340474 164400
rect 341338 163200 341394 164400
rect 342166 163200 342222 164400
rect 342994 163200 343050 164400
rect 343822 163200 343878 164400
rect 344650 163200 344706 164400
rect 345478 163200 345534 164400
rect 346306 163200 346362 164400
rect 347134 163200 347190 164400
rect 348054 163200 348110 164400
rect 348882 163200 348938 164400
rect 349710 163200 349766 164400
rect 350538 163200 350594 164400
rect 351366 163200 351422 164400
rect 352194 163200 352250 164400
rect 353022 163200 353078 164400
rect 353850 163200 353906 164400
rect 354770 163200 354826 164400
rect 355598 163200 355654 164400
rect 356426 163200 356482 164400
rect 357254 163200 357310 164400
rect 358082 163200 358138 164400
rect 358910 163200 358966 164400
rect 359738 163200 359794 164400
rect 360658 163200 360714 164400
rect 361486 163200 361542 164400
rect 362314 163200 362370 164400
rect 363142 163200 363198 164400
rect 363970 163200 364026 164400
rect 364798 163200 364854 164400
rect 365626 163200 365682 164400
rect 366454 163200 366510 164400
rect 367374 163200 367430 164400
rect 368202 163200 368258 164400
rect 369030 163200 369086 164400
rect 369858 163200 369914 164400
rect 370686 163200 370742 164400
rect 371514 163200 371570 164400
rect 372342 163200 372398 164400
rect 373170 163200 373226 164400
rect 374090 163200 374146 164400
rect 374918 163200 374974 164400
rect 375746 163200 375802 164400
rect 376574 163200 376630 164400
rect 377402 163200 377458 164400
rect 378230 163200 378286 164400
rect 379058 163200 379114 164400
rect 379886 163200 379942 164400
rect 380806 163200 380862 164400
rect 381634 163200 381690 164400
rect 382462 163200 382518 164400
rect 383290 163200 383346 164400
rect 384118 163200 384174 164400
rect 384946 163200 385002 164400
rect 385774 163200 385830 164400
rect 386602 163200 386658 164400
rect 387522 163200 387578 164400
rect 388350 163200 388406 164400
rect 389178 163200 389234 164400
rect 390006 163200 390062 164400
rect 390834 163200 390890 164400
rect 391662 163200 391718 164400
rect 392490 163200 392546 164400
rect 393410 163200 393466 164400
rect 394238 163200 394294 164400
rect 395066 163200 395122 164400
rect 395894 163200 395950 164400
rect 396722 163200 396778 164400
rect 397550 163200 397606 164400
rect 398378 163200 398434 164400
rect 399206 163200 399262 164400
rect 400126 163200 400182 164400
rect 400954 163200 401010 164400
rect 401782 163200 401838 164400
rect 402610 163200 402666 164400
rect 403438 163200 403494 164400
rect 404266 163200 404322 164400
rect 405094 163200 405150 164400
rect 405922 163200 405978 164400
rect 406842 163200 406898 164400
rect 407670 163200 407726 164400
rect 408498 163200 408554 164400
rect 409326 163200 409382 164400
rect 410154 163200 410210 164400
rect 410982 163200 411038 164400
rect 411810 163200 411866 164400
rect 412638 163200 412694 164400
rect 413558 163200 413614 164400
rect 414386 163200 414442 164400
rect 415214 163200 415270 164400
rect 416042 163200 416098 164400
rect 416870 163200 416926 164400
rect 417698 163200 417754 164400
rect 418526 163200 418582 164400
rect 419354 163200 419410 164400
rect 420274 163200 420330 164400
rect 421102 163200 421158 164400
rect 421930 163200 421986 164400
rect 422758 163200 422814 164400
rect 423586 163200 423642 164400
rect 424414 163200 424470 164400
rect 425242 163200 425298 164400
rect 426162 163200 426218 164400
rect 426990 163200 427046 164400
rect 427818 163200 427874 164400
rect 428646 163200 428702 164400
rect 429474 163200 429530 164400
rect 430302 163200 430358 164400
rect 431130 163200 431186 164400
rect 431958 163200 432014 164400
rect 432878 163200 432934 164400
rect 433706 163200 433762 164400
rect 434534 163200 434590 164400
rect 435362 163200 435418 164400
rect 436190 163200 436246 164400
rect 437018 163200 437074 164400
rect 437846 163200 437902 164400
rect 438674 163200 438730 164400
rect 439594 163200 439650 164400
rect 440422 163200 440478 164400
rect 441250 163200 441306 164400
rect 442078 163200 442134 164400
rect 442906 163200 442962 164400
rect 443734 163200 443790 164400
rect 444562 163200 444618 164400
rect 445390 163200 445446 164400
rect 446310 163200 446366 164400
rect 447138 163200 447194 164400
rect 447966 163200 448022 164400
rect 448794 163200 448850 164400
rect 449622 163200 449678 164400
rect 450450 163200 450506 164400
rect 451278 163200 451334 164400
rect 452106 163200 452162 164400
rect 453026 163200 453082 164400
rect 453854 163200 453910 164400
rect 454682 163200 454738 164400
rect 455510 163200 455566 164400
rect 456338 163200 456394 164400
rect 457166 163200 457222 164400
rect 457994 163200 458050 164400
rect 458914 163200 458970 164400
rect 459742 163200 459798 164400
rect 460570 163200 460626 164400
rect 461398 163200 461454 164400
rect 462226 163200 462282 164400
rect 463054 163200 463110 164400
rect 463882 163200 463938 164400
rect 464710 163200 464766 164400
rect 465630 163200 465686 164400
rect 466458 163200 466514 164400
rect 467286 163200 467342 164400
rect 468114 163200 468170 164400
rect 468942 163200 468998 164400
rect 469770 163200 469826 164400
rect 470598 163200 470654 164400
rect 471426 163200 471482 164400
rect 472346 163200 472402 164400
rect 473174 163200 473230 164400
rect 474002 163200 474058 164400
rect 474830 163200 474886 164400
rect 475658 163200 475714 164400
rect 476486 163200 476542 164400
rect 477314 163200 477370 164400
rect 478142 163200 478198 164400
rect 479062 163200 479118 164400
rect 479890 163200 479946 164400
rect 480718 163200 480774 164400
rect 481546 163200 481602 164400
rect 482374 163200 482430 164400
rect 483202 163200 483258 164400
rect 484030 163200 484086 164400
rect 484858 163200 484914 164400
rect 485778 163200 485834 164400
rect 486606 163200 486662 164400
rect 487434 163200 487490 164400
rect 488262 163200 488318 164400
rect 489090 163200 489146 164400
rect 489918 163200 489974 164400
rect 490746 163200 490802 164400
rect 491666 163200 491722 164400
rect 492494 163200 492550 164400
rect 493322 163200 493378 164400
rect 494150 163200 494206 164400
rect 494978 163200 495034 164400
rect 495806 163200 495862 164400
rect 496634 163200 496690 164400
rect 497462 163200 497518 164400
rect 498382 163200 498438 164400
rect 499210 163200 499266 164400
rect 500038 163200 500094 164400
rect 500866 163200 500922 164400
rect 501694 163200 501750 164400
rect 502522 163200 502578 164400
rect 503350 163200 503406 164400
rect 504178 163200 504234 164400
rect 505098 163200 505154 164400
rect 505926 163200 505982 164400
rect 506754 163200 506810 164400
rect 507582 163200 507638 164400
rect 508410 163200 508466 164400
rect 509238 163200 509294 164400
rect 510066 163200 510122 164400
rect 510894 163200 510950 164400
rect 511814 163200 511870 164400
rect 512642 163200 512698 164400
rect 513470 163200 513526 164400
rect 514298 163200 514354 164400
rect 515126 163200 515182 164400
rect 515954 163200 516010 164400
rect 516782 163200 516838 164400
rect 517610 163200 517666 164400
rect 518530 163200 518586 164400
rect 519358 163200 519414 164400
rect 520186 163200 520242 164400
rect 521014 163200 521070 164400
rect 521842 163200 521898 164400
rect 522670 163200 522726 164400
rect 523498 163200 523554 164400
rect 32770 -400 32826 800
rect 98274 -400 98330 800
rect 163778 -400 163834 800
rect 229282 -400 229338 800
rect 294786 -400 294842 800
rect 360290 -400 360346 800
rect 425794 -400 425850 800
rect 491298 -400 491354 800
<< obsm2 >>
rect 498 163144 1158 163282
rect 1326 163144 1986 163282
rect 2154 163144 2814 163282
rect 2982 163144 3642 163282
rect 3810 163144 4470 163282
rect 4638 163144 5298 163282
rect 5466 163144 6126 163282
rect 6294 163144 7046 163282
rect 7214 163144 7874 163282
rect 8042 163144 8702 163282
rect 8870 163144 9530 163282
rect 9698 163144 10358 163282
rect 10526 163144 11186 163282
rect 11354 163144 12014 163282
rect 12182 163144 12842 163282
rect 13010 163144 13762 163282
rect 13930 163144 14590 163282
rect 14758 163144 15418 163282
rect 15586 163144 16246 163282
rect 16414 163144 17074 163282
rect 17242 163144 17902 163282
rect 18070 163144 18730 163282
rect 18898 163144 19558 163282
rect 19726 163144 20478 163282
rect 20646 163144 21306 163282
rect 21474 163144 22134 163282
rect 22302 163144 22962 163282
rect 23130 163144 23790 163282
rect 23958 163144 24618 163282
rect 24786 163144 25446 163282
rect 25614 163144 26274 163282
rect 26442 163144 27194 163282
rect 27362 163144 28022 163282
rect 28190 163144 28850 163282
rect 29018 163144 29678 163282
rect 29846 163144 30506 163282
rect 30674 163144 31334 163282
rect 31502 163144 32162 163282
rect 32330 163144 33082 163282
rect 33250 163144 33910 163282
rect 34078 163144 34738 163282
rect 34906 163144 35566 163282
rect 35734 163144 36394 163282
rect 36562 163144 37222 163282
rect 37390 163144 38050 163282
rect 38218 163144 38878 163282
rect 39046 163144 39798 163282
rect 39966 163144 40626 163282
rect 40794 163144 41454 163282
rect 41622 163144 42282 163282
rect 42450 163144 43110 163282
rect 43278 163144 43938 163282
rect 44106 163144 44766 163282
rect 44934 163144 45594 163282
rect 45762 163144 46514 163282
rect 46682 163144 47342 163282
rect 47510 163144 48170 163282
rect 48338 163144 48998 163282
rect 49166 163144 49826 163282
rect 49994 163144 50654 163282
rect 50822 163144 51482 163282
rect 51650 163144 52310 163282
rect 52478 163144 53230 163282
rect 53398 163144 54058 163282
rect 54226 163144 54886 163282
rect 55054 163144 55714 163282
rect 55882 163144 56542 163282
rect 56710 163144 57370 163282
rect 57538 163144 58198 163282
rect 58366 163144 59026 163282
rect 59194 163144 59946 163282
rect 60114 163144 60774 163282
rect 60942 163144 61602 163282
rect 61770 163144 62430 163282
rect 62598 163144 63258 163282
rect 63426 163144 64086 163282
rect 64254 163144 64914 163282
rect 65082 163144 65834 163282
rect 66002 163144 66662 163282
rect 66830 163144 67490 163282
rect 67658 163144 68318 163282
rect 68486 163144 69146 163282
rect 69314 163144 69974 163282
rect 70142 163144 70802 163282
rect 70970 163144 71630 163282
rect 71798 163144 72550 163282
rect 72718 163144 73378 163282
rect 73546 163144 74206 163282
rect 74374 163144 75034 163282
rect 75202 163144 75862 163282
rect 76030 163144 76690 163282
rect 76858 163144 77518 163282
rect 77686 163144 78346 163282
rect 78514 163144 79266 163282
rect 79434 163144 80094 163282
rect 80262 163144 80922 163282
rect 81090 163144 81750 163282
rect 81918 163144 82578 163282
rect 82746 163144 83406 163282
rect 83574 163144 84234 163282
rect 84402 163144 85062 163282
rect 85230 163144 85982 163282
rect 86150 163144 86810 163282
rect 86978 163144 87638 163282
rect 87806 163144 88466 163282
rect 88634 163144 89294 163282
rect 89462 163144 90122 163282
rect 90290 163144 90950 163282
rect 91118 163144 91778 163282
rect 91946 163144 92698 163282
rect 92866 163144 93526 163282
rect 93694 163144 94354 163282
rect 94522 163144 95182 163282
rect 95350 163144 96010 163282
rect 96178 163144 96838 163282
rect 97006 163144 97666 163282
rect 97834 163144 98586 163282
rect 98754 163144 99414 163282
rect 99582 163144 100242 163282
rect 100410 163144 101070 163282
rect 101238 163144 101898 163282
rect 102066 163144 102726 163282
rect 102894 163144 103554 163282
rect 103722 163144 104382 163282
rect 104550 163144 105302 163282
rect 105470 163144 106130 163282
rect 106298 163144 106958 163282
rect 107126 163144 107786 163282
rect 107954 163144 108614 163282
rect 108782 163144 109442 163282
rect 109610 163144 110270 163282
rect 110438 163144 111098 163282
rect 111266 163144 112018 163282
rect 112186 163144 112846 163282
rect 113014 163144 113674 163282
rect 113842 163144 114502 163282
rect 114670 163144 115330 163282
rect 115498 163144 116158 163282
rect 116326 163144 116986 163282
rect 117154 163144 117814 163282
rect 117982 163144 118734 163282
rect 118902 163144 119562 163282
rect 119730 163144 120390 163282
rect 120558 163144 121218 163282
rect 121386 163144 122046 163282
rect 122214 163144 122874 163282
rect 123042 163144 123702 163282
rect 123870 163144 124530 163282
rect 124698 163144 125450 163282
rect 125618 163144 126278 163282
rect 126446 163144 127106 163282
rect 127274 163144 127934 163282
rect 128102 163144 128762 163282
rect 128930 163144 129590 163282
rect 129758 163144 130418 163282
rect 130586 163144 131338 163282
rect 131506 163144 132166 163282
rect 132334 163144 132994 163282
rect 133162 163144 133822 163282
rect 133990 163144 134650 163282
rect 134818 163144 135478 163282
rect 135646 163144 136306 163282
rect 136474 163144 137134 163282
rect 137302 163144 138054 163282
rect 138222 163144 138882 163282
rect 139050 163144 139710 163282
rect 139878 163144 140538 163282
rect 140706 163144 141366 163282
rect 141534 163144 142194 163282
rect 142362 163144 143022 163282
rect 143190 163144 143850 163282
rect 144018 163144 144770 163282
rect 144938 163144 145598 163282
rect 145766 163144 146426 163282
rect 146594 163144 147254 163282
rect 147422 163144 148082 163282
rect 148250 163144 148910 163282
rect 149078 163144 149738 163282
rect 149906 163144 150566 163282
rect 150734 163144 151486 163282
rect 151654 163144 152314 163282
rect 152482 163144 153142 163282
rect 153310 163144 153970 163282
rect 154138 163144 154798 163282
rect 154966 163144 155626 163282
rect 155794 163144 156454 163282
rect 156622 163144 157282 163282
rect 157450 163144 158202 163282
rect 158370 163144 159030 163282
rect 159198 163144 159858 163282
rect 160026 163144 160686 163282
rect 160854 163144 161514 163282
rect 161682 163144 162342 163282
rect 162510 163144 163170 163282
rect 163338 163144 164090 163282
rect 164258 163144 164918 163282
rect 165086 163144 165746 163282
rect 165914 163144 166574 163282
rect 166742 163144 167402 163282
rect 167570 163144 168230 163282
rect 168398 163144 169058 163282
rect 169226 163144 169886 163282
rect 170054 163144 170806 163282
rect 170974 163144 171634 163282
rect 171802 163144 172462 163282
rect 172630 163144 173290 163282
rect 173458 163144 174118 163282
rect 174286 163144 174946 163282
rect 175114 163144 175774 163282
rect 175942 163144 176602 163282
rect 176770 163144 177522 163282
rect 177690 163144 178350 163282
rect 178518 163144 179178 163282
rect 179346 163144 180006 163282
rect 180174 163144 180834 163282
rect 181002 163144 181662 163282
rect 181830 163144 182490 163282
rect 182658 163144 183318 163282
rect 183486 163144 184238 163282
rect 184406 163144 185066 163282
rect 185234 163144 185894 163282
rect 186062 163144 186722 163282
rect 186890 163144 187550 163282
rect 187718 163144 188378 163282
rect 188546 163144 189206 163282
rect 189374 163144 190034 163282
rect 190202 163144 190954 163282
rect 191122 163144 191782 163282
rect 191950 163144 192610 163282
rect 192778 163144 193438 163282
rect 193606 163144 194266 163282
rect 194434 163144 195094 163282
rect 195262 163144 195922 163282
rect 196090 163144 196842 163282
rect 197010 163144 197670 163282
rect 197838 163144 198498 163282
rect 198666 163144 199326 163282
rect 199494 163144 200154 163282
rect 200322 163144 200982 163282
rect 201150 163144 201810 163282
rect 201978 163144 202638 163282
rect 202806 163144 203558 163282
rect 203726 163144 204386 163282
rect 204554 163144 205214 163282
rect 205382 163144 206042 163282
rect 206210 163144 206870 163282
rect 207038 163144 207698 163282
rect 207866 163144 208526 163282
rect 208694 163144 209354 163282
rect 209522 163144 210274 163282
rect 210442 163144 211102 163282
rect 211270 163144 211930 163282
rect 212098 163144 212758 163282
rect 212926 163144 213586 163282
rect 213754 163144 214414 163282
rect 214582 163144 215242 163282
rect 215410 163144 216070 163282
rect 216238 163144 216990 163282
rect 217158 163144 217818 163282
rect 217986 163144 218646 163282
rect 218814 163144 219474 163282
rect 219642 163144 220302 163282
rect 220470 163144 221130 163282
rect 221298 163144 221958 163282
rect 222126 163144 222786 163282
rect 222954 163144 223706 163282
rect 223874 163144 224534 163282
rect 224702 163144 225362 163282
rect 225530 163144 226190 163282
rect 226358 163144 227018 163282
rect 227186 163144 227846 163282
rect 228014 163144 228674 163282
rect 228842 163144 229594 163282
rect 229762 163144 230422 163282
rect 230590 163144 231250 163282
rect 231418 163144 232078 163282
rect 232246 163144 232906 163282
rect 233074 163144 233734 163282
rect 233902 163144 234562 163282
rect 234730 163144 235390 163282
rect 235558 163144 236310 163282
rect 236478 163144 237138 163282
rect 237306 163144 237966 163282
rect 238134 163144 238794 163282
rect 238962 163144 239622 163282
rect 239790 163144 240450 163282
rect 240618 163144 241278 163282
rect 241446 163144 242106 163282
rect 242274 163144 243026 163282
rect 243194 163144 243854 163282
rect 244022 163144 244682 163282
rect 244850 163144 245510 163282
rect 245678 163144 246338 163282
rect 246506 163144 247166 163282
rect 247334 163144 247994 163282
rect 248162 163144 248822 163282
rect 248990 163144 249742 163282
rect 249910 163144 250570 163282
rect 250738 163144 251398 163282
rect 251566 163144 252226 163282
rect 252394 163144 253054 163282
rect 253222 163144 253882 163282
rect 254050 163144 254710 163282
rect 254878 163144 255538 163282
rect 255706 163144 256458 163282
rect 256626 163144 257286 163282
rect 257454 163144 258114 163282
rect 258282 163144 258942 163282
rect 259110 163144 259770 163282
rect 259938 163144 260598 163282
rect 260766 163144 261426 163282
rect 261594 163144 262346 163282
rect 262514 163144 263174 163282
rect 263342 163144 264002 163282
rect 264170 163144 264830 163282
rect 264998 163144 265658 163282
rect 265826 163144 266486 163282
rect 266654 163144 267314 163282
rect 267482 163144 268142 163282
rect 268310 163144 269062 163282
rect 269230 163144 269890 163282
rect 270058 163144 270718 163282
rect 270886 163144 271546 163282
rect 271714 163144 272374 163282
rect 272542 163144 273202 163282
rect 273370 163144 274030 163282
rect 274198 163144 274858 163282
rect 275026 163144 275778 163282
rect 275946 163144 276606 163282
rect 276774 163144 277434 163282
rect 277602 163144 278262 163282
rect 278430 163144 279090 163282
rect 279258 163144 279918 163282
rect 280086 163144 280746 163282
rect 280914 163144 281574 163282
rect 281742 163144 282494 163282
rect 282662 163144 283322 163282
rect 283490 163144 284150 163282
rect 284318 163144 284978 163282
rect 285146 163144 285806 163282
rect 285974 163144 286634 163282
rect 286802 163144 287462 163282
rect 287630 163144 288290 163282
rect 288458 163144 289210 163282
rect 289378 163144 290038 163282
rect 290206 163144 290866 163282
rect 291034 163144 291694 163282
rect 291862 163144 292522 163282
rect 292690 163144 293350 163282
rect 293518 163144 294178 163282
rect 294346 163144 295098 163282
rect 295266 163144 295926 163282
rect 296094 163144 296754 163282
rect 296922 163144 297582 163282
rect 297750 163144 298410 163282
rect 298578 163144 299238 163282
rect 299406 163144 300066 163282
rect 300234 163144 300894 163282
rect 301062 163144 301814 163282
rect 301982 163144 302642 163282
rect 302810 163144 303470 163282
rect 303638 163144 304298 163282
rect 304466 163144 305126 163282
rect 305294 163144 305954 163282
rect 306122 163144 306782 163282
rect 306950 163144 307610 163282
rect 307778 163144 308530 163282
rect 308698 163144 309358 163282
rect 309526 163144 310186 163282
rect 310354 163144 311014 163282
rect 311182 163144 311842 163282
rect 312010 163144 312670 163282
rect 312838 163144 313498 163282
rect 313666 163144 314326 163282
rect 314494 163144 315246 163282
rect 315414 163144 316074 163282
rect 316242 163144 316902 163282
rect 317070 163144 317730 163282
rect 317898 163144 318558 163282
rect 318726 163144 319386 163282
rect 319554 163144 320214 163282
rect 320382 163144 321042 163282
rect 321210 163144 321962 163282
rect 322130 163144 322790 163282
rect 322958 163144 323618 163282
rect 323786 163144 324446 163282
rect 324614 163144 325274 163282
rect 325442 163144 326102 163282
rect 326270 163144 326930 163282
rect 327098 163144 327850 163282
rect 328018 163144 328678 163282
rect 328846 163144 329506 163282
rect 329674 163144 330334 163282
rect 330502 163144 331162 163282
rect 331330 163144 331990 163282
rect 332158 163144 332818 163282
rect 332986 163144 333646 163282
rect 333814 163144 334566 163282
rect 334734 163144 335394 163282
rect 335562 163144 336222 163282
rect 336390 163144 337050 163282
rect 337218 163144 337878 163282
rect 338046 163144 338706 163282
rect 338874 163144 339534 163282
rect 339702 163144 340362 163282
rect 340530 163144 341282 163282
rect 341450 163144 342110 163282
rect 342278 163144 342938 163282
rect 343106 163144 343766 163282
rect 343934 163144 344594 163282
rect 344762 163144 345422 163282
rect 345590 163144 346250 163282
rect 346418 163144 347078 163282
rect 347246 163144 347998 163282
rect 348166 163144 348826 163282
rect 348994 163144 349654 163282
rect 349822 163144 350482 163282
rect 350650 163144 351310 163282
rect 351478 163144 352138 163282
rect 352306 163144 352966 163282
rect 353134 163144 353794 163282
rect 353962 163144 354714 163282
rect 354882 163144 355542 163282
rect 355710 163144 356370 163282
rect 356538 163144 357198 163282
rect 357366 163144 358026 163282
rect 358194 163144 358854 163282
rect 359022 163144 359682 163282
rect 359850 163144 360602 163282
rect 360770 163144 361430 163282
rect 361598 163144 362258 163282
rect 362426 163144 363086 163282
rect 363254 163144 363914 163282
rect 364082 163144 364742 163282
rect 364910 163144 365570 163282
rect 365738 163144 366398 163282
rect 366566 163144 367318 163282
rect 367486 163144 368146 163282
rect 368314 163144 368974 163282
rect 369142 163144 369802 163282
rect 369970 163144 370630 163282
rect 370798 163144 371458 163282
rect 371626 163144 372286 163282
rect 372454 163144 373114 163282
rect 373282 163144 374034 163282
rect 374202 163144 374862 163282
rect 375030 163144 375690 163282
rect 375858 163144 376518 163282
rect 376686 163144 377346 163282
rect 377514 163144 378174 163282
rect 378342 163144 379002 163282
rect 379170 163144 379830 163282
rect 379998 163144 380750 163282
rect 380918 163144 381578 163282
rect 381746 163144 382406 163282
rect 382574 163144 383234 163282
rect 383402 163144 384062 163282
rect 384230 163144 384890 163282
rect 385058 163144 385718 163282
rect 385886 163144 386546 163282
rect 386714 163144 387466 163282
rect 387634 163144 388294 163282
rect 388462 163144 389122 163282
rect 389290 163144 389950 163282
rect 390118 163144 390778 163282
rect 390946 163144 391606 163282
rect 391774 163144 392434 163282
rect 392602 163144 393354 163282
rect 393522 163144 394182 163282
rect 394350 163144 395010 163282
rect 395178 163144 395838 163282
rect 396006 163144 396666 163282
rect 396834 163144 397494 163282
rect 397662 163144 398322 163282
rect 398490 163144 399150 163282
rect 399318 163144 400070 163282
rect 400238 163144 400898 163282
rect 401066 163144 401726 163282
rect 401894 163144 402554 163282
rect 402722 163144 403382 163282
rect 403550 163144 404210 163282
rect 404378 163144 405038 163282
rect 405206 163144 405866 163282
rect 406034 163144 406786 163282
rect 406954 163144 407614 163282
rect 407782 163144 408442 163282
rect 408610 163144 409270 163282
rect 409438 163144 410098 163282
rect 410266 163144 410926 163282
rect 411094 163144 411754 163282
rect 411922 163144 412582 163282
rect 412750 163144 413502 163282
rect 413670 163144 414330 163282
rect 414498 163144 415158 163282
rect 415326 163144 415986 163282
rect 416154 163144 416814 163282
rect 416982 163144 417642 163282
rect 417810 163144 418470 163282
rect 418638 163144 419298 163282
rect 419466 163144 420218 163282
rect 420386 163144 421046 163282
rect 421214 163144 421874 163282
rect 422042 163144 422702 163282
rect 422870 163144 423530 163282
rect 423698 163144 424358 163282
rect 424526 163144 425186 163282
rect 425354 163144 426106 163282
rect 426274 163144 426934 163282
rect 427102 163144 427762 163282
rect 427930 163144 428590 163282
rect 428758 163144 429418 163282
rect 429586 163144 430246 163282
rect 430414 163144 431074 163282
rect 431242 163144 431902 163282
rect 432070 163144 432822 163282
rect 432990 163144 433650 163282
rect 433818 163144 434478 163282
rect 434646 163144 435306 163282
rect 435474 163144 436134 163282
rect 436302 163144 436962 163282
rect 437130 163144 437790 163282
rect 437958 163144 438618 163282
rect 438786 163144 439538 163282
rect 439706 163144 440366 163282
rect 440534 163144 441194 163282
rect 441362 163144 442022 163282
rect 442190 163144 442850 163282
rect 443018 163144 443678 163282
rect 443846 163144 444506 163282
rect 444674 163144 445334 163282
rect 445502 163144 446254 163282
rect 446422 163144 447082 163282
rect 447250 163144 447910 163282
rect 448078 163144 448738 163282
rect 448906 163144 449566 163282
rect 449734 163144 450394 163282
rect 450562 163144 451222 163282
rect 451390 163144 452050 163282
rect 452218 163144 452970 163282
rect 453138 163144 453798 163282
rect 453966 163144 454626 163282
rect 454794 163144 455454 163282
rect 455622 163144 456282 163282
rect 456450 163144 457110 163282
rect 457278 163144 457938 163282
rect 458106 163144 458858 163282
rect 459026 163144 459686 163282
rect 459854 163144 460514 163282
rect 460682 163144 461342 163282
rect 461510 163144 462170 163282
rect 462338 163144 462998 163282
rect 463166 163144 463826 163282
rect 463994 163144 464654 163282
rect 464822 163144 465574 163282
rect 465742 163144 466402 163282
rect 466570 163144 467230 163282
rect 467398 163144 468058 163282
rect 468226 163144 468886 163282
rect 469054 163144 469714 163282
rect 469882 163144 470542 163282
rect 470710 163144 471370 163282
rect 471538 163144 472290 163282
rect 472458 163144 473118 163282
rect 473286 163144 473946 163282
rect 474114 163144 474774 163282
rect 474942 163144 475602 163282
rect 475770 163144 476430 163282
rect 476598 163144 477258 163282
rect 477426 163144 478086 163282
rect 478254 163144 479006 163282
rect 479174 163144 479834 163282
rect 480002 163144 480662 163282
rect 480830 163144 481490 163282
rect 481658 163144 482318 163282
rect 482486 163144 483146 163282
rect 483314 163144 483974 163282
rect 484142 163144 484802 163282
rect 484970 163144 485722 163282
rect 485890 163144 486550 163282
rect 486718 163144 487378 163282
rect 487546 163144 488206 163282
rect 488374 163144 489034 163282
rect 489202 163144 489862 163282
rect 490030 163144 490690 163282
rect 490858 163144 491610 163282
rect 491778 163144 492438 163282
rect 492606 163144 493266 163282
rect 493434 163144 494094 163282
rect 494262 163144 494922 163282
rect 495090 163144 495750 163282
rect 495918 163144 496578 163282
rect 496746 163144 497406 163282
rect 497574 163144 498326 163282
rect 498494 163144 499154 163282
rect 499322 163144 499982 163282
rect 500150 163144 500810 163282
rect 500978 163144 501638 163282
rect 501806 163144 502466 163282
rect 502634 163144 503294 163282
rect 503462 163144 504122 163282
rect 504290 163144 505042 163282
rect 505210 163144 505870 163282
rect 506038 163144 506698 163282
rect 506866 163144 507526 163282
rect 507694 163144 508354 163282
rect 508522 163144 509182 163282
rect 509350 163144 510010 163282
rect 510178 163144 510838 163282
rect 511006 163144 511758 163282
rect 511926 163144 512586 163282
rect 512754 163144 513414 163282
rect 513582 163144 514242 163282
rect 514410 163144 515070 163282
rect 515238 163144 515898 163282
rect 516066 163144 516726 163282
rect 516894 163144 517554 163282
rect 517722 163144 518474 163282
rect 518642 163144 519302 163282
rect 519470 163144 520130 163282
rect 520298 163144 520958 163282
rect 521126 163144 521786 163282
rect 521954 163144 522614 163282
rect 522782 163144 523442 163282
rect 388 856 523552 163144
rect 388 682 32714 856
rect 32882 682 98218 856
rect 98386 682 163722 856
rect 163890 682 229226 856
rect 229394 682 294730 856
rect 294898 682 360234 856
rect 360402 682 425738 856
rect 425906 682 491242 856
rect 491410 682 523552 856
<< metal3 >>
rect 523200 163072 524400 163192
rect 523200 161576 524400 161696
rect 523200 160080 524400 160200
rect 523200 158584 524400 158704
rect 523200 157088 524400 157208
rect 523200 155592 524400 155712
rect 523200 153960 524400 154080
rect 523200 152464 524400 152584
rect 523200 150968 524400 151088
rect 523200 149472 524400 149592
rect 523200 147976 524400 148096
rect 523200 146480 524400 146600
rect 523200 144848 524400 144968
rect 523200 143352 524400 143472
rect 523200 141856 524400 141976
rect 523200 140360 524400 140480
rect 523200 138864 524400 138984
rect 523200 137368 524400 137488
rect 523200 135736 524400 135856
rect 523200 134240 524400 134360
rect 523200 132744 524400 132864
rect 523200 131248 524400 131368
rect 523200 129752 524400 129872
rect 523200 128256 524400 128376
rect 523200 126624 524400 126744
rect 523200 125128 524400 125248
rect 523200 123632 524400 123752
rect 523200 122136 524400 122256
rect 523200 120640 524400 120760
rect 523200 119144 524400 119264
rect 523200 117512 524400 117632
rect 523200 116016 524400 116136
rect 523200 114520 524400 114640
rect 523200 113024 524400 113144
rect 523200 111528 524400 111648
rect 523200 110032 524400 110152
rect 523200 108400 524400 108520
rect 523200 106904 524400 107024
rect 523200 105408 524400 105528
rect 523200 103912 524400 104032
rect 523200 102416 524400 102536
rect 523200 100920 524400 101040
rect 523200 99288 524400 99408
rect 523200 97792 524400 97912
rect 523200 96296 524400 96416
rect 523200 94800 524400 94920
rect 523200 93304 524400 93424
rect 523200 91808 524400 91928
rect 523200 90176 524400 90296
rect 523200 88680 524400 88800
rect 523200 87184 524400 87304
rect 523200 85688 524400 85808
rect 523200 84192 524400 84312
rect 523200 82696 524400 82816
rect 523200 81064 524400 81184
rect 523200 79568 524400 79688
rect 523200 78072 524400 78192
rect 523200 76576 524400 76696
rect 523200 75080 524400 75200
rect 523200 73584 524400 73704
rect 523200 71952 524400 72072
rect 523200 70456 524400 70576
rect 523200 68960 524400 69080
rect 523200 67464 524400 67584
rect 523200 65968 524400 66088
rect 523200 64472 524400 64592
rect 523200 62840 524400 62960
rect 523200 61344 524400 61464
rect 523200 59848 524400 59968
rect 523200 58352 524400 58472
rect 523200 56856 524400 56976
rect 523200 55360 524400 55480
rect 523200 53728 524400 53848
rect 523200 52232 524400 52352
rect 523200 50736 524400 50856
rect 523200 49240 524400 49360
rect 523200 47744 524400 47864
rect 523200 46248 524400 46368
rect 523200 44616 524400 44736
rect 523200 43120 524400 43240
rect 523200 41624 524400 41744
rect 523200 40128 524400 40248
rect 523200 38632 524400 38752
rect 523200 37136 524400 37256
rect 523200 35504 524400 35624
rect 523200 34008 524400 34128
rect 523200 32512 524400 32632
rect 523200 31016 524400 31136
rect 523200 29520 524400 29640
rect 523200 28024 524400 28144
rect 523200 26392 524400 26512
rect 523200 24896 524400 25016
rect 523200 23400 524400 23520
rect 523200 21904 524400 22024
rect 523200 20408 524400 20528
rect 523200 18912 524400 19032
rect 523200 17280 524400 17400
rect 523200 15784 524400 15904
rect 523200 14288 524400 14408
rect 523200 12792 524400 12912
rect 523200 11296 524400 11416
rect 523200 9800 524400 9920
rect 523200 8168 524400 8288
rect 523200 6672 524400 6792
rect 523200 5176 524400 5296
rect 523200 3680 524400 3800
rect 523200 2184 524400 2304
rect 523200 688 524400 808
<< obsm3 >>
rect 2669 162992 523120 163165
rect 2669 161776 523200 162992
rect 2669 161496 523120 161776
rect 2669 160280 523200 161496
rect 2669 160000 523120 160280
rect 2669 158784 523200 160000
rect 2669 158504 523120 158784
rect 2669 157288 523200 158504
rect 2669 157008 523120 157288
rect 2669 155792 523200 157008
rect 2669 155512 523120 155792
rect 2669 154160 523200 155512
rect 2669 153880 523120 154160
rect 2669 152664 523200 153880
rect 2669 152384 523120 152664
rect 2669 151168 523200 152384
rect 2669 150888 523120 151168
rect 2669 149672 523200 150888
rect 2669 149392 523120 149672
rect 2669 148176 523200 149392
rect 2669 147896 523120 148176
rect 2669 146680 523200 147896
rect 2669 146400 523120 146680
rect 2669 145048 523200 146400
rect 2669 144768 523120 145048
rect 2669 143552 523200 144768
rect 2669 143272 523120 143552
rect 2669 142056 523200 143272
rect 2669 141776 523120 142056
rect 2669 140560 523200 141776
rect 2669 140280 523120 140560
rect 2669 139064 523200 140280
rect 2669 138784 523120 139064
rect 2669 137568 523200 138784
rect 2669 137288 523120 137568
rect 2669 135936 523200 137288
rect 2669 135656 523120 135936
rect 2669 134440 523200 135656
rect 2669 134160 523120 134440
rect 2669 132944 523200 134160
rect 2669 132664 523120 132944
rect 2669 131448 523200 132664
rect 2669 131168 523120 131448
rect 2669 129952 523200 131168
rect 2669 129672 523120 129952
rect 2669 128456 523200 129672
rect 2669 128176 523120 128456
rect 2669 126824 523200 128176
rect 2669 126544 523120 126824
rect 2669 125328 523200 126544
rect 2669 125048 523120 125328
rect 2669 123832 523200 125048
rect 2669 123552 523120 123832
rect 2669 122336 523200 123552
rect 2669 122056 523120 122336
rect 2669 120840 523200 122056
rect 2669 120560 523120 120840
rect 2669 119344 523200 120560
rect 2669 119064 523120 119344
rect 2669 117712 523200 119064
rect 2669 117432 523120 117712
rect 2669 116216 523200 117432
rect 2669 115936 523120 116216
rect 2669 114720 523200 115936
rect 2669 114440 523120 114720
rect 2669 113224 523200 114440
rect 2669 112944 523120 113224
rect 2669 111728 523200 112944
rect 2669 111448 523120 111728
rect 2669 110232 523200 111448
rect 2669 109952 523120 110232
rect 2669 108600 523200 109952
rect 2669 108320 523120 108600
rect 2669 107104 523200 108320
rect 2669 106824 523120 107104
rect 2669 105608 523200 106824
rect 2669 105328 523120 105608
rect 2669 104112 523200 105328
rect 2669 103832 523120 104112
rect 2669 102616 523200 103832
rect 2669 102336 523120 102616
rect 2669 101120 523200 102336
rect 2669 100840 523120 101120
rect 2669 99488 523200 100840
rect 2669 99208 523120 99488
rect 2669 97992 523200 99208
rect 2669 97712 523120 97992
rect 2669 96496 523200 97712
rect 2669 96216 523120 96496
rect 2669 95000 523200 96216
rect 2669 94720 523120 95000
rect 2669 93504 523200 94720
rect 2669 93224 523120 93504
rect 2669 92008 523200 93224
rect 2669 91728 523120 92008
rect 2669 90376 523200 91728
rect 2669 90096 523120 90376
rect 2669 88880 523200 90096
rect 2669 88600 523120 88880
rect 2669 87384 523200 88600
rect 2669 87104 523120 87384
rect 2669 85888 523200 87104
rect 2669 85608 523120 85888
rect 2669 84392 523200 85608
rect 2669 84112 523120 84392
rect 2669 82896 523200 84112
rect 2669 82616 523120 82896
rect 2669 81264 523200 82616
rect 2669 80984 523120 81264
rect 2669 79768 523200 80984
rect 2669 79488 523120 79768
rect 2669 78272 523200 79488
rect 2669 77992 523120 78272
rect 2669 76776 523200 77992
rect 2669 76496 523120 76776
rect 2669 75280 523200 76496
rect 2669 75000 523120 75280
rect 2669 73784 523200 75000
rect 2669 73504 523120 73784
rect 2669 72152 523200 73504
rect 2669 71872 523120 72152
rect 2669 70656 523200 71872
rect 2669 70376 523120 70656
rect 2669 69160 523200 70376
rect 2669 68880 523120 69160
rect 2669 67664 523200 68880
rect 2669 67384 523120 67664
rect 2669 66168 523200 67384
rect 2669 65888 523120 66168
rect 2669 64672 523200 65888
rect 2669 64392 523120 64672
rect 2669 63040 523200 64392
rect 2669 62760 523120 63040
rect 2669 61544 523200 62760
rect 2669 61264 523120 61544
rect 2669 60048 523200 61264
rect 2669 59768 523120 60048
rect 2669 58552 523200 59768
rect 2669 58272 523120 58552
rect 2669 57056 523200 58272
rect 2669 56776 523120 57056
rect 2669 55560 523200 56776
rect 2669 55280 523120 55560
rect 2669 53928 523200 55280
rect 2669 53648 523120 53928
rect 2669 52432 523200 53648
rect 2669 52152 523120 52432
rect 2669 50936 523200 52152
rect 2669 50656 523120 50936
rect 2669 49440 523200 50656
rect 2669 49160 523120 49440
rect 2669 47944 523200 49160
rect 2669 47664 523120 47944
rect 2669 46448 523200 47664
rect 2669 46168 523120 46448
rect 2669 44816 523200 46168
rect 2669 44536 523120 44816
rect 2669 43320 523200 44536
rect 2669 43040 523120 43320
rect 2669 41824 523200 43040
rect 2669 41544 523120 41824
rect 2669 40328 523200 41544
rect 2669 40048 523120 40328
rect 2669 38832 523200 40048
rect 2669 38552 523120 38832
rect 2669 37336 523200 38552
rect 2669 37056 523120 37336
rect 2669 35704 523200 37056
rect 2669 35424 523120 35704
rect 2669 34208 523200 35424
rect 2669 33928 523120 34208
rect 2669 32712 523200 33928
rect 2669 32432 523120 32712
rect 2669 31216 523200 32432
rect 2669 30936 523120 31216
rect 2669 29720 523200 30936
rect 2669 29440 523120 29720
rect 2669 28224 523200 29440
rect 2669 27944 523120 28224
rect 2669 26592 523200 27944
rect 2669 26312 523120 26592
rect 2669 25096 523200 26312
rect 2669 24816 523120 25096
rect 2669 23600 523200 24816
rect 2669 23320 523120 23600
rect 2669 22104 523200 23320
rect 2669 21824 523120 22104
rect 2669 20608 523200 21824
rect 2669 20328 523120 20608
rect 2669 19112 523200 20328
rect 2669 18832 523120 19112
rect 2669 17480 523200 18832
rect 2669 17200 523120 17480
rect 2669 15984 523200 17200
rect 2669 15704 523120 15984
rect 2669 14488 523200 15704
rect 2669 14208 523120 14488
rect 2669 12992 523200 14208
rect 2669 12712 523120 12992
rect 2669 11496 523200 12712
rect 2669 11216 523120 11496
rect 2669 10000 523200 11216
rect 2669 9720 523120 10000
rect 2669 8368 523200 9720
rect 2669 8088 523120 8368
rect 2669 6872 523200 8088
rect 2669 6592 523120 6872
rect 2669 5376 523200 6592
rect 2669 5096 523120 5376
rect 2669 3880 523200 5096
rect 2669 3600 523120 3880
rect 2669 2384 523200 3600
rect 2669 2104 523120 2384
rect 2669 888 523200 2104
rect 2669 715 523120 888
<< obsm4 >>
rect 1004 1531 518920 149812
<< metal5 >>
rect 1104 156856 522836 157496
rect 1104 143856 2200 144496
rect 109800 143856 120200 144496
rect 517800 143856 522836 144496
rect 1104 130856 2200 131496
rect 109800 130856 120200 131496
rect 517800 130856 522836 131496
rect 1104 117856 2200 118496
rect 109800 117856 120200 118496
rect 517800 117856 522836 118496
rect 1104 104856 2200 105496
rect 109800 104856 120200 105496
rect 517800 104856 522836 105496
rect 1104 91856 2200 92496
rect 109800 91856 120200 92496
rect 517800 91856 522836 92496
rect 1104 78856 2200 79496
rect 109800 78856 120200 79496
rect 517800 78856 522836 79496
rect 1104 65856 2200 66496
rect 109800 65856 120200 66496
rect 517800 65856 522836 66496
rect 1104 52856 2200 53496
rect 109800 52856 120200 53496
rect 517800 52856 522836 53496
rect 1104 39856 2200 40496
rect 109800 39856 120200 40496
rect 517800 39856 522836 40496
rect 1104 26856 2200 27496
rect 109800 26856 120200 27496
rect 517800 26856 522836 27496
rect 1104 13856 2200 14496
rect 109800 13856 120200 14496
rect 517800 13856 522836 14496
<< obsm5 >>
rect 1004 144816 518920 149812
rect 2520 143536 109480 144816
rect 120520 143536 517480 144816
rect 1004 131816 518920 143536
rect 2520 130536 109480 131816
rect 120520 130536 517480 131816
rect 1004 118816 518920 130536
rect 2520 117536 109480 118816
rect 120520 117536 517480 118816
rect 1004 105816 518920 117536
rect 2520 104536 109480 105816
rect 120520 104536 517480 105816
rect 1004 92816 518920 104536
rect 2520 91536 109480 92816
rect 120520 91536 517480 92816
rect 1004 79816 518920 91536
rect 2520 78536 109480 79816
rect 120520 78536 517480 79816
rect 1004 66816 518920 78536
rect 2520 65536 109480 66816
rect 120520 65536 517480 66816
rect 1004 53816 518920 65536
rect 2520 52536 109480 53816
rect 120520 52536 517480 53816
rect 1004 40816 518920 52536
rect 2520 39536 109480 40816
rect 120520 39536 517480 40816
rect 1004 27816 518920 39536
rect 2520 26536 109480 27816
rect 120520 26536 517480 27816
rect 1004 14816 518920 26536
rect 2520 13536 109480 14816
rect 120520 13536 517480 14816
rect 1004 2156 518920 13536
<< labels >>
rlabel metal5 s 1104 26856 2200 27496 6 VGND
port 1 nsew ground input
rlabel metal5 s 109800 26856 120200 27496 6 VGND
port 1 nsew ground input
rlabel metal5 s 517800 26856 522836 27496 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 52856 2200 53496 6 VGND
port 1 nsew ground input
rlabel metal5 s 109800 52856 120200 53496 6 VGND
port 1 nsew ground input
rlabel metal5 s 517800 52856 522836 53496 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 78856 2200 79496 6 VGND
port 1 nsew ground input
rlabel metal5 s 109800 78856 120200 79496 6 VGND
port 1 nsew ground input
rlabel metal5 s 517800 78856 522836 79496 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 104856 2200 105496 6 VGND
port 1 nsew ground input
rlabel metal5 s 109800 104856 120200 105496 6 VGND
port 1 nsew ground input
rlabel metal5 s 517800 104856 522836 105496 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 130856 2200 131496 6 VGND
port 1 nsew ground input
rlabel metal5 s 109800 130856 120200 131496 6 VGND
port 1 nsew ground input
rlabel metal5 s 517800 130856 522836 131496 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 156856 522836 157496 6 VGND
port 1 nsew ground input
rlabel metal5 s 1104 13856 2200 14496 6 VPWR
port 2 nsew power input
rlabel metal5 s 109800 13856 120200 14496 6 VPWR
port 2 nsew power input
rlabel metal5 s 517800 13856 522836 14496 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 39856 2200 40496 6 VPWR
port 2 nsew power input
rlabel metal5 s 109800 39856 120200 40496 6 VPWR
port 2 nsew power input
rlabel metal5 s 517800 39856 522836 40496 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 65856 2200 66496 6 VPWR
port 2 nsew power input
rlabel metal5 s 109800 65856 120200 66496 6 VPWR
port 2 nsew power input
rlabel metal5 s 517800 65856 522836 66496 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 91856 2200 92496 6 VPWR
port 2 nsew power input
rlabel metal5 s 109800 91856 120200 92496 6 VPWR
port 2 nsew power input
rlabel metal5 s 517800 91856 522836 92496 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 117856 2200 118496 6 VPWR
port 2 nsew power input
rlabel metal5 s 109800 117856 120200 118496 6 VPWR
port 2 nsew power input
rlabel metal5 s 517800 117856 522836 118496 6 VPWR
port 2 nsew power input
rlabel metal5 s 1104 143856 2200 144496 6 VPWR
port 2 nsew power input
rlabel metal5 s 109800 143856 120200 144496 6 VPWR
port 2 nsew power input
rlabel metal5 s 517800 143856 522836 144496 6 VPWR
port 2 nsew power input
rlabel metal2 s 294786 -400 294842 800 6 core_clk
port 3 nsew signal input
rlabel metal2 s 98274 -400 98330 800 6 core_rstn
port 4 nsew signal input
rlabel metal3 s 523200 64472 524400 64592 6 debug_in
port 5 nsew signal input
rlabel metal3 s 523200 65968 524400 66088 6 debug_mode
port 6 nsew signal output
rlabel metal3 s 523200 67464 524400 67584 6 debug_oeb
port 7 nsew signal output
rlabel metal3 s 523200 68960 524400 69080 6 debug_out
port 8 nsew signal output
rlabel metal3 s 523200 144848 524400 144968 6 flash_clk
port 9 nsew signal output
rlabel metal3 s 523200 143352 524400 143472 6 flash_csb
port 10 nsew signal output
rlabel metal3 s 523200 146480 524400 146600 6 flash_io0_di
port 11 nsew signal input
rlabel metal3 s 523200 147976 524400 148096 6 flash_io0_do
port 12 nsew signal output
rlabel metal3 s 523200 149472 524400 149592 6 flash_io0_oeb
port 13 nsew signal output
rlabel metal3 s 523200 150968 524400 151088 6 flash_io1_di
port 14 nsew signal input
rlabel metal3 s 523200 152464 524400 152584 6 flash_io1_do
port 15 nsew signal output
rlabel metal3 s 523200 153960 524400 154080 6 flash_io1_oeb
port 16 nsew signal output
rlabel metal3 s 523200 155592 524400 155712 6 flash_io2_di
port 17 nsew signal input
rlabel metal3 s 523200 157088 524400 157208 6 flash_io2_do
port 18 nsew signal output
rlabel metal3 s 523200 158584 524400 158704 6 flash_io2_oeb
port 19 nsew signal output
rlabel metal3 s 523200 160080 524400 160200 6 flash_io3_di
port 20 nsew signal input
rlabel metal3 s 523200 161576 524400 161696 6 flash_io3_do
port 21 nsew signal output
rlabel metal3 s 523200 163072 524400 163192 6 flash_io3_oeb
port 22 nsew signal output
rlabel metal2 s 32770 -400 32826 800 6 gpio_in_pad
port 23 nsew signal input
rlabel metal2 s 163778 -400 163834 800 6 gpio_inenb_pad
port 24 nsew signal output
rlabel metal2 s 229282 -400 229338 800 6 gpio_mode0_pad
port 25 nsew signal output
rlabel metal2 s 360290 -400 360346 800 6 gpio_mode1_pad
port 26 nsew signal output
rlabel metal2 s 425794 -400 425850 800 6 gpio_out_pad
port 27 nsew signal output
rlabel metal2 s 491298 -400 491354 800 6 gpio_outenb_pad
port 28 nsew signal output
rlabel metal3 s 523200 91808 524400 91928 6 hk_ack_i
port 29 nsew signal input
rlabel metal2 s 523498 163200 523554 164400 6 hk_cyc_o
port 30 nsew signal output
rlabel metal3 s 523200 94800 524400 94920 6 hk_dat_i[0]
port 31 nsew signal input
rlabel metal3 s 523200 110032 524400 110152 6 hk_dat_i[10]
port 32 nsew signal input
rlabel metal3 s 523200 111528 524400 111648 6 hk_dat_i[11]
port 33 nsew signal input
rlabel metal3 s 523200 113024 524400 113144 6 hk_dat_i[12]
port 34 nsew signal input
rlabel metal3 s 523200 114520 524400 114640 6 hk_dat_i[13]
port 35 nsew signal input
rlabel metal3 s 523200 116016 524400 116136 6 hk_dat_i[14]
port 36 nsew signal input
rlabel metal3 s 523200 117512 524400 117632 6 hk_dat_i[15]
port 37 nsew signal input
rlabel metal3 s 523200 119144 524400 119264 6 hk_dat_i[16]
port 38 nsew signal input
rlabel metal3 s 523200 120640 524400 120760 6 hk_dat_i[17]
port 39 nsew signal input
rlabel metal3 s 523200 122136 524400 122256 6 hk_dat_i[18]
port 40 nsew signal input
rlabel metal3 s 523200 123632 524400 123752 6 hk_dat_i[19]
port 41 nsew signal input
rlabel metal3 s 523200 96296 524400 96416 6 hk_dat_i[1]
port 42 nsew signal input
rlabel metal3 s 523200 125128 524400 125248 6 hk_dat_i[20]
port 43 nsew signal input
rlabel metal3 s 523200 126624 524400 126744 6 hk_dat_i[21]
port 44 nsew signal input
rlabel metal3 s 523200 128256 524400 128376 6 hk_dat_i[22]
port 45 nsew signal input
rlabel metal3 s 523200 129752 524400 129872 6 hk_dat_i[23]
port 46 nsew signal input
rlabel metal3 s 523200 131248 524400 131368 6 hk_dat_i[24]
port 47 nsew signal input
rlabel metal3 s 523200 132744 524400 132864 6 hk_dat_i[25]
port 48 nsew signal input
rlabel metal3 s 523200 134240 524400 134360 6 hk_dat_i[26]
port 49 nsew signal input
rlabel metal3 s 523200 135736 524400 135856 6 hk_dat_i[27]
port 50 nsew signal input
rlabel metal3 s 523200 137368 524400 137488 6 hk_dat_i[28]
port 51 nsew signal input
rlabel metal3 s 523200 138864 524400 138984 6 hk_dat_i[29]
port 52 nsew signal input
rlabel metal3 s 523200 97792 524400 97912 6 hk_dat_i[2]
port 53 nsew signal input
rlabel metal3 s 523200 140360 524400 140480 6 hk_dat_i[30]
port 54 nsew signal input
rlabel metal3 s 523200 141856 524400 141976 6 hk_dat_i[31]
port 55 nsew signal input
rlabel metal3 s 523200 99288 524400 99408 6 hk_dat_i[3]
port 56 nsew signal input
rlabel metal3 s 523200 100920 524400 101040 6 hk_dat_i[4]
port 57 nsew signal input
rlabel metal3 s 523200 102416 524400 102536 6 hk_dat_i[5]
port 58 nsew signal input
rlabel metal3 s 523200 103912 524400 104032 6 hk_dat_i[6]
port 59 nsew signal input
rlabel metal3 s 523200 105408 524400 105528 6 hk_dat_i[7]
port 60 nsew signal input
rlabel metal3 s 523200 106904 524400 107024 6 hk_dat_i[8]
port 61 nsew signal input
rlabel metal3 s 523200 108400 524400 108520 6 hk_dat_i[9]
port 62 nsew signal input
rlabel metal3 s 523200 93304 524400 93424 6 hk_stb_o
port 63 nsew signal output
rlabel metal2 s 521014 163200 521070 164400 6 irq[0]
port 64 nsew signal input
rlabel metal2 s 521842 163200 521898 164400 6 irq[1]
port 65 nsew signal input
rlabel metal2 s 522670 163200 522726 164400 6 irq[2]
port 66 nsew signal input
rlabel metal3 s 523200 75080 524400 75200 6 irq[3]
port 67 nsew signal input
rlabel metal3 s 523200 73584 524400 73704 6 irq[4]
port 68 nsew signal input
rlabel metal3 s 523200 71952 524400 72072 6 irq[5]
port 69 nsew signal input
rlabel metal2 s 386 163200 442 164400 6 la_iena[0]
port 70 nsew signal output
rlabel metal2 s 336278 163200 336334 164400 6 la_iena[100]
port 71 nsew signal output
rlabel metal2 s 339590 163200 339646 164400 6 la_iena[101]
port 72 nsew signal output
rlabel metal2 s 342994 163200 343050 164400 6 la_iena[102]
port 73 nsew signal output
rlabel metal2 s 346306 163200 346362 164400 6 la_iena[103]
port 74 nsew signal output
rlabel metal2 s 349710 163200 349766 164400 6 la_iena[104]
port 75 nsew signal output
rlabel metal2 s 353022 163200 353078 164400 6 la_iena[105]
port 76 nsew signal output
rlabel metal2 s 356426 163200 356482 164400 6 la_iena[106]
port 77 nsew signal output
rlabel metal2 s 359738 163200 359794 164400 6 la_iena[107]
port 78 nsew signal output
rlabel metal2 s 363142 163200 363198 164400 6 la_iena[108]
port 79 nsew signal output
rlabel metal2 s 366454 163200 366510 164400 6 la_iena[109]
port 80 nsew signal output
rlabel metal2 s 33966 163200 34022 164400 6 la_iena[10]
port 81 nsew signal output
rlabel metal2 s 369858 163200 369914 164400 6 la_iena[110]
port 82 nsew signal output
rlabel metal2 s 373170 163200 373226 164400 6 la_iena[111]
port 83 nsew signal output
rlabel metal2 s 376574 163200 376630 164400 6 la_iena[112]
port 84 nsew signal output
rlabel metal2 s 379886 163200 379942 164400 6 la_iena[113]
port 85 nsew signal output
rlabel metal2 s 383290 163200 383346 164400 6 la_iena[114]
port 86 nsew signal output
rlabel metal2 s 386602 163200 386658 164400 6 la_iena[115]
port 87 nsew signal output
rlabel metal2 s 390006 163200 390062 164400 6 la_iena[116]
port 88 nsew signal output
rlabel metal2 s 393410 163200 393466 164400 6 la_iena[117]
port 89 nsew signal output
rlabel metal2 s 396722 163200 396778 164400 6 la_iena[118]
port 90 nsew signal output
rlabel metal2 s 400126 163200 400182 164400 6 la_iena[119]
port 91 nsew signal output
rlabel metal2 s 37278 163200 37334 164400 6 la_iena[11]
port 92 nsew signal output
rlabel metal2 s 403438 163200 403494 164400 6 la_iena[120]
port 93 nsew signal output
rlabel metal2 s 406842 163200 406898 164400 6 la_iena[121]
port 94 nsew signal output
rlabel metal2 s 410154 163200 410210 164400 6 la_iena[122]
port 95 nsew signal output
rlabel metal2 s 413558 163200 413614 164400 6 la_iena[123]
port 96 nsew signal output
rlabel metal2 s 416870 163200 416926 164400 6 la_iena[124]
port 97 nsew signal output
rlabel metal2 s 420274 163200 420330 164400 6 la_iena[125]
port 98 nsew signal output
rlabel metal2 s 423586 163200 423642 164400 6 la_iena[126]
port 99 nsew signal output
rlabel metal2 s 426990 163200 427046 164400 6 la_iena[127]
port 100 nsew signal output
rlabel metal2 s 40682 163200 40738 164400 6 la_iena[12]
port 101 nsew signal output
rlabel metal2 s 43994 163200 44050 164400 6 la_iena[13]
port 102 nsew signal output
rlabel metal2 s 47398 163200 47454 164400 6 la_iena[14]
port 103 nsew signal output
rlabel metal2 s 50710 163200 50766 164400 6 la_iena[15]
port 104 nsew signal output
rlabel metal2 s 54114 163200 54170 164400 6 la_iena[16]
port 105 nsew signal output
rlabel metal2 s 57426 163200 57482 164400 6 la_iena[17]
port 106 nsew signal output
rlabel metal2 s 60830 163200 60886 164400 6 la_iena[18]
port 107 nsew signal output
rlabel metal2 s 64142 163200 64198 164400 6 la_iena[19]
port 108 nsew signal output
rlabel metal2 s 3698 163200 3754 164400 6 la_iena[1]
port 109 nsew signal output
rlabel metal2 s 67546 163200 67602 164400 6 la_iena[20]
port 110 nsew signal output
rlabel metal2 s 70858 163200 70914 164400 6 la_iena[21]
port 111 nsew signal output
rlabel metal2 s 74262 163200 74318 164400 6 la_iena[22]
port 112 nsew signal output
rlabel metal2 s 77574 163200 77630 164400 6 la_iena[23]
port 113 nsew signal output
rlabel metal2 s 80978 163200 81034 164400 6 la_iena[24]
port 114 nsew signal output
rlabel metal2 s 84290 163200 84346 164400 6 la_iena[25]
port 115 nsew signal output
rlabel metal2 s 87694 163200 87750 164400 6 la_iena[26]
port 116 nsew signal output
rlabel metal2 s 91006 163200 91062 164400 6 la_iena[27]
port 117 nsew signal output
rlabel metal2 s 94410 163200 94466 164400 6 la_iena[28]
port 118 nsew signal output
rlabel metal2 s 97722 163200 97778 164400 6 la_iena[29]
port 119 nsew signal output
rlabel metal2 s 7102 163200 7158 164400 6 la_iena[2]
port 120 nsew signal output
rlabel metal2 s 101126 163200 101182 164400 6 la_iena[30]
port 121 nsew signal output
rlabel metal2 s 104438 163200 104494 164400 6 la_iena[31]
port 122 nsew signal output
rlabel metal2 s 107842 163200 107898 164400 6 la_iena[32]
port 123 nsew signal output
rlabel metal2 s 111154 163200 111210 164400 6 la_iena[33]
port 124 nsew signal output
rlabel metal2 s 114558 163200 114614 164400 6 la_iena[34]
port 125 nsew signal output
rlabel metal2 s 117870 163200 117926 164400 6 la_iena[35]
port 126 nsew signal output
rlabel metal2 s 121274 163200 121330 164400 6 la_iena[36]
port 127 nsew signal output
rlabel metal2 s 124586 163200 124642 164400 6 la_iena[37]
port 128 nsew signal output
rlabel metal2 s 127990 163200 128046 164400 6 la_iena[38]
port 129 nsew signal output
rlabel metal2 s 131394 163200 131450 164400 6 la_iena[39]
port 130 nsew signal output
rlabel metal2 s 10414 163200 10470 164400 6 la_iena[3]
port 131 nsew signal output
rlabel metal2 s 134706 163200 134762 164400 6 la_iena[40]
port 132 nsew signal output
rlabel metal2 s 138110 163200 138166 164400 6 la_iena[41]
port 133 nsew signal output
rlabel metal2 s 141422 163200 141478 164400 6 la_iena[42]
port 134 nsew signal output
rlabel metal2 s 144826 163200 144882 164400 6 la_iena[43]
port 135 nsew signal output
rlabel metal2 s 148138 163200 148194 164400 6 la_iena[44]
port 136 nsew signal output
rlabel metal2 s 151542 163200 151598 164400 6 la_iena[45]
port 137 nsew signal output
rlabel metal2 s 154854 163200 154910 164400 6 la_iena[46]
port 138 nsew signal output
rlabel metal2 s 158258 163200 158314 164400 6 la_iena[47]
port 139 nsew signal output
rlabel metal2 s 161570 163200 161626 164400 6 la_iena[48]
port 140 nsew signal output
rlabel metal2 s 164974 163200 165030 164400 6 la_iena[49]
port 141 nsew signal output
rlabel metal2 s 13818 163200 13874 164400 6 la_iena[4]
port 142 nsew signal output
rlabel metal2 s 168286 163200 168342 164400 6 la_iena[50]
port 143 nsew signal output
rlabel metal2 s 171690 163200 171746 164400 6 la_iena[51]
port 144 nsew signal output
rlabel metal2 s 175002 163200 175058 164400 6 la_iena[52]
port 145 nsew signal output
rlabel metal2 s 178406 163200 178462 164400 6 la_iena[53]
port 146 nsew signal output
rlabel metal2 s 181718 163200 181774 164400 6 la_iena[54]
port 147 nsew signal output
rlabel metal2 s 185122 163200 185178 164400 6 la_iena[55]
port 148 nsew signal output
rlabel metal2 s 188434 163200 188490 164400 6 la_iena[56]
port 149 nsew signal output
rlabel metal2 s 191838 163200 191894 164400 6 la_iena[57]
port 150 nsew signal output
rlabel metal2 s 195150 163200 195206 164400 6 la_iena[58]
port 151 nsew signal output
rlabel metal2 s 198554 163200 198610 164400 6 la_iena[59]
port 152 nsew signal output
rlabel metal2 s 17130 163200 17186 164400 6 la_iena[5]
port 153 nsew signal output
rlabel metal2 s 201866 163200 201922 164400 6 la_iena[60]
port 154 nsew signal output
rlabel metal2 s 205270 163200 205326 164400 6 la_iena[61]
port 155 nsew signal output
rlabel metal2 s 208582 163200 208638 164400 6 la_iena[62]
port 156 nsew signal output
rlabel metal2 s 211986 163200 212042 164400 6 la_iena[63]
port 157 nsew signal output
rlabel metal2 s 215298 163200 215354 164400 6 la_iena[64]
port 158 nsew signal output
rlabel metal2 s 218702 163200 218758 164400 6 la_iena[65]
port 159 nsew signal output
rlabel metal2 s 222014 163200 222070 164400 6 la_iena[66]
port 160 nsew signal output
rlabel metal2 s 225418 163200 225474 164400 6 la_iena[67]
port 161 nsew signal output
rlabel metal2 s 228730 163200 228786 164400 6 la_iena[68]
port 162 nsew signal output
rlabel metal2 s 232134 163200 232190 164400 6 la_iena[69]
port 163 nsew signal output
rlabel metal2 s 20534 163200 20590 164400 6 la_iena[6]
port 164 nsew signal output
rlabel metal2 s 235446 163200 235502 164400 6 la_iena[70]
port 165 nsew signal output
rlabel metal2 s 238850 163200 238906 164400 6 la_iena[71]
port 166 nsew signal output
rlabel metal2 s 242162 163200 242218 164400 6 la_iena[72]
port 167 nsew signal output
rlabel metal2 s 245566 163200 245622 164400 6 la_iena[73]
port 168 nsew signal output
rlabel metal2 s 248878 163200 248934 164400 6 la_iena[74]
port 169 nsew signal output
rlabel metal2 s 252282 163200 252338 164400 6 la_iena[75]
port 170 nsew signal output
rlabel metal2 s 255594 163200 255650 164400 6 la_iena[76]
port 171 nsew signal output
rlabel metal2 s 258998 163200 259054 164400 6 la_iena[77]
port 172 nsew signal output
rlabel metal2 s 262402 163200 262458 164400 6 la_iena[78]
port 173 nsew signal output
rlabel metal2 s 265714 163200 265770 164400 6 la_iena[79]
port 174 nsew signal output
rlabel metal2 s 23846 163200 23902 164400 6 la_iena[7]
port 175 nsew signal output
rlabel metal2 s 269118 163200 269174 164400 6 la_iena[80]
port 176 nsew signal output
rlabel metal2 s 272430 163200 272486 164400 6 la_iena[81]
port 177 nsew signal output
rlabel metal2 s 275834 163200 275890 164400 6 la_iena[82]
port 178 nsew signal output
rlabel metal2 s 279146 163200 279202 164400 6 la_iena[83]
port 179 nsew signal output
rlabel metal2 s 282550 163200 282606 164400 6 la_iena[84]
port 180 nsew signal output
rlabel metal2 s 285862 163200 285918 164400 6 la_iena[85]
port 181 nsew signal output
rlabel metal2 s 289266 163200 289322 164400 6 la_iena[86]
port 182 nsew signal output
rlabel metal2 s 292578 163200 292634 164400 6 la_iena[87]
port 183 nsew signal output
rlabel metal2 s 295982 163200 296038 164400 6 la_iena[88]
port 184 nsew signal output
rlabel metal2 s 299294 163200 299350 164400 6 la_iena[89]
port 185 nsew signal output
rlabel metal2 s 27250 163200 27306 164400 6 la_iena[8]
port 186 nsew signal output
rlabel metal2 s 302698 163200 302754 164400 6 la_iena[90]
port 187 nsew signal output
rlabel metal2 s 306010 163200 306066 164400 6 la_iena[91]
port 188 nsew signal output
rlabel metal2 s 309414 163200 309470 164400 6 la_iena[92]
port 189 nsew signal output
rlabel metal2 s 312726 163200 312782 164400 6 la_iena[93]
port 190 nsew signal output
rlabel metal2 s 316130 163200 316186 164400 6 la_iena[94]
port 191 nsew signal output
rlabel metal2 s 319442 163200 319498 164400 6 la_iena[95]
port 192 nsew signal output
rlabel metal2 s 322846 163200 322902 164400 6 la_iena[96]
port 193 nsew signal output
rlabel metal2 s 326158 163200 326214 164400 6 la_iena[97]
port 194 nsew signal output
rlabel metal2 s 329562 163200 329618 164400 6 la_iena[98]
port 195 nsew signal output
rlabel metal2 s 332874 163200 332930 164400 6 la_iena[99]
port 196 nsew signal output
rlabel metal2 s 30562 163200 30618 164400 6 la_iena[9]
port 197 nsew signal output
rlabel metal2 s 1214 163200 1270 164400 6 la_input[0]
port 198 nsew signal input
rlabel metal2 s 337106 163200 337162 164400 6 la_input[100]
port 199 nsew signal input
rlabel metal2 s 340418 163200 340474 164400 6 la_input[101]
port 200 nsew signal input
rlabel metal2 s 343822 163200 343878 164400 6 la_input[102]
port 201 nsew signal input
rlabel metal2 s 347134 163200 347190 164400 6 la_input[103]
port 202 nsew signal input
rlabel metal2 s 350538 163200 350594 164400 6 la_input[104]
port 203 nsew signal input
rlabel metal2 s 353850 163200 353906 164400 6 la_input[105]
port 204 nsew signal input
rlabel metal2 s 357254 163200 357310 164400 6 la_input[106]
port 205 nsew signal input
rlabel metal2 s 360658 163200 360714 164400 6 la_input[107]
port 206 nsew signal input
rlabel metal2 s 363970 163200 364026 164400 6 la_input[108]
port 207 nsew signal input
rlabel metal2 s 367374 163200 367430 164400 6 la_input[109]
port 208 nsew signal input
rlabel metal2 s 34794 163200 34850 164400 6 la_input[10]
port 209 nsew signal input
rlabel metal2 s 370686 163200 370742 164400 6 la_input[110]
port 210 nsew signal input
rlabel metal2 s 374090 163200 374146 164400 6 la_input[111]
port 211 nsew signal input
rlabel metal2 s 377402 163200 377458 164400 6 la_input[112]
port 212 nsew signal input
rlabel metal2 s 380806 163200 380862 164400 6 la_input[113]
port 213 nsew signal input
rlabel metal2 s 384118 163200 384174 164400 6 la_input[114]
port 214 nsew signal input
rlabel metal2 s 387522 163200 387578 164400 6 la_input[115]
port 215 nsew signal input
rlabel metal2 s 390834 163200 390890 164400 6 la_input[116]
port 216 nsew signal input
rlabel metal2 s 394238 163200 394294 164400 6 la_input[117]
port 217 nsew signal input
rlabel metal2 s 397550 163200 397606 164400 6 la_input[118]
port 218 nsew signal input
rlabel metal2 s 400954 163200 401010 164400 6 la_input[119]
port 219 nsew signal input
rlabel metal2 s 38106 163200 38162 164400 6 la_input[11]
port 220 nsew signal input
rlabel metal2 s 404266 163200 404322 164400 6 la_input[120]
port 221 nsew signal input
rlabel metal2 s 407670 163200 407726 164400 6 la_input[121]
port 222 nsew signal input
rlabel metal2 s 410982 163200 411038 164400 6 la_input[122]
port 223 nsew signal input
rlabel metal2 s 414386 163200 414442 164400 6 la_input[123]
port 224 nsew signal input
rlabel metal2 s 417698 163200 417754 164400 6 la_input[124]
port 225 nsew signal input
rlabel metal2 s 421102 163200 421158 164400 6 la_input[125]
port 226 nsew signal input
rlabel metal2 s 424414 163200 424470 164400 6 la_input[126]
port 227 nsew signal input
rlabel metal2 s 427818 163200 427874 164400 6 la_input[127]
port 228 nsew signal input
rlabel metal2 s 41510 163200 41566 164400 6 la_input[12]
port 229 nsew signal input
rlabel metal2 s 44822 163200 44878 164400 6 la_input[13]
port 230 nsew signal input
rlabel metal2 s 48226 163200 48282 164400 6 la_input[14]
port 231 nsew signal input
rlabel metal2 s 51538 163200 51594 164400 6 la_input[15]
port 232 nsew signal input
rlabel metal2 s 54942 163200 54998 164400 6 la_input[16]
port 233 nsew signal input
rlabel metal2 s 58254 163200 58310 164400 6 la_input[17]
port 234 nsew signal input
rlabel metal2 s 61658 163200 61714 164400 6 la_input[18]
port 235 nsew signal input
rlabel metal2 s 64970 163200 65026 164400 6 la_input[19]
port 236 nsew signal input
rlabel metal2 s 4526 163200 4582 164400 6 la_input[1]
port 237 nsew signal input
rlabel metal2 s 68374 163200 68430 164400 6 la_input[20]
port 238 nsew signal input
rlabel metal2 s 71686 163200 71742 164400 6 la_input[21]
port 239 nsew signal input
rlabel metal2 s 75090 163200 75146 164400 6 la_input[22]
port 240 nsew signal input
rlabel metal2 s 78402 163200 78458 164400 6 la_input[23]
port 241 nsew signal input
rlabel metal2 s 81806 163200 81862 164400 6 la_input[24]
port 242 nsew signal input
rlabel metal2 s 85118 163200 85174 164400 6 la_input[25]
port 243 nsew signal input
rlabel metal2 s 88522 163200 88578 164400 6 la_input[26]
port 244 nsew signal input
rlabel metal2 s 91834 163200 91890 164400 6 la_input[27]
port 245 nsew signal input
rlabel metal2 s 95238 163200 95294 164400 6 la_input[28]
port 246 nsew signal input
rlabel metal2 s 98642 163200 98698 164400 6 la_input[29]
port 247 nsew signal input
rlabel metal2 s 7930 163200 7986 164400 6 la_input[2]
port 248 nsew signal input
rlabel metal2 s 101954 163200 102010 164400 6 la_input[30]
port 249 nsew signal input
rlabel metal2 s 105358 163200 105414 164400 6 la_input[31]
port 250 nsew signal input
rlabel metal2 s 108670 163200 108726 164400 6 la_input[32]
port 251 nsew signal input
rlabel metal2 s 112074 163200 112130 164400 6 la_input[33]
port 252 nsew signal input
rlabel metal2 s 115386 163200 115442 164400 6 la_input[34]
port 253 nsew signal input
rlabel metal2 s 118790 163200 118846 164400 6 la_input[35]
port 254 nsew signal input
rlabel metal2 s 122102 163200 122158 164400 6 la_input[36]
port 255 nsew signal input
rlabel metal2 s 125506 163200 125562 164400 6 la_input[37]
port 256 nsew signal input
rlabel metal2 s 128818 163200 128874 164400 6 la_input[38]
port 257 nsew signal input
rlabel metal2 s 132222 163200 132278 164400 6 la_input[39]
port 258 nsew signal input
rlabel metal2 s 11242 163200 11298 164400 6 la_input[3]
port 259 nsew signal input
rlabel metal2 s 135534 163200 135590 164400 6 la_input[40]
port 260 nsew signal input
rlabel metal2 s 138938 163200 138994 164400 6 la_input[41]
port 261 nsew signal input
rlabel metal2 s 142250 163200 142306 164400 6 la_input[42]
port 262 nsew signal input
rlabel metal2 s 145654 163200 145710 164400 6 la_input[43]
port 263 nsew signal input
rlabel metal2 s 148966 163200 149022 164400 6 la_input[44]
port 264 nsew signal input
rlabel metal2 s 152370 163200 152426 164400 6 la_input[45]
port 265 nsew signal input
rlabel metal2 s 155682 163200 155738 164400 6 la_input[46]
port 266 nsew signal input
rlabel metal2 s 159086 163200 159142 164400 6 la_input[47]
port 267 nsew signal input
rlabel metal2 s 162398 163200 162454 164400 6 la_input[48]
port 268 nsew signal input
rlabel metal2 s 165802 163200 165858 164400 6 la_input[49]
port 269 nsew signal input
rlabel metal2 s 14646 163200 14702 164400 6 la_input[4]
port 270 nsew signal input
rlabel metal2 s 169114 163200 169170 164400 6 la_input[50]
port 271 nsew signal input
rlabel metal2 s 172518 163200 172574 164400 6 la_input[51]
port 272 nsew signal input
rlabel metal2 s 175830 163200 175886 164400 6 la_input[52]
port 273 nsew signal input
rlabel metal2 s 179234 163200 179290 164400 6 la_input[53]
port 274 nsew signal input
rlabel metal2 s 182546 163200 182602 164400 6 la_input[54]
port 275 nsew signal input
rlabel metal2 s 185950 163200 186006 164400 6 la_input[55]
port 276 nsew signal input
rlabel metal2 s 189262 163200 189318 164400 6 la_input[56]
port 277 nsew signal input
rlabel metal2 s 192666 163200 192722 164400 6 la_input[57]
port 278 nsew signal input
rlabel metal2 s 195978 163200 196034 164400 6 la_input[58]
port 279 nsew signal input
rlabel metal2 s 199382 163200 199438 164400 6 la_input[59]
port 280 nsew signal input
rlabel metal2 s 17958 163200 18014 164400 6 la_input[5]
port 281 nsew signal input
rlabel metal2 s 202694 163200 202750 164400 6 la_input[60]
port 282 nsew signal input
rlabel metal2 s 206098 163200 206154 164400 6 la_input[61]
port 283 nsew signal input
rlabel metal2 s 209410 163200 209466 164400 6 la_input[62]
port 284 nsew signal input
rlabel metal2 s 212814 163200 212870 164400 6 la_input[63]
port 285 nsew signal input
rlabel metal2 s 216126 163200 216182 164400 6 la_input[64]
port 286 nsew signal input
rlabel metal2 s 219530 163200 219586 164400 6 la_input[65]
port 287 nsew signal input
rlabel metal2 s 222842 163200 222898 164400 6 la_input[66]
port 288 nsew signal input
rlabel metal2 s 226246 163200 226302 164400 6 la_input[67]
port 289 nsew signal input
rlabel metal2 s 229650 163200 229706 164400 6 la_input[68]
port 290 nsew signal input
rlabel metal2 s 232962 163200 233018 164400 6 la_input[69]
port 291 nsew signal input
rlabel metal2 s 21362 163200 21418 164400 6 la_input[6]
port 292 nsew signal input
rlabel metal2 s 236366 163200 236422 164400 6 la_input[70]
port 293 nsew signal input
rlabel metal2 s 239678 163200 239734 164400 6 la_input[71]
port 294 nsew signal input
rlabel metal2 s 243082 163200 243138 164400 6 la_input[72]
port 295 nsew signal input
rlabel metal2 s 246394 163200 246450 164400 6 la_input[73]
port 296 nsew signal input
rlabel metal2 s 249798 163200 249854 164400 6 la_input[74]
port 297 nsew signal input
rlabel metal2 s 253110 163200 253166 164400 6 la_input[75]
port 298 nsew signal input
rlabel metal2 s 256514 163200 256570 164400 6 la_input[76]
port 299 nsew signal input
rlabel metal2 s 259826 163200 259882 164400 6 la_input[77]
port 300 nsew signal input
rlabel metal2 s 263230 163200 263286 164400 6 la_input[78]
port 301 nsew signal input
rlabel metal2 s 266542 163200 266598 164400 6 la_input[79]
port 302 nsew signal input
rlabel metal2 s 24674 163200 24730 164400 6 la_input[7]
port 303 nsew signal input
rlabel metal2 s 269946 163200 270002 164400 6 la_input[80]
port 304 nsew signal input
rlabel metal2 s 273258 163200 273314 164400 6 la_input[81]
port 305 nsew signal input
rlabel metal2 s 276662 163200 276718 164400 6 la_input[82]
port 306 nsew signal input
rlabel metal2 s 279974 163200 280030 164400 6 la_input[83]
port 307 nsew signal input
rlabel metal2 s 283378 163200 283434 164400 6 la_input[84]
port 308 nsew signal input
rlabel metal2 s 286690 163200 286746 164400 6 la_input[85]
port 309 nsew signal input
rlabel metal2 s 290094 163200 290150 164400 6 la_input[86]
port 310 nsew signal input
rlabel metal2 s 293406 163200 293462 164400 6 la_input[87]
port 311 nsew signal input
rlabel metal2 s 296810 163200 296866 164400 6 la_input[88]
port 312 nsew signal input
rlabel metal2 s 300122 163200 300178 164400 6 la_input[89]
port 313 nsew signal input
rlabel metal2 s 28078 163200 28134 164400 6 la_input[8]
port 314 nsew signal input
rlabel metal2 s 303526 163200 303582 164400 6 la_input[90]
port 315 nsew signal input
rlabel metal2 s 306838 163200 306894 164400 6 la_input[91]
port 316 nsew signal input
rlabel metal2 s 310242 163200 310298 164400 6 la_input[92]
port 317 nsew signal input
rlabel metal2 s 313554 163200 313610 164400 6 la_input[93]
port 318 nsew signal input
rlabel metal2 s 316958 163200 317014 164400 6 la_input[94]
port 319 nsew signal input
rlabel metal2 s 320270 163200 320326 164400 6 la_input[95]
port 320 nsew signal input
rlabel metal2 s 323674 163200 323730 164400 6 la_input[96]
port 321 nsew signal input
rlabel metal2 s 326986 163200 327042 164400 6 la_input[97]
port 322 nsew signal input
rlabel metal2 s 330390 163200 330446 164400 6 la_input[98]
port 323 nsew signal input
rlabel metal2 s 333702 163200 333758 164400 6 la_input[99]
port 324 nsew signal input
rlabel metal2 s 31390 163200 31446 164400 6 la_input[9]
port 325 nsew signal input
rlabel metal2 s 2042 163200 2098 164400 6 la_oenb[0]
port 326 nsew signal output
rlabel metal2 s 337934 163200 337990 164400 6 la_oenb[100]
port 327 nsew signal output
rlabel metal2 s 341338 163200 341394 164400 6 la_oenb[101]
port 328 nsew signal output
rlabel metal2 s 344650 163200 344706 164400 6 la_oenb[102]
port 329 nsew signal output
rlabel metal2 s 348054 163200 348110 164400 6 la_oenb[103]
port 330 nsew signal output
rlabel metal2 s 351366 163200 351422 164400 6 la_oenb[104]
port 331 nsew signal output
rlabel metal2 s 354770 163200 354826 164400 6 la_oenb[105]
port 332 nsew signal output
rlabel metal2 s 358082 163200 358138 164400 6 la_oenb[106]
port 333 nsew signal output
rlabel metal2 s 361486 163200 361542 164400 6 la_oenb[107]
port 334 nsew signal output
rlabel metal2 s 364798 163200 364854 164400 6 la_oenb[108]
port 335 nsew signal output
rlabel metal2 s 368202 163200 368258 164400 6 la_oenb[109]
port 336 nsew signal output
rlabel metal2 s 35622 163200 35678 164400 6 la_oenb[10]
port 337 nsew signal output
rlabel metal2 s 371514 163200 371570 164400 6 la_oenb[110]
port 338 nsew signal output
rlabel metal2 s 374918 163200 374974 164400 6 la_oenb[111]
port 339 nsew signal output
rlabel metal2 s 378230 163200 378286 164400 6 la_oenb[112]
port 340 nsew signal output
rlabel metal2 s 381634 163200 381690 164400 6 la_oenb[113]
port 341 nsew signal output
rlabel metal2 s 384946 163200 385002 164400 6 la_oenb[114]
port 342 nsew signal output
rlabel metal2 s 388350 163200 388406 164400 6 la_oenb[115]
port 343 nsew signal output
rlabel metal2 s 391662 163200 391718 164400 6 la_oenb[116]
port 344 nsew signal output
rlabel metal2 s 395066 163200 395122 164400 6 la_oenb[117]
port 345 nsew signal output
rlabel metal2 s 398378 163200 398434 164400 6 la_oenb[118]
port 346 nsew signal output
rlabel metal2 s 401782 163200 401838 164400 6 la_oenb[119]
port 347 nsew signal output
rlabel metal2 s 38934 163200 38990 164400 6 la_oenb[11]
port 348 nsew signal output
rlabel metal2 s 405094 163200 405150 164400 6 la_oenb[120]
port 349 nsew signal output
rlabel metal2 s 408498 163200 408554 164400 6 la_oenb[121]
port 350 nsew signal output
rlabel metal2 s 411810 163200 411866 164400 6 la_oenb[122]
port 351 nsew signal output
rlabel metal2 s 415214 163200 415270 164400 6 la_oenb[123]
port 352 nsew signal output
rlabel metal2 s 418526 163200 418582 164400 6 la_oenb[124]
port 353 nsew signal output
rlabel metal2 s 421930 163200 421986 164400 6 la_oenb[125]
port 354 nsew signal output
rlabel metal2 s 425242 163200 425298 164400 6 la_oenb[126]
port 355 nsew signal output
rlabel metal2 s 428646 163200 428702 164400 6 la_oenb[127]
port 356 nsew signal output
rlabel metal2 s 42338 163200 42394 164400 6 la_oenb[12]
port 357 nsew signal output
rlabel metal2 s 45650 163200 45706 164400 6 la_oenb[13]
port 358 nsew signal output
rlabel metal2 s 49054 163200 49110 164400 6 la_oenb[14]
port 359 nsew signal output
rlabel metal2 s 52366 163200 52422 164400 6 la_oenb[15]
port 360 nsew signal output
rlabel metal2 s 55770 163200 55826 164400 6 la_oenb[16]
port 361 nsew signal output
rlabel metal2 s 59082 163200 59138 164400 6 la_oenb[17]
port 362 nsew signal output
rlabel metal2 s 62486 163200 62542 164400 6 la_oenb[18]
port 363 nsew signal output
rlabel metal2 s 65890 163200 65946 164400 6 la_oenb[19]
port 364 nsew signal output
rlabel metal2 s 5354 163200 5410 164400 6 la_oenb[1]
port 365 nsew signal output
rlabel metal2 s 69202 163200 69258 164400 6 la_oenb[20]
port 366 nsew signal output
rlabel metal2 s 72606 163200 72662 164400 6 la_oenb[21]
port 367 nsew signal output
rlabel metal2 s 75918 163200 75974 164400 6 la_oenb[22]
port 368 nsew signal output
rlabel metal2 s 79322 163200 79378 164400 6 la_oenb[23]
port 369 nsew signal output
rlabel metal2 s 82634 163200 82690 164400 6 la_oenb[24]
port 370 nsew signal output
rlabel metal2 s 86038 163200 86094 164400 6 la_oenb[25]
port 371 nsew signal output
rlabel metal2 s 89350 163200 89406 164400 6 la_oenb[26]
port 372 nsew signal output
rlabel metal2 s 92754 163200 92810 164400 6 la_oenb[27]
port 373 nsew signal output
rlabel metal2 s 96066 163200 96122 164400 6 la_oenb[28]
port 374 nsew signal output
rlabel metal2 s 99470 163200 99526 164400 6 la_oenb[29]
port 375 nsew signal output
rlabel metal2 s 8758 163200 8814 164400 6 la_oenb[2]
port 376 nsew signal output
rlabel metal2 s 102782 163200 102838 164400 6 la_oenb[30]
port 377 nsew signal output
rlabel metal2 s 106186 163200 106242 164400 6 la_oenb[31]
port 378 nsew signal output
rlabel metal2 s 109498 163200 109554 164400 6 la_oenb[32]
port 379 nsew signal output
rlabel metal2 s 112902 163200 112958 164400 6 la_oenb[33]
port 380 nsew signal output
rlabel metal2 s 116214 163200 116270 164400 6 la_oenb[34]
port 381 nsew signal output
rlabel metal2 s 119618 163200 119674 164400 6 la_oenb[35]
port 382 nsew signal output
rlabel metal2 s 122930 163200 122986 164400 6 la_oenb[36]
port 383 nsew signal output
rlabel metal2 s 126334 163200 126390 164400 6 la_oenb[37]
port 384 nsew signal output
rlabel metal2 s 129646 163200 129702 164400 6 la_oenb[38]
port 385 nsew signal output
rlabel metal2 s 133050 163200 133106 164400 6 la_oenb[39]
port 386 nsew signal output
rlabel metal2 s 12070 163200 12126 164400 6 la_oenb[3]
port 387 nsew signal output
rlabel metal2 s 136362 163200 136418 164400 6 la_oenb[40]
port 388 nsew signal output
rlabel metal2 s 139766 163200 139822 164400 6 la_oenb[41]
port 389 nsew signal output
rlabel metal2 s 143078 163200 143134 164400 6 la_oenb[42]
port 390 nsew signal output
rlabel metal2 s 146482 163200 146538 164400 6 la_oenb[43]
port 391 nsew signal output
rlabel metal2 s 149794 163200 149850 164400 6 la_oenb[44]
port 392 nsew signal output
rlabel metal2 s 153198 163200 153254 164400 6 la_oenb[45]
port 393 nsew signal output
rlabel metal2 s 156510 163200 156566 164400 6 la_oenb[46]
port 394 nsew signal output
rlabel metal2 s 159914 163200 159970 164400 6 la_oenb[47]
port 395 nsew signal output
rlabel metal2 s 163226 163200 163282 164400 6 la_oenb[48]
port 396 nsew signal output
rlabel metal2 s 166630 163200 166686 164400 6 la_oenb[49]
port 397 nsew signal output
rlabel metal2 s 15474 163200 15530 164400 6 la_oenb[4]
port 398 nsew signal output
rlabel metal2 s 169942 163200 169998 164400 6 la_oenb[50]
port 399 nsew signal output
rlabel metal2 s 173346 163200 173402 164400 6 la_oenb[51]
port 400 nsew signal output
rlabel metal2 s 176658 163200 176714 164400 6 la_oenb[52]
port 401 nsew signal output
rlabel metal2 s 180062 163200 180118 164400 6 la_oenb[53]
port 402 nsew signal output
rlabel metal2 s 183374 163200 183430 164400 6 la_oenb[54]
port 403 nsew signal output
rlabel metal2 s 186778 163200 186834 164400 6 la_oenb[55]
port 404 nsew signal output
rlabel metal2 s 190090 163200 190146 164400 6 la_oenb[56]
port 405 nsew signal output
rlabel metal2 s 193494 163200 193550 164400 6 la_oenb[57]
port 406 nsew signal output
rlabel metal2 s 196898 163200 196954 164400 6 la_oenb[58]
port 407 nsew signal output
rlabel metal2 s 200210 163200 200266 164400 6 la_oenb[59]
port 408 nsew signal output
rlabel metal2 s 18786 163200 18842 164400 6 la_oenb[5]
port 409 nsew signal output
rlabel metal2 s 203614 163200 203670 164400 6 la_oenb[60]
port 410 nsew signal output
rlabel metal2 s 206926 163200 206982 164400 6 la_oenb[61]
port 411 nsew signal output
rlabel metal2 s 210330 163200 210386 164400 6 la_oenb[62]
port 412 nsew signal output
rlabel metal2 s 213642 163200 213698 164400 6 la_oenb[63]
port 413 nsew signal output
rlabel metal2 s 217046 163200 217102 164400 6 la_oenb[64]
port 414 nsew signal output
rlabel metal2 s 220358 163200 220414 164400 6 la_oenb[65]
port 415 nsew signal output
rlabel metal2 s 223762 163200 223818 164400 6 la_oenb[66]
port 416 nsew signal output
rlabel metal2 s 227074 163200 227130 164400 6 la_oenb[67]
port 417 nsew signal output
rlabel metal2 s 230478 163200 230534 164400 6 la_oenb[68]
port 418 nsew signal output
rlabel metal2 s 233790 163200 233846 164400 6 la_oenb[69]
port 419 nsew signal output
rlabel metal2 s 22190 163200 22246 164400 6 la_oenb[6]
port 420 nsew signal output
rlabel metal2 s 237194 163200 237250 164400 6 la_oenb[70]
port 421 nsew signal output
rlabel metal2 s 240506 163200 240562 164400 6 la_oenb[71]
port 422 nsew signal output
rlabel metal2 s 243910 163200 243966 164400 6 la_oenb[72]
port 423 nsew signal output
rlabel metal2 s 247222 163200 247278 164400 6 la_oenb[73]
port 424 nsew signal output
rlabel metal2 s 250626 163200 250682 164400 6 la_oenb[74]
port 425 nsew signal output
rlabel metal2 s 253938 163200 253994 164400 6 la_oenb[75]
port 426 nsew signal output
rlabel metal2 s 257342 163200 257398 164400 6 la_oenb[76]
port 427 nsew signal output
rlabel metal2 s 260654 163200 260710 164400 6 la_oenb[77]
port 428 nsew signal output
rlabel metal2 s 264058 163200 264114 164400 6 la_oenb[78]
port 429 nsew signal output
rlabel metal2 s 267370 163200 267426 164400 6 la_oenb[79]
port 430 nsew signal output
rlabel metal2 s 25502 163200 25558 164400 6 la_oenb[7]
port 431 nsew signal output
rlabel metal2 s 270774 163200 270830 164400 6 la_oenb[80]
port 432 nsew signal output
rlabel metal2 s 274086 163200 274142 164400 6 la_oenb[81]
port 433 nsew signal output
rlabel metal2 s 277490 163200 277546 164400 6 la_oenb[82]
port 434 nsew signal output
rlabel metal2 s 280802 163200 280858 164400 6 la_oenb[83]
port 435 nsew signal output
rlabel metal2 s 284206 163200 284262 164400 6 la_oenb[84]
port 436 nsew signal output
rlabel metal2 s 287518 163200 287574 164400 6 la_oenb[85]
port 437 nsew signal output
rlabel metal2 s 290922 163200 290978 164400 6 la_oenb[86]
port 438 nsew signal output
rlabel metal2 s 294234 163200 294290 164400 6 la_oenb[87]
port 439 nsew signal output
rlabel metal2 s 297638 163200 297694 164400 6 la_oenb[88]
port 440 nsew signal output
rlabel metal2 s 300950 163200 301006 164400 6 la_oenb[89]
port 441 nsew signal output
rlabel metal2 s 28906 163200 28962 164400 6 la_oenb[8]
port 442 nsew signal output
rlabel metal2 s 304354 163200 304410 164400 6 la_oenb[90]
port 443 nsew signal output
rlabel metal2 s 307666 163200 307722 164400 6 la_oenb[91]
port 444 nsew signal output
rlabel metal2 s 311070 163200 311126 164400 6 la_oenb[92]
port 445 nsew signal output
rlabel metal2 s 314382 163200 314438 164400 6 la_oenb[93]
port 446 nsew signal output
rlabel metal2 s 317786 163200 317842 164400 6 la_oenb[94]
port 447 nsew signal output
rlabel metal2 s 321098 163200 321154 164400 6 la_oenb[95]
port 448 nsew signal output
rlabel metal2 s 324502 163200 324558 164400 6 la_oenb[96]
port 449 nsew signal output
rlabel metal2 s 327906 163200 327962 164400 6 la_oenb[97]
port 450 nsew signal output
rlabel metal2 s 331218 163200 331274 164400 6 la_oenb[98]
port 451 nsew signal output
rlabel metal2 s 334622 163200 334678 164400 6 la_oenb[99]
port 452 nsew signal output
rlabel metal2 s 32218 163200 32274 164400 6 la_oenb[9]
port 453 nsew signal output
rlabel metal2 s 2870 163200 2926 164400 6 la_output[0]
port 454 nsew signal output
rlabel metal2 s 338762 163200 338818 164400 6 la_output[100]
port 455 nsew signal output
rlabel metal2 s 342166 163200 342222 164400 6 la_output[101]
port 456 nsew signal output
rlabel metal2 s 345478 163200 345534 164400 6 la_output[102]
port 457 nsew signal output
rlabel metal2 s 348882 163200 348938 164400 6 la_output[103]
port 458 nsew signal output
rlabel metal2 s 352194 163200 352250 164400 6 la_output[104]
port 459 nsew signal output
rlabel metal2 s 355598 163200 355654 164400 6 la_output[105]
port 460 nsew signal output
rlabel metal2 s 358910 163200 358966 164400 6 la_output[106]
port 461 nsew signal output
rlabel metal2 s 362314 163200 362370 164400 6 la_output[107]
port 462 nsew signal output
rlabel metal2 s 365626 163200 365682 164400 6 la_output[108]
port 463 nsew signal output
rlabel metal2 s 369030 163200 369086 164400 6 la_output[109]
port 464 nsew signal output
rlabel metal2 s 36450 163200 36506 164400 6 la_output[10]
port 465 nsew signal output
rlabel metal2 s 372342 163200 372398 164400 6 la_output[110]
port 466 nsew signal output
rlabel metal2 s 375746 163200 375802 164400 6 la_output[111]
port 467 nsew signal output
rlabel metal2 s 379058 163200 379114 164400 6 la_output[112]
port 468 nsew signal output
rlabel metal2 s 382462 163200 382518 164400 6 la_output[113]
port 469 nsew signal output
rlabel metal2 s 385774 163200 385830 164400 6 la_output[114]
port 470 nsew signal output
rlabel metal2 s 389178 163200 389234 164400 6 la_output[115]
port 471 nsew signal output
rlabel metal2 s 392490 163200 392546 164400 6 la_output[116]
port 472 nsew signal output
rlabel metal2 s 395894 163200 395950 164400 6 la_output[117]
port 473 nsew signal output
rlabel metal2 s 399206 163200 399262 164400 6 la_output[118]
port 474 nsew signal output
rlabel metal2 s 402610 163200 402666 164400 6 la_output[119]
port 475 nsew signal output
rlabel metal2 s 39854 163200 39910 164400 6 la_output[11]
port 476 nsew signal output
rlabel metal2 s 405922 163200 405978 164400 6 la_output[120]
port 477 nsew signal output
rlabel metal2 s 409326 163200 409382 164400 6 la_output[121]
port 478 nsew signal output
rlabel metal2 s 412638 163200 412694 164400 6 la_output[122]
port 479 nsew signal output
rlabel metal2 s 416042 163200 416098 164400 6 la_output[123]
port 480 nsew signal output
rlabel metal2 s 419354 163200 419410 164400 6 la_output[124]
port 481 nsew signal output
rlabel metal2 s 422758 163200 422814 164400 6 la_output[125]
port 482 nsew signal output
rlabel metal2 s 426162 163200 426218 164400 6 la_output[126]
port 483 nsew signal output
rlabel metal2 s 429474 163200 429530 164400 6 la_output[127]
port 484 nsew signal output
rlabel metal2 s 43166 163200 43222 164400 6 la_output[12]
port 485 nsew signal output
rlabel metal2 s 46570 163200 46626 164400 6 la_output[13]
port 486 nsew signal output
rlabel metal2 s 49882 163200 49938 164400 6 la_output[14]
port 487 nsew signal output
rlabel metal2 s 53286 163200 53342 164400 6 la_output[15]
port 488 nsew signal output
rlabel metal2 s 56598 163200 56654 164400 6 la_output[16]
port 489 nsew signal output
rlabel metal2 s 60002 163200 60058 164400 6 la_output[17]
port 490 nsew signal output
rlabel metal2 s 63314 163200 63370 164400 6 la_output[18]
port 491 nsew signal output
rlabel metal2 s 66718 163200 66774 164400 6 la_output[19]
port 492 nsew signal output
rlabel metal2 s 6182 163200 6238 164400 6 la_output[1]
port 493 nsew signal output
rlabel metal2 s 70030 163200 70086 164400 6 la_output[20]
port 494 nsew signal output
rlabel metal2 s 73434 163200 73490 164400 6 la_output[21]
port 495 nsew signal output
rlabel metal2 s 76746 163200 76802 164400 6 la_output[22]
port 496 nsew signal output
rlabel metal2 s 80150 163200 80206 164400 6 la_output[23]
port 497 nsew signal output
rlabel metal2 s 83462 163200 83518 164400 6 la_output[24]
port 498 nsew signal output
rlabel metal2 s 86866 163200 86922 164400 6 la_output[25]
port 499 nsew signal output
rlabel metal2 s 90178 163200 90234 164400 6 la_output[26]
port 500 nsew signal output
rlabel metal2 s 93582 163200 93638 164400 6 la_output[27]
port 501 nsew signal output
rlabel metal2 s 96894 163200 96950 164400 6 la_output[28]
port 502 nsew signal output
rlabel metal2 s 100298 163200 100354 164400 6 la_output[29]
port 503 nsew signal output
rlabel metal2 s 9586 163200 9642 164400 6 la_output[2]
port 504 nsew signal output
rlabel metal2 s 103610 163200 103666 164400 6 la_output[30]
port 505 nsew signal output
rlabel metal2 s 107014 163200 107070 164400 6 la_output[31]
port 506 nsew signal output
rlabel metal2 s 110326 163200 110382 164400 6 la_output[32]
port 507 nsew signal output
rlabel metal2 s 113730 163200 113786 164400 6 la_output[33]
port 508 nsew signal output
rlabel metal2 s 117042 163200 117098 164400 6 la_output[34]
port 509 nsew signal output
rlabel metal2 s 120446 163200 120502 164400 6 la_output[35]
port 510 nsew signal output
rlabel metal2 s 123758 163200 123814 164400 6 la_output[36]
port 511 nsew signal output
rlabel metal2 s 127162 163200 127218 164400 6 la_output[37]
port 512 nsew signal output
rlabel metal2 s 130474 163200 130530 164400 6 la_output[38]
port 513 nsew signal output
rlabel metal2 s 133878 163200 133934 164400 6 la_output[39]
port 514 nsew signal output
rlabel metal2 s 12898 163200 12954 164400 6 la_output[3]
port 515 nsew signal output
rlabel metal2 s 137190 163200 137246 164400 6 la_output[40]
port 516 nsew signal output
rlabel metal2 s 140594 163200 140650 164400 6 la_output[41]
port 517 nsew signal output
rlabel metal2 s 143906 163200 143962 164400 6 la_output[42]
port 518 nsew signal output
rlabel metal2 s 147310 163200 147366 164400 6 la_output[43]
port 519 nsew signal output
rlabel metal2 s 150622 163200 150678 164400 6 la_output[44]
port 520 nsew signal output
rlabel metal2 s 154026 163200 154082 164400 6 la_output[45]
port 521 nsew signal output
rlabel metal2 s 157338 163200 157394 164400 6 la_output[46]
port 522 nsew signal output
rlabel metal2 s 160742 163200 160798 164400 6 la_output[47]
port 523 nsew signal output
rlabel metal2 s 164146 163200 164202 164400 6 la_output[48]
port 524 nsew signal output
rlabel metal2 s 167458 163200 167514 164400 6 la_output[49]
port 525 nsew signal output
rlabel metal2 s 16302 163200 16358 164400 6 la_output[4]
port 526 nsew signal output
rlabel metal2 s 170862 163200 170918 164400 6 la_output[50]
port 527 nsew signal output
rlabel metal2 s 174174 163200 174230 164400 6 la_output[51]
port 528 nsew signal output
rlabel metal2 s 177578 163200 177634 164400 6 la_output[52]
port 529 nsew signal output
rlabel metal2 s 180890 163200 180946 164400 6 la_output[53]
port 530 nsew signal output
rlabel metal2 s 184294 163200 184350 164400 6 la_output[54]
port 531 nsew signal output
rlabel metal2 s 187606 163200 187662 164400 6 la_output[55]
port 532 nsew signal output
rlabel metal2 s 191010 163200 191066 164400 6 la_output[56]
port 533 nsew signal output
rlabel metal2 s 194322 163200 194378 164400 6 la_output[57]
port 534 nsew signal output
rlabel metal2 s 197726 163200 197782 164400 6 la_output[58]
port 535 nsew signal output
rlabel metal2 s 201038 163200 201094 164400 6 la_output[59]
port 536 nsew signal output
rlabel metal2 s 19614 163200 19670 164400 6 la_output[5]
port 537 nsew signal output
rlabel metal2 s 204442 163200 204498 164400 6 la_output[60]
port 538 nsew signal output
rlabel metal2 s 207754 163200 207810 164400 6 la_output[61]
port 539 nsew signal output
rlabel metal2 s 211158 163200 211214 164400 6 la_output[62]
port 540 nsew signal output
rlabel metal2 s 214470 163200 214526 164400 6 la_output[63]
port 541 nsew signal output
rlabel metal2 s 217874 163200 217930 164400 6 la_output[64]
port 542 nsew signal output
rlabel metal2 s 221186 163200 221242 164400 6 la_output[65]
port 543 nsew signal output
rlabel metal2 s 224590 163200 224646 164400 6 la_output[66]
port 544 nsew signal output
rlabel metal2 s 227902 163200 227958 164400 6 la_output[67]
port 545 nsew signal output
rlabel metal2 s 231306 163200 231362 164400 6 la_output[68]
port 546 nsew signal output
rlabel metal2 s 234618 163200 234674 164400 6 la_output[69]
port 547 nsew signal output
rlabel metal2 s 23018 163200 23074 164400 6 la_output[6]
port 548 nsew signal output
rlabel metal2 s 238022 163200 238078 164400 6 la_output[70]
port 549 nsew signal output
rlabel metal2 s 241334 163200 241390 164400 6 la_output[71]
port 550 nsew signal output
rlabel metal2 s 244738 163200 244794 164400 6 la_output[72]
port 551 nsew signal output
rlabel metal2 s 248050 163200 248106 164400 6 la_output[73]
port 552 nsew signal output
rlabel metal2 s 251454 163200 251510 164400 6 la_output[74]
port 553 nsew signal output
rlabel metal2 s 254766 163200 254822 164400 6 la_output[75]
port 554 nsew signal output
rlabel metal2 s 258170 163200 258226 164400 6 la_output[76]
port 555 nsew signal output
rlabel metal2 s 261482 163200 261538 164400 6 la_output[77]
port 556 nsew signal output
rlabel metal2 s 264886 163200 264942 164400 6 la_output[78]
port 557 nsew signal output
rlabel metal2 s 268198 163200 268254 164400 6 la_output[79]
port 558 nsew signal output
rlabel metal2 s 26330 163200 26386 164400 6 la_output[7]
port 559 nsew signal output
rlabel metal2 s 271602 163200 271658 164400 6 la_output[80]
port 560 nsew signal output
rlabel metal2 s 274914 163200 274970 164400 6 la_output[81]
port 561 nsew signal output
rlabel metal2 s 278318 163200 278374 164400 6 la_output[82]
port 562 nsew signal output
rlabel metal2 s 281630 163200 281686 164400 6 la_output[83]
port 563 nsew signal output
rlabel metal2 s 285034 163200 285090 164400 6 la_output[84]
port 564 nsew signal output
rlabel metal2 s 288346 163200 288402 164400 6 la_output[85]
port 565 nsew signal output
rlabel metal2 s 291750 163200 291806 164400 6 la_output[86]
port 566 nsew signal output
rlabel metal2 s 295154 163200 295210 164400 6 la_output[87]
port 567 nsew signal output
rlabel metal2 s 298466 163200 298522 164400 6 la_output[88]
port 568 nsew signal output
rlabel metal2 s 301870 163200 301926 164400 6 la_output[89]
port 569 nsew signal output
rlabel metal2 s 29734 163200 29790 164400 6 la_output[8]
port 570 nsew signal output
rlabel metal2 s 305182 163200 305238 164400 6 la_output[90]
port 571 nsew signal output
rlabel metal2 s 308586 163200 308642 164400 6 la_output[91]
port 572 nsew signal output
rlabel metal2 s 311898 163200 311954 164400 6 la_output[92]
port 573 nsew signal output
rlabel metal2 s 315302 163200 315358 164400 6 la_output[93]
port 574 nsew signal output
rlabel metal2 s 318614 163200 318670 164400 6 la_output[94]
port 575 nsew signal output
rlabel metal2 s 322018 163200 322074 164400 6 la_output[95]
port 576 nsew signal output
rlabel metal2 s 325330 163200 325386 164400 6 la_output[96]
port 577 nsew signal output
rlabel metal2 s 328734 163200 328790 164400 6 la_output[97]
port 578 nsew signal output
rlabel metal2 s 332046 163200 332102 164400 6 la_output[98]
port 579 nsew signal output
rlabel metal2 s 335450 163200 335506 164400 6 la_output[99]
port 580 nsew signal output
rlabel metal2 s 33138 163200 33194 164400 6 la_output[9]
port 581 nsew signal output
rlabel metal2 s 430302 163200 430358 164400 6 mprj_ack_i
port 582 nsew signal input
rlabel metal2 s 434534 163200 434590 164400 6 mprj_adr_o[0]
port 583 nsew signal output
rlabel metal2 s 463054 163200 463110 164400 6 mprj_adr_o[10]
port 584 nsew signal output
rlabel metal2 s 465630 163200 465686 164400 6 mprj_adr_o[11]
port 585 nsew signal output
rlabel metal2 s 468114 163200 468170 164400 6 mprj_adr_o[12]
port 586 nsew signal output
rlabel metal2 s 470598 163200 470654 164400 6 mprj_adr_o[13]
port 587 nsew signal output
rlabel metal2 s 473174 163200 473230 164400 6 mprj_adr_o[14]
port 588 nsew signal output
rlabel metal2 s 475658 163200 475714 164400 6 mprj_adr_o[15]
port 589 nsew signal output
rlabel metal2 s 478142 163200 478198 164400 6 mprj_adr_o[16]
port 590 nsew signal output
rlabel metal2 s 480718 163200 480774 164400 6 mprj_adr_o[17]
port 591 nsew signal output
rlabel metal2 s 483202 163200 483258 164400 6 mprj_adr_o[18]
port 592 nsew signal output
rlabel metal2 s 485778 163200 485834 164400 6 mprj_adr_o[19]
port 593 nsew signal output
rlabel metal2 s 437846 163200 437902 164400 6 mprj_adr_o[1]
port 594 nsew signal output
rlabel metal2 s 488262 163200 488318 164400 6 mprj_adr_o[20]
port 595 nsew signal output
rlabel metal2 s 490746 163200 490802 164400 6 mprj_adr_o[21]
port 596 nsew signal output
rlabel metal2 s 493322 163200 493378 164400 6 mprj_adr_o[22]
port 597 nsew signal output
rlabel metal2 s 495806 163200 495862 164400 6 mprj_adr_o[23]
port 598 nsew signal output
rlabel metal2 s 498382 163200 498438 164400 6 mprj_adr_o[24]
port 599 nsew signal output
rlabel metal2 s 500866 163200 500922 164400 6 mprj_adr_o[25]
port 600 nsew signal output
rlabel metal2 s 503350 163200 503406 164400 6 mprj_adr_o[26]
port 601 nsew signal output
rlabel metal2 s 505926 163200 505982 164400 6 mprj_adr_o[27]
port 602 nsew signal output
rlabel metal2 s 508410 163200 508466 164400 6 mprj_adr_o[28]
port 603 nsew signal output
rlabel metal2 s 510894 163200 510950 164400 6 mprj_adr_o[29]
port 604 nsew signal output
rlabel metal2 s 441250 163200 441306 164400 6 mprj_adr_o[2]
port 605 nsew signal output
rlabel metal2 s 513470 163200 513526 164400 6 mprj_adr_o[30]
port 606 nsew signal output
rlabel metal2 s 515954 163200 516010 164400 6 mprj_adr_o[31]
port 607 nsew signal output
rlabel metal2 s 444562 163200 444618 164400 6 mprj_adr_o[3]
port 608 nsew signal output
rlabel metal2 s 447966 163200 448022 164400 6 mprj_adr_o[4]
port 609 nsew signal output
rlabel metal2 s 450450 163200 450506 164400 6 mprj_adr_o[5]
port 610 nsew signal output
rlabel metal2 s 453026 163200 453082 164400 6 mprj_adr_o[6]
port 611 nsew signal output
rlabel metal2 s 455510 163200 455566 164400 6 mprj_adr_o[7]
port 612 nsew signal output
rlabel metal2 s 457994 163200 458050 164400 6 mprj_adr_o[8]
port 613 nsew signal output
rlabel metal2 s 460570 163200 460626 164400 6 mprj_adr_o[9]
port 614 nsew signal output
rlabel metal2 s 431130 163200 431186 164400 6 mprj_cyc_o
port 615 nsew signal output
rlabel metal2 s 435362 163200 435418 164400 6 mprj_dat_i[0]
port 616 nsew signal input
rlabel metal2 s 463882 163200 463938 164400 6 mprj_dat_i[10]
port 617 nsew signal input
rlabel metal2 s 466458 163200 466514 164400 6 mprj_dat_i[11]
port 618 nsew signal input
rlabel metal2 s 468942 163200 468998 164400 6 mprj_dat_i[12]
port 619 nsew signal input
rlabel metal2 s 471426 163200 471482 164400 6 mprj_dat_i[13]
port 620 nsew signal input
rlabel metal2 s 474002 163200 474058 164400 6 mprj_dat_i[14]
port 621 nsew signal input
rlabel metal2 s 476486 163200 476542 164400 6 mprj_dat_i[15]
port 622 nsew signal input
rlabel metal2 s 479062 163200 479118 164400 6 mprj_dat_i[16]
port 623 nsew signal input
rlabel metal2 s 481546 163200 481602 164400 6 mprj_dat_i[17]
port 624 nsew signal input
rlabel metal2 s 484030 163200 484086 164400 6 mprj_dat_i[18]
port 625 nsew signal input
rlabel metal2 s 486606 163200 486662 164400 6 mprj_dat_i[19]
port 626 nsew signal input
rlabel metal2 s 438674 163200 438730 164400 6 mprj_dat_i[1]
port 627 nsew signal input
rlabel metal2 s 489090 163200 489146 164400 6 mprj_dat_i[20]
port 628 nsew signal input
rlabel metal2 s 491666 163200 491722 164400 6 mprj_dat_i[21]
port 629 nsew signal input
rlabel metal2 s 494150 163200 494206 164400 6 mprj_dat_i[22]
port 630 nsew signal input
rlabel metal2 s 496634 163200 496690 164400 6 mprj_dat_i[23]
port 631 nsew signal input
rlabel metal2 s 499210 163200 499266 164400 6 mprj_dat_i[24]
port 632 nsew signal input
rlabel metal2 s 501694 163200 501750 164400 6 mprj_dat_i[25]
port 633 nsew signal input
rlabel metal2 s 504178 163200 504234 164400 6 mprj_dat_i[26]
port 634 nsew signal input
rlabel metal2 s 506754 163200 506810 164400 6 mprj_dat_i[27]
port 635 nsew signal input
rlabel metal2 s 509238 163200 509294 164400 6 mprj_dat_i[28]
port 636 nsew signal input
rlabel metal2 s 511814 163200 511870 164400 6 mprj_dat_i[29]
port 637 nsew signal input
rlabel metal2 s 442078 163200 442134 164400 6 mprj_dat_i[2]
port 638 nsew signal input
rlabel metal2 s 514298 163200 514354 164400 6 mprj_dat_i[30]
port 639 nsew signal input
rlabel metal2 s 516782 163200 516838 164400 6 mprj_dat_i[31]
port 640 nsew signal input
rlabel metal2 s 445390 163200 445446 164400 6 mprj_dat_i[3]
port 641 nsew signal input
rlabel metal2 s 448794 163200 448850 164400 6 mprj_dat_i[4]
port 642 nsew signal input
rlabel metal2 s 451278 163200 451334 164400 6 mprj_dat_i[5]
port 643 nsew signal input
rlabel metal2 s 453854 163200 453910 164400 6 mprj_dat_i[6]
port 644 nsew signal input
rlabel metal2 s 456338 163200 456394 164400 6 mprj_dat_i[7]
port 645 nsew signal input
rlabel metal2 s 458914 163200 458970 164400 6 mprj_dat_i[8]
port 646 nsew signal input
rlabel metal2 s 461398 163200 461454 164400 6 mprj_dat_i[9]
port 647 nsew signal input
rlabel metal2 s 436190 163200 436246 164400 6 mprj_dat_o[0]
port 648 nsew signal output
rlabel metal2 s 464710 163200 464766 164400 6 mprj_dat_o[10]
port 649 nsew signal output
rlabel metal2 s 467286 163200 467342 164400 6 mprj_dat_o[11]
port 650 nsew signal output
rlabel metal2 s 469770 163200 469826 164400 6 mprj_dat_o[12]
port 651 nsew signal output
rlabel metal2 s 472346 163200 472402 164400 6 mprj_dat_o[13]
port 652 nsew signal output
rlabel metal2 s 474830 163200 474886 164400 6 mprj_dat_o[14]
port 653 nsew signal output
rlabel metal2 s 477314 163200 477370 164400 6 mprj_dat_o[15]
port 654 nsew signal output
rlabel metal2 s 479890 163200 479946 164400 6 mprj_dat_o[16]
port 655 nsew signal output
rlabel metal2 s 482374 163200 482430 164400 6 mprj_dat_o[17]
port 656 nsew signal output
rlabel metal2 s 484858 163200 484914 164400 6 mprj_dat_o[18]
port 657 nsew signal output
rlabel metal2 s 487434 163200 487490 164400 6 mprj_dat_o[19]
port 658 nsew signal output
rlabel metal2 s 439594 163200 439650 164400 6 mprj_dat_o[1]
port 659 nsew signal output
rlabel metal2 s 489918 163200 489974 164400 6 mprj_dat_o[20]
port 660 nsew signal output
rlabel metal2 s 492494 163200 492550 164400 6 mprj_dat_o[21]
port 661 nsew signal output
rlabel metal2 s 494978 163200 495034 164400 6 mprj_dat_o[22]
port 662 nsew signal output
rlabel metal2 s 497462 163200 497518 164400 6 mprj_dat_o[23]
port 663 nsew signal output
rlabel metal2 s 500038 163200 500094 164400 6 mprj_dat_o[24]
port 664 nsew signal output
rlabel metal2 s 502522 163200 502578 164400 6 mprj_dat_o[25]
port 665 nsew signal output
rlabel metal2 s 505098 163200 505154 164400 6 mprj_dat_o[26]
port 666 nsew signal output
rlabel metal2 s 507582 163200 507638 164400 6 mprj_dat_o[27]
port 667 nsew signal output
rlabel metal2 s 510066 163200 510122 164400 6 mprj_dat_o[28]
port 668 nsew signal output
rlabel metal2 s 512642 163200 512698 164400 6 mprj_dat_o[29]
port 669 nsew signal output
rlabel metal2 s 442906 163200 442962 164400 6 mprj_dat_o[2]
port 670 nsew signal output
rlabel metal2 s 515126 163200 515182 164400 6 mprj_dat_o[30]
port 671 nsew signal output
rlabel metal2 s 517610 163200 517666 164400 6 mprj_dat_o[31]
port 672 nsew signal output
rlabel metal2 s 446310 163200 446366 164400 6 mprj_dat_o[3]
port 673 nsew signal output
rlabel metal2 s 449622 163200 449678 164400 6 mprj_dat_o[4]
port 674 nsew signal output
rlabel metal2 s 452106 163200 452162 164400 6 mprj_dat_o[5]
port 675 nsew signal output
rlabel metal2 s 454682 163200 454738 164400 6 mprj_dat_o[6]
port 676 nsew signal output
rlabel metal2 s 457166 163200 457222 164400 6 mprj_dat_o[7]
port 677 nsew signal output
rlabel metal2 s 459742 163200 459798 164400 6 mprj_dat_o[8]
port 678 nsew signal output
rlabel metal2 s 462226 163200 462282 164400 6 mprj_dat_o[9]
port 679 nsew signal output
rlabel metal2 s 437018 163200 437074 164400 6 mprj_sel_o[0]
port 680 nsew signal output
rlabel metal2 s 440422 163200 440478 164400 6 mprj_sel_o[1]
port 681 nsew signal output
rlabel metal2 s 443734 163200 443790 164400 6 mprj_sel_o[2]
port 682 nsew signal output
rlabel metal2 s 447138 163200 447194 164400 6 mprj_sel_o[3]
port 683 nsew signal output
rlabel metal2 s 431958 163200 432014 164400 6 mprj_stb_o
port 684 nsew signal output
rlabel metal2 s 432878 163200 432934 164400 6 mprj_wb_iena
port 685 nsew signal output
rlabel metal2 s 433706 163200 433762 164400 6 mprj_we_o
port 686 nsew signal output
rlabel metal3 s 523200 90176 524400 90296 6 qspi_enabled
port 687 nsew signal output
rlabel metal3 s 523200 84192 524400 84312 6 ser_rx
port 688 nsew signal input
rlabel metal3 s 523200 85688 524400 85808 6 ser_tx
port 689 nsew signal output
rlabel metal3 s 523200 81064 524400 81184 6 spi_csb
port 690 nsew signal output
rlabel metal3 s 523200 87184 524400 87304 6 spi_enabled
port 691 nsew signal output
rlabel metal3 s 523200 79568 524400 79688 6 spi_sck
port 692 nsew signal output
rlabel metal3 s 523200 82696 524400 82816 6 spi_sdi
port 693 nsew signal input
rlabel metal3 s 523200 78072 524400 78192 6 spi_sdo
port 694 nsew signal output
rlabel metal3 s 523200 76576 524400 76696 6 spi_sdoenb
port 695 nsew signal output
rlabel metal3 s 523200 2184 524400 2304 6 sram_ro_addr[0]
port 696 nsew signal input
rlabel metal3 s 523200 3680 524400 3800 6 sram_ro_addr[1]
port 697 nsew signal input
rlabel metal3 s 523200 5176 524400 5296 6 sram_ro_addr[2]
port 698 nsew signal input
rlabel metal3 s 523200 6672 524400 6792 6 sram_ro_addr[3]
port 699 nsew signal input
rlabel metal3 s 523200 8168 524400 8288 6 sram_ro_addr[4]
port 700 nsew signal input
rlabel metal3 s 523200 9800 524400 9920 6 sram_ro_addr[5]
port 701 nsew signal input
rlabel metal3 s 523200 11296 524400 11416 6 sram_ro_addr[6]
port 702 nsew signal input
rlabel metal3 s 523200 12792 524400 12912 6 sram_ro_addr[7]
port 703 nsew signal input
rlabel metal3 s 523200 14288 524400 14408 6 sram_ro_clk
port 704 nsew signal input
rlabel metal3 s 523200 688 524400 808 6 sram_ro_csb
port 705 nsew signal input
rlabel metal3 s 523200 15784 524400 15904 6 sram_ro_data[0]
port 706 nsew signal output
rlabel metal3 s 523200 31016 524400 31136 6 sram_ro_data[10]
port 707 nsew signal output
rlabel metal3 s 523200 32512 524400 32632 6 sram_ro_data[11]
port 708 nsew signal output
rlabel metal3 s 523200 34008 524400 34128 6 sram_ro_data[12]
port 709 nsew signal output
rlabel metal3 s 523200 35504 524400 35624 6 sram_ro_data[13]
port 710 nsew signal output
rlabel metal3 s 523200 37136 524400 37256 6 sram_ro_data[14]
port 711 nsew signal output
rlabel metal3 s 523200 38632 524400 38752 6 sram_ro_data[15]
port 712 nsew signal output
rlabel metal3 s 523200 40128 524400 40248 6 sram_ro_data[16]
port 713 nsew signal output
rlabel metal3 s 523200 41624 524400 41744 6 sram_ro_data[17]
port 714 nsew signal output
rlabel metal3 s 523200 43120 524400 43240 6 sram_ro_data[18]
port 715 nsew signal output
rlabel metal3 s 523200 44616 524400 44736 6 sram_ro_data[19]
port 716 nsew signal output
rlabel metal3 s 523200 17280 524400 17400 6 sram_ro_data[1]
port 717 nsew signal output
rlabel metal3 s 523200 46248 524400 46368 6 sram_ro_data[20]
port 718 nsew signal output
rlabel metal3 s 523200 47744 524400 47864 6 sram_ro_data[21]
port 719 nsew signal output
rlabel metal3 s 523200 49240 524400 49360 6 sram_ro_data[22]
port 720 nsew signal output
rlabel metal3 s 523200 50736 524400 50856 6 sram_ro_data[23]
port 721 nsew signal output
rlabel metal3 s 523200 52232 524400 52352 6 sram_ro_data[24]
port 722 nsew signal output
rlabel metal3 s 523200 53728 524400 53848 6 sram_ro_data[25]
port 723 nsew signal output
rlabel metal3 s 523200 55360 524400 55480 6 sram_ro_data[26]
port 724 nsew signal output
rlabel metal3 s 523200 56856 524400 56976 6 sram_ro_data[27]
port 725 nsew signal output
rlabel metal3 s 523200 58352 524400 58472 6 sram_ro_data[28]
port 726 nsew signal output
rlabel metal3 s 523200 59848 524400 59968 6 sram_ro_data[29]
port 727 nsew signal output
rlabel metal3 s 523200 18912 524400 19032 6 sram_ro_data[2]
port 728 nsew signal output
rlabel metal3 s 523200 61344 524400 61464 6 sram_ro_data[30]
port 729 nsew signal output
rlabel metal3 s 523200 62840 524400 62960 6 sram_ro_data[31]
port 730 nsew signal output
rlabel metal3 s 523200 20408 524400 20528 6 sram_ro_data[3]
port 731 nsew signal output
rlabel metal3 s 523200 21904 524400 22024 6 sram_ro_data[4]
port 732 nsew signal output
rlabel metal3 s 523200 23400 524400 23520 6 sram_ro_data[5]
port 733 nsew signal output
rlabel metal3 s 523200 24896 524400 25016 6 sram_ro_data[6]
port 734 nsew signal output
rlabel metal3 s 523200 26392 524400 26512 6 sram_ro_data[7]
port 735 nsew signal output
rlabel metal3 s 523200 28024 524400 28144 6 sram_ro_data[8]
port 736 nsew signal output
rlabel metal3 s 523200 29520 524400 29640 6 sram_ro_data[9]
port 737 nsew signal output
rlabel metal3 s 523200 70456 524400 70576 6 trap
port 738 nsew signal output
rlabel metal3 s 523200 88680 524400 88800 6 uart_enabled
port 739 nsew signal output
rlabel metal2 s 518530 163200 518586 164400 6 user_irq_ena[0]
port 740 nsew signal output
rlabel metal2 s 519358 163200 519414 164400 6 user_irq_ena[1]
port 741 nsew signal output
rlabel metal2 s 520186 163200 520242 164400 6 user_irq_ena[2]
port 742 nsew signal output
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 524000 164000
string LEFview TRUE
string GDS_FILE /project/openlane/mgmt_core_wrapper/runs/mgmt_core_wrapper/results/finishing/mgmt_core_wrapper.gds
string GDS_END 177804292
string GDS_START 176646198
<< end >>

