VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_core
  CLASS BLOCK ;
  FOREIGN mgmt_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 2000.000 BY 740.000 ;
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.020 0.780 1999.600 2.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 91.490 1999.600 93.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 221.490 1999.600 223.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 351.490 1999.600 353.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 481.490 1999.600 483.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 611.490 1999.600 613.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 737.460 1999.600 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 100.640 0.780 102.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 150.640 0.780 152.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 200.640 0.780 202.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 250.640 0.780 252.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 300.640 0.780 302.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 350.640 0.780 352.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 400.640 0.780 402.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 450.640 0.780 452.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 500.640 0.780 502.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 550.640 0.780 552.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 600.640 0.780 602.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 650.640 0.780 652.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 700.640 0.780 702.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 750.640 0.780 752.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.020 0.780 1.620 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.640 0.780 52.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 100.640 537.300 102.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 150.640 537.300 152.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 200.640 537.300 202.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 250.640 537.300 252.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 300.640 537.300 302.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 350.640 537.300 352.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 400.640 537.300 402.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 450.640 537.300 452.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 500.640 537.300 502.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 550.640 537.300 552.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 600.640 537.300 602.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 650.640 537.300 652.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 700.640 537.300 702.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 750.640 537.300 752.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 800.640 0.780 802.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 850.640 0.780 852.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 900.640 0.780 902.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 950.640 0.780 952.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1000.640 0.780 1002.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1050.640 0.780 1052.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1100.640 0.780 1102.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1150.640 0.780 1152.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1200.640 0.780 1202.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1250.640 0.780 1252.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1300.640 0.780 1302.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1350.640 0.780 1352.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1400.640 0.780 1402.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1450.640 0.780 1452.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1500.640 0.780 1502.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1550.640 0.780 1552.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1600.640 0.780 1602.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1650.640 0.780 1652.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1700.640 0.780 1702.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1750.640 0.780 1752.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1800.640 0.780 1802.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1850.640 0.780 1852.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1900.640 0.780 1902.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1950.640 0.780 1952.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1998.000 0.780 1999.600 739.060 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 3.320 4.080 1996.300 5.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 26.490 1999.600 28.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 156.490 1999.600 158.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 286.490 1999.600 288.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 416.490 1999.600 418.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 546.490 1999.600 548.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 676.490 1999.600 678.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 3.320 734.160 1996.300 735.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.640 0.780 127.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 175.640 0.780 177.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 225.640 0.780 227.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 275.640 0.780 277.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.640 0.780 327.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 375.640 0.780 377.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 425.640 0.780 427.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 475.640 0.780 477.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 525.640 0.780 527.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.640 0.780 577.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 625.640 0.780 627.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.640 0.780 677.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 725.640 0.780 727.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 775.640 0.780 777.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 3.320 4.080 4.920 735.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1994.700 4.080 1996.300 735.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 25.640 0.780 27.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 75.640 0.780 77.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.640 537.300 127.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 175.640 537.300 177.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 225.640 537.300 227.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 275.640 537.300 277.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.640 537.300 327.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 375.640 537.300 377.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 425.640 537.300 427.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 475.640 537.300 477.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 525.640 537.300 527.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.640 537.300 577.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 625.640 537.300 627.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.640 537.300 677.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 725.640 537.300 727.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 775.640 537.300 777.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 825.640 0.780 827.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 875.640 0.780 877.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 925.640 0.780 927.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 975.640 0.780 977.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.640 0.780 1027.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1075.640 0.780 1077.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1125.640 0.780 1127.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1175.640 0.780 1177.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1225.640 0.780 1227.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.640 0.780 1277.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1325.640 0.780 1327.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1375.640 0.780 1377.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1425.640 0.780 1427.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.640 0.780 1477.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1525.640 0.780 1527.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1575.640 0.780 1577.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1625.640 0.780 1627.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1675.640 0.780 1677.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1725.640 0.780 1727.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1775.640 0.780 1777.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1825.640 0.780 1827.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1875.640 0.780 1877.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1925.640 0.780 1927.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1975.640 0.780 1977.240 739.060 ;
    END
  END VPWR
  PIN core_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.790 0.000 1125.070 4.000 ;
    END
  END core_clk
  PIN core_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END core_rstn
  PIN debug_mode
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 287.680 2000.000 288.280 ;
    END
  END debug_mode
  PIN debug_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 294.480 2000.000 295.080 ;
    END
  END debug_oeb
  PIN debug_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 301.280 2000.000 301.880 ;
    END
  END debug_rx
  PIN debug_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 308.080 2000.000 308.680 ;
    END
  END debug_tx
  PIN flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 654.200 2000.000 654.800 ;
    END
  END flash_clk
  PIN flash_cs_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 647.400 2000.000 648.000 ;
    END
  END flash_cs_n
  PIN flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 661.000 2000.000 661.600 ;
    END
  END flash_io0_di
  PIN flash_io0_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 667.800 2000.000 668.400 ;
    END
  END flash_io0_do
  PIN flash_io0_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 674.600 2000.000 675.200 ;
    END
  END flash_io0_oeb
  PIN flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 681.400 2000.000 682.000 ;
    END
  END flash_io1_di
  PIN flash_io1_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 688.200 2000.000 688.800 ;
    END
  END flash_io1_do
  PIN flash_io1_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 695.000 2000.000 695.600 ;
    END
  END flash_io1_oeb
  PIN flash_io2_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 701.800 2000.000 702.400 ;
    END
  END flash_io2_di
  PIN flash_io2_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 708.600 2000.000 709.200 ;
    END
  END flash_io2_do
  PIN flash_io2_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 715.400 2000.000 716.000 ;
    END
  END flash_io2_oeb
  PIN flash_io3_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 722.200 2000.000 722.800 ;
    END
  END flash_io3_di
  PIN flash_io3_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 729.000 2000.000 729.600 ;
    END
  END flash_io3_do
  PIN flash_io3_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 735.800 2000.000 736.400 ;
    END
  END flash_io3_oeb
  PIN gpio_in_pad
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 0.000 125.030 4.000 ;
    END
  END gpio_in_pad
  PIN gpio_inenb_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.770 0.000 625.050 4.000 ;
    END
  END gpio_inenb_pad
  PIN gpio_mode0_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.550 0.000 874.830 4.000 ;
    END
  END gpio_mode0_pad
  PIN gpio_mode1_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1374.570 0.000 1374.850 4.000 ;
    END
  END gpio_mode1_pad
  PIN gpio_out_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1624.810 0.000 1625.090 4.000 ;
    END
  END gpio_out_pad
  PIN gpio_outenb_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1874.590 0.000 1874.870 4.000 ;
    END
  END gpio_outenb_pad
  PIN hk_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 409.400 2000.000 410.000 ;
    END
  END hk_ack_i
  PIN hk_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 423.000 2000.000 423.600 ;
    END
  END hk_cyc_o
  PIN hk_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 429.800 2000.000 430.400 ;
    END
  END hk_dat_i[0]
  PIN hk_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 497.800 2000.000 498.400 ;
    END
  END hk_dat_i[10]
  PIN hk_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 504.600 2000.000 505.200 ;
    END
  END hk_dat_i[11]
  PIN hk_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 511.400 2000.000 512.000 ;
    END
  END hk_dat_i[12]
  PIN hk_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 518.200 2000.000 518.800 ;
    END
  END hk_dat_i[13]
  PIN hk_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 525.000 2000.000 525.600 ;
    END
  END hk_dat_i[14]
  PIN hk_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 531.800 2000.000 532.400 ;
    END
  END hk_dat_i[15]
  PIN hk_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 538.600 2000.000 539.200 ;
    END
  END hk_dat_i[16]
  PIN hk_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 545.400 2000.000 546.000 ;
    END
  END hk_dat_i[17]
  PIN hk_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 552.200 2000.000 552.800 ;
    END
  END hk_dat_i[18]
  PIN hk_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 559.000 2000.000 559.600 ;
    END
  END hk_dat_i[19]
  PIN hk_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 436.600 2000.000 437.200 ;
    END
  END hk_dat_i[1]
  PIN hk_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 565.800 2000.000 566.400 ;
    END
  END hk_dat_i[20]
  PIN hk_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 572.600 2000.000 573.200 ;
    END
  END hk_dat_i[21]
  PIN hk_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 579.400 2000.000 580.000 ;
    END
  END hk_dat_i[22]
  PIN hk_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 586.200 2000.000 586.800 ;
    END
  END hk_dat_i[23]
  PIN hk_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 593.000 2000.000 593.600 ;
    END
  END hk_dat_i[24]
  PIN hk_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 599.800 2000.000 600.400 ;
    END
  END hk_dat_i[25]
  PIN hk_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 606.600 2000.000 607.200 ;
    END
  END hk_dat_i[26]
  PIN hk_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 613.400 2000.000 614.000 ;
    END
  END hk_dat_i[27]
  PIN hk_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 620.200 2000.000 620.800 ;
    END
  END hk_dat_i[28]
  PIN hk_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 627.000 2000.000 627.600 ;
    END
  END hk_dat_i[29]
  PIN hk_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 443.400 2000.000 444.000 ;
    END
  END hk_dat_i[2]
  PIN hk_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 633.800 2000.000 634.400 ;
    END
  END hk_dat_i[30]
  PIN hk_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 640.600 2000.000 641.200 ;
    END
  END hk_dat_i[31]
  PIN hk_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 450.200 2000.000 450.800 ;
    END
  END hk_dat_i[3]
  PIN hk_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 457.000 2000.000 457.600 ;
    END
  END hk_dat_i[4]
  PIN hk_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 463.800 2000.000 464.400 ;
    END
  END hk_dat_i[5]
  PIN hk_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 470.600 2000.000 471.200 ;
    END
  END hk_dat_i[6]
  PIN hk_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 477.400 2000.000 478.000 ;
    END
  END hk_dat_i[7]
  PIN hk_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 484.200 2000.000 484.800 ;
    END
  END hk_dat_i[8]
  PIN hk_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 491.000 2000.000 491.600 ;
    END
  END hk_dat_i[9]
  PIN hk_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 416.200 2000.000 416.800 ;
    END
  END hk_stb_o
  PIN la_iena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 736.000 1.750 740.000 ;
    END
  END la_iena[0]
  PIN la_iena[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.330 736.000 1285.610 740.000 ;
    END
  END la_iena[100]
  PIN la_iena[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.210 736.000 1298.490 740.000 ;
    END
  END la_iena[101]
  PIN la_iena[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1311.090 736.000 1311.370 740.000 ;
    END
  END la_iena[102]
  PIN la_iena[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.970 736.000 1324.250 740.000 ;
    END
  END la_iena[103]
  PIN la_iena[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1336.850 736.000 1337.130 740.000 ;
    END
  END la_iena[104]
  PIN la_iena[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.730 736.000 1350.010 740.000 ;
    END
  END la_iena[105]
  PIN la_iena[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.610 736.000 1362.890 740.000 ;
    END
  END la_iena[106]
  PIN la_iena[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.490 736.000 1375.770 740.000 ;
    END
  END la_iena[107]
  PIN la_iena[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.910 736.000 1388.190 740.000 ;
    END
  END la_iena[108]
  PIN la_iena[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.790 736.000 1401.070 740.000 ;
    END
  END la_iena[109]
  PIN la_iena[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 736.000 130.090 740.000 ;
    END
  END la_iena[10]
  PIN la_iena[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.670 736.000 1413.950 740.000 ;
    END
  END la_iena[110]
  PIN la_iena[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.550 736.000 1426.830 740.000 ;
    END
  END la_iena[111]
  PIN la_iena[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.430 736.000 1439.710 740.000 ;
    END
  END la_iena[112]
  PIN la_iena[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1452.310 736.000 1452.590 740.000 ;
    END
  END la_iena[113]
  PIN la_iena[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1465.190 736.000 1465.470 740.000 ;
    END
  END la_iena[114]
  PIN la_iena[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.070 736.000 1478.350 740.000 ;
    END
  END la_iena[115]
  PIN la_iena[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 736.000 1491.230 740.000 ;
    END
  END la_iena[116]
  PIN la_iena[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.830 736.000 1504.110 740.000 ;
    END
  END la_iena[117]
  PIN la_iena[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1516.710 736.000 1516.990 740.000 ;
    END
  END la_iena[118]
  PIN la_iena[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1529.590 736.000 1529.870 740.000 ;
    END
  END la_iena[119]
  PIN la_iena[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 736.000 142.970 740.000 ;
    END
  END la_iena[11]
  PIN la_iena[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.010 736.000 1542.290 740.000 ;
    END
  END la_iena[120]
  PIN la_iena[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1554.890 736.000 1555.170 740.000 ;
    END
  END la_iena[121]
  PIN la_iena[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1567.770 736.000 1568.050 740.000 ;
    END
  END la_iena[122]
  PIN la_iena[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.650 736.000 1580.930 740.000 ;
    END
  END la_iena[123]
  PIN la_iena[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1593.530 736.000 1593.810 740.000 ;
    END
  END la_iena[124]
  PIN la_iena[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1606.410 736.000 1606.690 740.000 ;
    END
  END la_iena[125]
  PIN la_iena[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1619.290 736.000 1619.570 740.000 ;
    END
  END la_iena[126]
  PIN la_iena[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.170 736.000 1632.450 740.000 ;
    END
  END la_iena[127]
  PIN la_iena[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 736.000 155.390 740.000 ;
    END
  END la_iena[12]
  PIN la_iena[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 736.000 168.270 740.000 ;
    END
  END la_iena[13]
  PIN la_iena[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 736.000 181.150 740.000 ;
    END
  END la_iena[14]
  PIN la_iena[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 736.000 194.030 740.000 ;
    END
  END la_iena[15]
  PIN la_iena[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.630 736.000 206.910 740.000 ;
    END
  END la_iena[16]
  PIN la_iena[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 736.000 219.790 740.000 ;
    END
  END la_iena[17]
  PIN la_iena[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 736.000 232.670 740.000 ;
    END
  END la_iena[18]
  PIN la_iena[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 736.000 245.550 740.000 ;
    END
  END la_iena[19]
  PIN la_iena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 736.000 14.170 740.000 ;
    END
  END la_iena[1]
  PIN la_iena[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 736.000 258.430 740.000 ;
    END
  END la_iena[20]
  PIN la_iena[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 736.000 271.310 740.000 ;
    END
  END la_iena[21]
  PIN la_iena[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.910 736.000 284.190 740.000 ;
    END
  END la_iena[22]
  PIN la_iena[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 736.000 297.070 740.000 ;
    END
  END la_iena[23]
  PIN la_iena[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 736.000 309.490 740.000 ;
    END
  END la_iena[24]
  PIN la_iena[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 736.000 322.370 740.000 ;
    END
  END la_iena[25]
  PIN la_iena[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 736.000 335.250 740.000 ;
    END
  END la_iena[26]
  PIN la_iena[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 736.000 348.130 740.000 ;
    END
  END la_iena[27]
  PIN la_iena[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 736.000 361.010 740.000 ;
    END
  END la_iena[28]
  PIN la_iena[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.610 736.000 373.890 740.000 ;
    END
  END la_iena[29]
  PIN la_iena[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 736.000 27.050 740.000 ;
    END
  END la_iena[2]
  PIN la_iena[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 736.000 386.770 740.000 ;
    END
  END la_iena[30]
  PIN la_iena[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 736.000 399.650 740.000 ;
    END
  END la_iena[31]
  PIN la_iena[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 736.000 412.530 740.000 ;
    END
  END la_iena[32]
  PIN la_iena[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 736.000 425.410 740.000 ;
    END
  END la_iena[33]
  PIN la_iena[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 736.000 438.290 740.000 ;
    END
  END la_iena[34]
  PIN la_iena[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 736.000 451.170 740.000 ;
    END
  END la_iena[35]
  PIN la_iena[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.310 736.000 463.590 740.000 ;
    END
  END la_iena[36]
  PIN la_iena[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 736.000 476.470 740.000 ;
    END
  END la_iena[37]
  PIN la_iena[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 736.000 489.350 740.000 ;
    END
  END la_iena[38]
  PIN la_iena[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 736.000 502.230 740.000 ;
    END
  END la_iena[39]
  PIN la_iena[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 736.000 39.930 740.000 ;
    END
  END la_iena[3]
  PIN la_iena[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 736.000 515.110 740.000 ;
    END
  END la_iena[40]
  PIN la_iena[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.710 736.000 527.990 740.000 ;
    END
  END la_iena[41]
  PIN la_iena[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 736.000 540.870 740.000 ;
    END
  END la_iena[42]
  PIN la_iena[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.470 736.000 553.750 740.000 ;
    END
  END la_iena[43]
  PIN la_iena[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.350 736.000 566.630 740.000 ;
    END
  END la_iena[44]
  PIN la_iena[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 736.000 579.510 740.000 ;
    END
  END la_iena[45]
  PIN la_iena[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.110 736.000 592.390 740.000 ;
    END
  END la_iena[46]
  PIN la_iena[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.990 736.000 605.270 740.000 ;
    END
  END la_iena[47]
  PIN la_iena[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 736.000 617.690 740.000 ;
    END
  END la_iena[48]
  PIN la_iena[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.290 736.000 630.570 740.000 ;
    END
  END la_iena[49]
  PIN la_iena[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 736.000 52.810 740.000 ;
    END
  END la_iena[4]
  PIN la_iena[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 736.000 643.450 740.000 ;
    END
  END la_iena[50]
  PIN la_iena[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.050 736.000 656.330 740.000 ;
    END
  END la_iena[51]
  PIN la_iena[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 736.000 669.210 740.000 ;
    END
  END la_iena[52]
  PIN la_iena[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.810 736.000 682.090 740.000 ;
    END
  END la_iena[53]
  PIN la_iena[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.690 736.000 694.970 740.000 ;
    END
  END la_iena[54]
  PIN la_iena[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 736.000 707.850 740.000 ;
    END
  END la_iena[55]
  PIN la_iena[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.450 736.000 720.730 740.000 ;
    END
  END la_iena[56]
  PIN la_iena[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.330 736.000 733.610 740.000 ;
    END
  END la_iena[57]
  PIN la_iena[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 736.000 746.490 740.000 ;
    END
  END la_iena[58]
  PIN la_iena[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 736.000 759.370 740.000 ;
    END
  END la_iena[59]
  PIN la_iena[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 736.000 65.690 740.000 ;
    END
  END la_iena[5]
  PIN la_iena[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 736.000 771.790 740.000 ;
    END
  END la_iena[60]
  PIN la_iena[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 736.000 784.670 740.000 ;
    END
  END la_iena[61]
  PIN la_iena[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.270 736.000 797.550 740.000 ;
    END
  END la_iena[62]
  PIN la_iena[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.150 736.000 810.430 740.000 ;
    END
  END la_iena[63]
  PIN la_iena[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.030 736.000 823.310 740.000 ;
    END
  END la_iena[64]
  PIN la_iena[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.910 736.000 836.190 740.000 ;
    END
  END la_iena[65]
  PIN la_iena[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 736.000 849.070 740.000 ;
    END
  END la_iena[66]
  PIN la_iena[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.670 736.000 861.950 740.000 ;
    END
  END la_iena[67]
  PIN la_iena[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.550 736.000 874.830 740.000 ;
    END
  END la_iena[68]
  PIN la_iena[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.430 736.000 887.710 740.000 ;
    END
  END la_iena[69]
  PIN la_iena[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.290 736.000 78.570 740.000 ;
    END
  END la_iena[6]
  PIN la_iena[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.310 736.000 900.590 740.000 ;
    END
  END la_iena[70]
  PIN la_iena[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 913.190 736.000 913.470 740.000 ;
    END
  END la_iena[71]
  PIN la_iena[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 925.610 736.000 925.890 740.000 ;
    END
  END la_iena[72]
  PIN la_iena[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.490 736.000 938.770 740.000 ;
    END
  END la_iena[73]
  PIN la_iena[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.370 736.000 951.650 740.000 ;
    END
  END la_iena[74]
  PIN la_iena[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 964.250 736.000 964.530 740.000 ;
    END
  END la_iena[75]
  PIN la_iena[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.130 736.000 977.410 740.000 ;
    END
  END la_iena[76]
  PIN la_iena[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.010 736.000 990.290 740.000 ;
    END
  END la_iena[77]
  PIN la_iena[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.890 736.000 1003.170 740.000 ;
    END
  END la_iena[78]
  PIN la_iena[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.770 736.000 1016.050 740.000 ;
    END
  END la_iena[79]
  PIN la_iena[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.170 736.000 91.450 740.000 ;
    END
  END la_iena[7]
  PIN la_iena[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1028.650 736.000 1028.930 740.000 ;
    END
  END la_iena[80]
  PIN la_iena[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.530 736.000 1041.810 740.000 ;
    END
  END la_iena[81]
  PIN la_iena[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.410 736.000 1054.690 740.000 ;
    END
  END la_iena[82]
  PIN la_iena[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.290 736.000 1067.570 740.000 ;
    END
  END la_iena[83]
  PIN la_iena[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1079.710 736.000 1079.990 740.000 ;
    END
  END la_iena[84]
  PIN la_iena[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.590 736.000 1092.870 740.000 ;
    END
  END la_iena[85]
  PIN la_iena[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.470 736.000 1105.750 740.000 ;
    END
  END la_iena[86]
  PIN la_iena[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1118.350 736.000 1118.630 740.000 ;
    END
  END la_iena[87]
  PIN la_iena[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.230 736.000 1131.510 740.000 ;
    END
  END la_iena[88]
  PIN la_iena[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1144.110 736.000 1144.390 740.000 ;
    END
  END la_iena[89]
  PIN la_iena[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 736.000 104.330 740.000 ;
    END
  END la_iena[8]
  PIN la_iena[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.990 736.000 1157.270 740.000 ;
    END
  END la_iena[90]
  PIN la_iena[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.870 736.000 1170.150 740.000 ;
    END
  END la_iena[91]
  PIN la_iena[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1182.750 736.000 1183.030 740.000 ;
    END
  END la_iena[92]
  PIN la_iena[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1195.630 736.000 1195.910 740.000 ;
    END
  END la_iena[93]
  PIN la_iena[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.510 736.000 1208.790 740.000 ;
    END
  END la_iena[94]
  PIN la_iena[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.390 736.000 1221.670 740.000 ;
    END
  END la_iena[95]
  PIN la_iena[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.810 736.000 1234.090 740.000 ;
    END
  END la_iena[96]
  PIN la_iena[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.690 736.000 1246.970 740.000 ;
    END
  END la_iena[97]
  PIN la_iena[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1259.570 736.000 1259.850 740.000 ;
    END
  END la_iena[98]
  PIN la_iena[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1272.450 736.000 1272.730 740.000 ;
    END
  END la_iena[99]
  PIN la_iena[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 736.000 117.210 740.000 ;
    END
  END la_iena[9]
  PIN la_input[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 736.000 4.510 740.000 ;
    END
  END la_input[0]
  PIN la_input[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1288.550 736.000 1288.830 740.000 ;
    END
  END la_input[100]
  PIN la_input[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.430 736.000 1301.710 740.000 ;
    END
  END la_input[101]
  PIN la_input[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.310 736.000 1314.590 740.000 ;
    END
  END la_input[102]
  PIN la_input[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1327.190 736.000 1327.470 740.000 ;
    END
  END la_input[103]
  PIN la_input[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.070 736.000 1340.350 740.000 ;
    END
  END la_input[104]
  PIN la_input[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.950 736.000 1353.230 740.000 ;
    END
  END la_input[105]
  PIN la_input[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1365.830 736.000 1366.110 740.000 ;
    END
  END la_input[106]
  PIN la_input[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.710 736.000 1378.990 740.000 ;
    END
  END la_input[107]
  PIN la_input[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.130 736.000 1391.410 740.000 ;
    END
  END la_input[108]
  PIN la_input[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.010 736.000 1404.290 740.000 ;
    END
  END la_input[109]
  PIN la_input[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.030 736.000 133.310 740.000 ;
    END
  END la_input[10]
  PIN la_input[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1416.890 736.000 1417.170 740.000 ;
    END
  END la_input[110]
  PIN la_input[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.770 736.000 1430.050 740.000 ;
    END
  END la_input[111]
  PIN la_input[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.650 736.000 1442.930 740.000 ;
    END
  END la_input[112]
  PIN la_input[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.530 736.000 1455.810 740.000 ;
    END
  END la_input[113]
  PIN la_input[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.410 736.000 1468.690 740.000 ;
    END
  END la_input[114]
  PIN la_input[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.290 736.000 1481.570 740.000 ;
    END
  END la_input[115]
  PIN la_input[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.170 736.000 1494.450 740.000 ;
    END
  END la_input[116]
  PIN la_input[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.050 736.000 1507.330 740.000 ;
    END
  END la_input[117]
  PIN la_input[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.930 736.000 1520.210 740.000 ;
    END
  END la_input[118]
  PIN la_input[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1532.810 736.000 1533.090 740.000 ;
    END
  END la_input[119]
  PIN la_input[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 736.000 146.190 740.000 ;
    END
  END la_input[11]
  PIN la_input[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.230 736.000 1545.510 740.000 ;
    END
  END la_input[120]
  PIN la_input[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1558.110 736.000 1558.390 740.000 ;
    END
  END la_input[121]
  PIN la_input[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1570.990 736.000 1571.270 740.000 ;
    END
  END la_input[122]
  PIN la_input[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1583.870 736.000 1584.150 740.000 ;
    END
  END la_input[123]
  PIN la_input[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1596.750 736.000 1597.030 740.000 ;
    END
  END la_input[124]
  PIN la_input[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1609.630 736.000 1609.910 740.000 ;
    END
  END la_input[125]
  PIN la_input[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.510 736.000 1622.790 740.000 ;
    END
  END la_input[126]
  PIN la_input[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.390 736.000 1635.670 740.000 ;
    END
  END la_input[127]
  PIN la_input[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 736.000 158.610 740.000 ;
    END
  END la_input[12]
  PIN la_input[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 736.000 171.490 740.000 ;
    END
  END la_input[13]
  PIN la_input[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 736.000 184.370 740.000 ;
    END
  END la_input[14]
  PIN la_input[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 736.000 197.250 740.000 ;
    END
  END la_input[15]
  PIN la_input[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 736.000 210.130 740.000 ;
    END
  END la_input[16]
  PIN la_input[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.730 736.000 223.010 740.000 ;
    END
  END la_input[17]
  PIN la_input[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 736.000 235.890 740.000 ;
    END
  END la_input[18]
  PIN la_input[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 736.000 248.770 740.000 ;
    END
  END la_input[19]
  PIN la_input[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.110 736.000 17.390 740.000 ;
    END
  END la_input[1]
  PIN la_input[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 736.000 261.650 740.000 ;
    END
  END la_input[20]
  PIN la_input[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 736.000 274.530 740.000 ;
    END
  END la_input[21]
  PIN la_input[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 736.000 287.410 740.000 ;
    END
  END la_input[22]
  PIN la_input[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 736.000 300.290 740.000 ;
    END
  END la_input[23]
  PIN la_input[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 736.000 312.710 740.000 ;
    END
  END la_input[24]
  PIN la_input[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 736.000 325.590 740.000 ;
    END
  END la_input[25]
  PIN la_input[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 736.000 338.470 740.000 ;
    END
  END la_input[26]
  PIN la_input[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.070 736.000 351.350 740.000 ;
    END
  END la_input[27]
  PIN la_input[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 736.000 364.230 740.000 ;
    END
  END la_input[28]
  PIN la_input[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 736.000 377.110 740.000 ;
    END
  END la_input[29]
  PIN la_input[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.990 736.000 30.270 740.000 ;
    END
  END la_input[2]
  PIN la_input[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 736.000 389.990 740.000 ;
    END
  END la_input[30]
  PIN la_input[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 736.000 402.870 740.000 ;
    END
  END la_input[31]
  PIN la_input[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 736.000 415.750 740.000 ;
    END
  END la_input[32]
  PIN la_input[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 736.000 428.630 740.000 ;
    END
  END la_input[33]
  PIN la_input[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 736.000 441.510 740.000 ;
    END
  END la_input[34]
  PIN la_input[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 736.000 454.390 740.000 ;
    END
  END la_input[35]
  PIN la_input[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.530 736.000 466.810 740.000 ;
    END
  END la_input[36]
  PIN la_input[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 736.000 479.690 740.000 ;
    END
  END la_input[37]
  PIN la_input[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 736.000 492.570 740.000 ;
    END
  END la_input[38]
  PIN la_input[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 736.000 505.450 740.000 ;
    END
  END la_input[39]
  PIN la_input[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 736.000 43.150 740.000 ;
    END
  END la_input[3]
  PIN la_input[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 736.000 518.330 740.000 ;
    END
  END la_input[40]
  PIN la_input[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.930 736.000 531.210 740.000 ;
    END
  END la_input[41]
  PIN la_input[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 736.000 544.090 740.000 ;
    END
  END la_input[42]
  PIN la_input[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 736.000 556.970 740.000 ;
    END
  END la_input[43]
  PIN la_input[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 736.000 569.850 740.000 ;
    END
  END la_input[44]
  PIN la_input[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.450 736.000 582.730 740.000 ;
    END
  END la_input[45]
  PIN la_input[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 736.000 595.610 740.000 ;
    END
  END la_input[46]
  PIN la_input[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.210 736.000 608.490 740.000 ;
    END
  END la_input[47]
  PIN la_input[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 736.000 620.910 740.000 ;
    END
  END la_input[48]
  PIN la_input[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.510 736.000 633.790 740.000 ;
    END
  END la_input[49]
  PIN la_input[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 736.000 56.030 740.000 ;
    END
  END la_input[4]
  PIN la_input[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 736.000 646.670 740.000 ;
    END
  END la_input[50]
  PIN la_input[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.270 736.000 659.550 740.000 ;
    END
  END la_input[51]
  PIN la_input[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.150 736.000 672.430 740.000 ;
    END
  END la_input[52]
  PIN la_input[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.030 736.000 685.310 740.000 ;
    END
  END la_input[53]
  PIN la_input[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.910 736.000 698.190 740.000 ;
    END
  END la_input[54]
  PIN la_input[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.790 736.000 711.070 740.000 ;
    END
  END la_input[55]
  PIN la_input[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.670 736.000 723.950 740.000 ;
    END
  END la_input[56]
  PIN la_input[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.550 736.000 736.830 740.000 ;
    END
  END la_input[57]
  PIN la_input[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 736.000 749.710 740.000 ;
    END
  END la_input[58]
  PIN la_input[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.310 736.000 762.590 740.000 ;
    END
  END la_input[59]
  PIN la_input[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.630 736.000 68.910 740.000 ;
    END
  END la_input[5]
  PIN la_input[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.730 736.000 775.010 740.000 ;
    END
  END la_input[60]
  PIN la_input[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.610 736.000 787.890 740.000 ;
    END
  END la_input[61]
  PIN la_input[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.490 736.000 800.770 740.000 ;
    END
  END la_input[62]
  PIN la_input[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.370 736.000 813.650 740.000 ;
    END
  END la_input[63]
  PIN la_input[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.250 736.000 826.530 740.000 ;
    END
  END la_input[64]
  PIN la_input[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.130 736.000 839.410 740.000 ;
    END
  END la_input[65]
  PIN la_input[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.010 736.000 852.290 740.000 ;
    END
  END la_input[66]
  PIN la_input[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 864.890 736.000 865.170 740.000 ;
    END
  END la_input[67]
  PIN la_input[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.770 736.000 878.050 740.000 ;
    END
  END la_input[68]
  PIN la_input[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.650 736.000 890.930 740.000 ;
    END
  END la_input[69]
  PIN la_input[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.510 736.000 81.790 740.000 ;
    END
  END la_input[6]
  PIN la_input[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.530 736.000 903.810 740.000 ;
    END
  END la_input[70]
  PIN la_input[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.410 736.000 916.690 740.000 ;
    END
  END la_input[71]
  PIN la_input[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.830 736.000 929.110 740.000 ;
    END
  END la_input[72]
  PIN la_input[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.710 736.000 941.990 740.000 ;
    END
  END la_input[73]
  PIN la_input[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.590 736.000 954.870 740.000 ;
    END
  END la_input[74]
  PIN la_input[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.470 736.000 967.750 740.000 ;
    END
  END la_input[75]
  PIN la_input[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.350 736.000 980.630 740.000 ;
    END
  END la_input[76]
  PIN la_input[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.230 736.000 993.510 740.000 ;
    END
  END la_input[77]
  PIN la_input[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1006.110 736.000 1006.390 740.000 ;
    END
  END la_input[78]
  PIN la_input[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.990 736.000 1019.270 740.000 ;
    END
  END la_input[79]
  PIN la_input[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 736.000 94.670 740.000 ;
    END
  END la_input[7]
  PIN la_input[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.870 736.000 1032.150 740.000 ;
    END
  END la_input[80]
  PIN la_input[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.750 736.000 1045.030 740.000 ;
    END
  END la_input[81]
  PIN la_input[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1057.630 736.000 1057.910 740.000 ;
    END
  END la_input[82]
  PIN la_input[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.510 736.000 1070.790 740.000 ;
    END
  END la_input[83]
  PIN la_input[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.930 736.000 1083.210 740.000 ;
    END
  END la_input[84]
  PIN la_input[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.810 736.000 1096.090 740.000 ;
    END
  END la_input[85]
  PIN la_input[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.690 736.000 1108.970 740.000 ;
    END
  END la_input[86]
  PIN la_input[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.570 736.000 1121.850 740.000 ;
    END
  END la_input[87]
  PIN la_input[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.450 736.000 1134.730 740.000 ;
    END
  END la_input[88]
  PIN la_input[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.330 736.000 1147.610 740.000 ;
    END
  END la_input[89]
  PIN la_input[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 736.000 107.550 740.000 ;
    END
  END la_input[8]
  PIN la_input[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.210 736.000 1160.490 740.000 ;
    END
  END la_input[90]
  PIN la_input[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.090 736.000 1173.370 740.000 ;
    END
  END la_input[91]
  PIN la_input[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.970 736.000 1186.250 740.000 ;
    END
  END la_input[92]
  PIN la_input[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1198.850 736.000 1199.130 740.000 ;
    END
  END la_input[93]
  PIN la_input[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1211.730 736.000 1212.010 740.000 ;
    END
  END la_input[94]
  PIN la_input[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.610 736.000 1224.890 740.000 ;
    END
  END la_input[95]
  PIN la_input[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.030 736.000 1237.310 740.000 ;
    END
  END la_input[96]
  PIN la_input[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.910 736.000 1250.190 740.000 ;
    END
  END la_input[97]
  PIN la_input[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1262.790 736.000 1263.070 740.000 ;
    END
  END la_input[98]
  PIN la_input[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.670 736.000 1275.950 740.000 ;
    END
  END la_input[99]
  PIN la_input[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 736.000 120.430 740.000 ;
    END
  END la_input[9]
  PIN la_oenb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 736.000 7.730 740.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.770 736.000 1292.050 740.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.650 736.000 1304.930 740.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.530 736.000 1317.810 740.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1330.410 736.000 1330.690 740.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1343.290 736.000 1343.570 740.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.170 736.000 1356.450 740.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1369.050 736.000 1369.330 740.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.930 736.000 1382.210 740.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1394.350 736.000 1394.630 740.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.230 736.000 1407.510 740.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 736.000 136.530 740.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.110 736.000 1420.390 740.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.990 736.000 1433.270 740.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.870 736.000 1446.150 740.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.750 736.000 1459.030 740.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.630 736.000 1471.910 740.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.510 736.000 1484.790 740.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.390 736.000 1497.670 740.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1510.270 736.000 1510.550 740.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.150 736.000 1523.430 740.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.030 736.000 1536.310 740.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.130 736.000 149.410 740.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1548.450 736.000 1548.730 740.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.330 736.000 1561.610 740.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.210 736.000 1574.490 740.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1587.090 736.000 1587.370 740.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1599.970 736.000 1600.250 740.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1612.850 736.000 1613.130 740.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1625.730 736.000 1626.010 740.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1638.610 736.000 1638.890 740.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 736.000 161.830 740.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 736.000 174.710 740.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.310 736.000 187.590 740.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 736.000 200.470 740.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.070 736.000 213.350 740.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 736.000 226.230 740.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 736.000 239.110 740.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 736.000 251.990 740.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.330 736.000 20.610 740.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 736.000 264.870 740.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 736.000 277.750 740.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 736.000 290.630 740.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.230 736.000 303.510 740.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 736.000 315.930 740.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 736.000 328.810 740.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 736.000 341.690 740.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 736.000 354.570 740.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 736.000 367.450 740.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 736.000 380.330 740.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.210 736.000 33.490 740.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 736.000 393.210 740.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 736.000 406.090 740.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.690 736.000 418.970 740.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 736.000 431.850 740.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 736.000 444.730 740.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 736.000 457.610 740.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 736.000 470.030 740.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 736.000 482.910 740.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 736.000 495.790 740.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 736.000 508.670 740.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.090 736.000 46.370 740.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 736.000 521.550 740.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.150 736.000 534.430 740.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 736.000 547.310 740.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.910 736.000 560.190 740.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 736.000 573.070 740.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 736.000 585.950 740.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.550 736.000 598.830 740.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.430 736.000 611.710 740.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 736.000 624.130 740.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.730 736.000 637.010 740.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 736.000 59.250 740.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 736.000 649.890 740.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 736.000 662.770 740.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.370 736.000 675.650 740.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.250 736.000 688.530 740.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.130 736.000 701.410 740.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.010 736.000 714.290 740.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.890 736.000 727.170 740.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.770 736.000 740.050 740.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 736.000 752.930 740.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.530 736.000 765.810 740.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 736.000 72.130 740.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.950 736.000 778.230 740.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 790.830 736.000 791.110 740.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 803.710 736.000 803.990 740.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.590 736.000 816.870 740.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.470 736.000 829.750 740.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.350 736.000 842.630 740.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.230 736.000 855.510 740.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.110 736.000 868.390 740.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.990 736.000 881.270 740.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.870 736.000 894.150 740.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 736.000 85.010 740.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 906.750 736.000 907.030 740.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.630 736.000 919.910 740.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.050 736.000 932.330 740.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.930 736.000 945.210 740.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.810 736.000 958.090 740.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.690 736.000 970.970 740.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.570 736.000 983.850 740.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.450 736.000 996.730 740.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.330 736.000 1009.610 740.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.210 736.000 1022.490 740.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 736.000 97.890 740.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.090 736.000 1035.370 740.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.970 736.000 1048.250 740.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.850 736.000 1061.130 740.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.730 736.000 1074.010 740.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.150 736.000 1086.430 740.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.030 736.000 1099.310 740.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.910 736.000 1112.190 740.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.790 736.000 1125.070 740.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.670 736.000 1137.950 740.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.550 736.000 1150.830 740.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.490 736.000 110.770 740.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1163.430 736.000 1163.710 740.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.310 736.000 1176.590 740.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1189.190 736.000 1189.470 740.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.070 736.000 1202.350 740.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.950 736.000 1215.230 740.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.830 736.000 1228.110 740.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1240.250 736.000 1240.530 740.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.130 736.000 1253.410 740.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.010 736.000 1266.290 740.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1278.890 736.000 1279.170 740.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 736.000 123.650 740.000 ;
    END
  END la_oenb[9]
  PIN la_output[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 10.670 736.000 10.950 740.000 ;
    END
  END la_output[0]
  PIN la_output[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.990 736.000 1295.270 740.000 ;
    END
  END la_output[100]
  PIN la_output[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.870 736.000 1308.150 740.000 ;
    END
  END la_output[101]
  PIN la_output[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.750 736.000 1321.030 740.000 ;
    END
  END la_output[102]
  PIN la_output[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.630 736.000 1333.910 740.000 ;
    END
  END la_output[103]
  PIN la_output[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.510 736.000 1346.790 740.000 ;
    END
  END la_output[104]
  PIN la_output[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1359.390 736.000 1359.670 740.000 ;
    END
  END la_output[105]
  PIN la_output[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1372.270 736.000 1372.550 740.000 ;
    END
  END la_output[106]
  PIN la_output[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.150 736.000 1385.430 740.000 ;
    END
  END la_output[107]
  PIN la_output[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.570 736.000 1397.850 740.000 ;
    END
  END la_output[108]
  PIN la_output[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1410.450 736.000 1410.730 740.000 ;
    END
  END la_output[109]
  PIN la_output[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 736.000 139.750 740.000 ;
    END
  END la_output[10]
  PIN la_output[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.330 736.000 1423.610 740.000 ;
    END
  END la_output[110]
  PIN la_output[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.210 736.000 1436.490 740.000 ;
    END
  END la_output[111]
  PIN la_output[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1449.090 736.000 1449.370 740.000 ;
    END
  END la_output[112]
  PIN la_output[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.970 736.000 1462.250 740.000 ;
    END
  END la_output[113]
  PIN la_output[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.850 736.000 1475.130 740.000 ;
    END
  END la_output[114]
  PIN la_output[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1487.730 736.000 1488.010 740.000 ;
    END
  END la_output[115]
  PIN la_output[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.610 736.000 1500.890 740.000 ;
    END
  END la_output[116]
  PIN la_output[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.490 736.000 1513.770 740.000 ;
    END
  END la_output[117]
  PIN la_output[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.370 736.000 1526.650 740.000 ;
    END
  END la_output[118]
  PIN la_output[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.250 736.000 1539.530 740.000 ;
    END
  END la_output[119]
  PIN la_output[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 736.000 152.630 740.000 ;
    END
  END la_output[11]
  PIN la_output[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.670 736.000 1551.950 740.000 ;
    END
  END la_output[120]
  PIN la_output[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1564.550 736.000 1564.830 740.000 ;
    END
  END la_output[121]
  PIN la_output[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1577.430 736.000 1577.710 740.000 ;
    END
  END la_output[122]
  PIN la_output[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1590.310 736.000 1590.590 740.000 ;
    END
  END la_output[123]
  PIN la_output[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.190 736.000 1603.470 740.000 ;
    END
  END la_output[124]
  PIN la_output[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.070 736.000 1616.350 740.000 ;
    END
  END la_output[125]
  PIN la_output[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1628.950 736.000 1629.230 740.000 ;
    END
  END la_output[126]
  PIN la_output[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1641.830 736.000 1642.110 740.000 ;
    END
  END la_output[127]
  PIN la_output[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 736.000 165.050 740.000 ;
    END
  END la_output[12]
  PIN la_output[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 736.000 177.930 740.000 ;
    END
  END la_output[13]
  PIN la_output[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.530 736.000 190.810 740.000 ;
    END
  END la_output[14]
  PIN la_output[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.410 736.000 203.690 740.000 ;
    END
  END la_output[15]
  PIN la_output[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 736.000 216.570 740.000 ;
    END
  END la_output[16]
  PIN la_output[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 736.000 229.450 740.000 ;
    END
  END la_output[17]
  PIN la_output[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 736.000 242.330 740.000 ;
    END
  END la_output[18]
  PIN la_output[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 736.000 255.210 740.000 ;
    END
  END la_output[19]
  PIN la_output[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 736.000 23.830 740.000 ;
    END
  END la_output[1]
  PIN la_output[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 736.000 268.090 740.000 ;
    END
  END la_output[20]
  PIN la_output[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 736.000 280.970 740.000 ;
    END
  END la_output[21]
  PIN la_output[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 736.000 293.850 740.000 ;
    END
  END la_output[22]
  PIN la_output[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.450 736.000 306.730 740.000 ;
    END
  END la_output[23]
  PIN la_output[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 736.000 319.150 740.000 ;
    END
  END la_output[24]
  PIN la_output[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 736.000 332.030 740.000 ;
    END
  END la_output[25]
  PIN la_output[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 736.000 344.910 740.000 ;
    END
  END la_output[26]
  PIN la_output[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 736.000 357.790 740.000 ;
    END
  END la_output[27]
  PIN la_output[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 736.000 370.670 740.000 ;
    END
  END la_output[28]
  PIN la_output[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 736.000 383.550 740.000 ;
    END
  END la_output[29]
  PIN la_output[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 736.000 36.710 740.000 ;
    END
  END la_output[2]
  PIN la_output[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 736.000 396.430 740.000 ;
    END
  END la_output[30]
  PIN la_output[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 736.000 409.310 740.000 ;
    END
  END la_output[31]
  PIN la_output[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 736.000 422.190 740.000 ;
    END
  END la_output[32]
  PIN la_output[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 736.000 435.070 740.000 ;
    END
  END la_output[33]
  PIN la_output[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 736.000 447.950 740.000 ;
    END
  END la_output[34]
  PIN la_output[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 736.000 460.830 740.000 ;
    END
  END la_output[35]
  PIN la_output[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 736.000 473.250 740.000 ;
    END
  END la_output[36]
  PIN la_output[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 736.000 486.130 740.000 ;
    END
  END la_output[37]
  PIN la_output[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 736.000 499.010 740.000 ;
    END
  END la_output[38]
  PIN la_output[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.610 736.000 511.890 740.000 ;
    END
  END la_output[39]
  PIN la_output[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 736.000 49.590 740.000 ;
    END
  END la_output[3]
  PIN la_output[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.490 736.000 524.770 740.000 ;
    END
  END la_output[40]
  PIN la_output[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.370 736.000 537.650 740.000 ;
    END
  END la_output[41]
  PIN la_output[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.250 736.000 550.530 740.000 ;
    END
  END la_output[42]
  PIN la_output[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.130 736.000 563.410 740.000 ;
    END
  END la_output[43]
  PIN la_output[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 736.000 576.290 740.000 ;
    END
  END la_output[44]
  PIN la_output[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.890 736.000 589.170 740.000 ;
    END
  END la_output[45]
  PIN la_output[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.770 736.000 602.050 740.000 ;
    END
  END la_output[46]
  PIN la_output[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.650 736.000 614.930 740.000 ;
    END
  END la_output[47]
  PIN la_output[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.070 736.000 627.350 740.000 ;
    END
  END la_output[48]
  PIN la_output[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.950 736.000 640.230 740.000 ;
    END
  END la_output[49]
  PIN la_output[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.190 736.000 62.470 740.000 ;
    END
  END la_output[4]
  PIN la_output[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 736.000 653.110 740.000 ;
    END
  END la_output[50]
  PIN la_output[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.710 736.000 665.990 740.000 ;
    END
  END la_output[51]
  PIN la_output[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.590 736.000 678.870 740.000 ;
    END
  END la_output[52]
  PIN la_output[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.470 736.000 691.750 740.000 ;
    END
  END la_output[53]
  PIN la_output[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 704.350 736.000 704.630 740.000 ;
    END
  END la_output[54]
  PIN la_output[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.230 736.000 717.510 740.000 ;
    END
  END la_output[55]
  PIN la_output[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 736.000 730.390 740.000 ;
    END
  END la_output[56]
  PIN la_output[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.990 736.000 743.270 740.000 ;
    END
  END la_output[57]
  PIN la_output[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.870 736.000 756.150 740.000 ;
    END
  END la_output[58]
  PIN la_output[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 736.000 769.030 740.000 ;
    END
  END la_output[59]
  PIN la_output[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.070 736.000 75.350 740.000 ;
    END
  END la_output[5]
  PIN la_output[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 736.000 781.450 740.000 ;
    END
  END la_output[60]
  PIN la_output[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.050 736.000 794.330 740.000 ;
    END
  END la_output[61]
  PIN la_output[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.930 736.000 807.210 740.000 ;
    END
  END la_output[62]
  PIN la_output[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.810 736.000 820.090 740.000 ;
    END
  END la_output[63]
  PIN la_output[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.690 736.000 832.970 740.000 ;
    END
  END la_output[64]
  PIN la_output[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.570 736.000 845.850 740.000 ;
    END
  END la_output[65]
  PIN la_output[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.450 736.000 858.730 740.000 ;
    END
  END la_output[66]
  PIN la_output[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.330 736.000 871.610 740.000 ;
    END
  END la_output[67]
  PIN la_output[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.210 736.000 884.490 740.000 ;
    END
  END la_output[68]
  PIN la_output[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 897.090 736.000 897.370 740.000 ;
    END
  END la_output[69]
  PIN la_output[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 736.000 88.230 740.000 ;
    END
  END la_output[6]
  PIN la_output[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.970 736.000 910.250 740.000 ;
    END
  END la_output[70]
  PIN la_output[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.850 736.000 923.130 740.000 ;
    END
  END la_output[71]
  PIN la_output[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 935.270 736.000 935.550 740.000 ;
    END
  END la_output[72]
  PIN la_output[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.150 736.000 948.430 740.000 ;
    END
  END la_output[73]
  PIN la_output[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.030 736.000 961.310 740.000 ;
    END
  END la_output[74]
  PIN la_output[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 973.910 736.000 974.190 740.000 ;
    END
  END la_output[75]
  PIN la_output[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.790 736.000 987.070 740.000 ;
    END
  END la_output[76]
  PIN la_output[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.670 736.000 999.950 740.000 ;
    END
  END la_output[77]
  PIN la_output[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.550 736.000 1012.830 740.000 ;
    END
  END la_output[78]
  PIN la_output[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.430 736.000 1025.710 740.000 ;
    END
  END la_output[79]
  PIN la_output[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 736.000 101.110 740.000 ;
    END
  END la_output[7]
  PIN la_output[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1038.310 736.000 1038.590 740.000 ;
    END
  END la_output[80]
  PIN la_output[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.190 736.000 1051.470 740.000 ;
    END
  END la_output[81]
  PIN la_output[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.070 736.000 1064.350 740.000 ;
    END
  END la_output[82]
  PIN la_output[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.950 736.000 1077.230 740.000 ;
    END
  END la_output[83]
  PIN la_output[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1089.370 736.000 1089.650 740.000 ;
    END
  END la_output[84]
  PIN la_output[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.250 736.000 1102.530 740.000 ;
    END
  END la_output[85]
  PIN la_output[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1115.130 736.000 1115.410 740.000 ;
    END
  END la_output[86]
  PIN la_output[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.010 736.000 1128.290 740.000 ;
    END
  END la_output[87]
  PIN la_output[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1140.890 736.000 1141.170 740.000 ;
    END
  END la_output[88]
  PIN la_output[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1153.770 736.000 1154.050 740.000 ;
    END
  END la_output[89]
  PIN la_output[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.710 736.000 113.990 740.000 ;
    END
  END la_output[8]
  PIN la_output[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.650 736.000 1166.930 740.000 ;
    END
  END la_output[90]
  PIN la_output[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.530 736.000 1179.810 740.000 ;
    END
  END la_output[91]
  PIN la_output[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1192.410 736.000 1192.690 740.000 ;
    END
  END la_output[92]
  PIN la_output[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.290 736.000 1205.570 740.000 ;
    END
  END la_output[93]
  PIN la_output[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.170 736.000 1218.450 740.000 ;
    END
  END la_output[94]
  PIN la_output[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.050 736.000 1231.330 740.000 ;
    END
  END la_output[95]
  PIN la_output[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.470 736.000 1243.750 740.000 ;
    END
  END la_output[96]
  PIN la_output[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1256.350 736.000 1256.630 740.000 ;
    END
  END la_output[97]
  PIN la_output[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.230 736.000 1269.510 740.000 ;
    END
  END la_output[98]
  PIN la_output[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1282.110 736.000 1282.390 740.000 ;
    END
  END la_output[99]
  PIN la_output[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 736.000 126.870 740.000 ;
    END
  END la_output[9]
  PIN mgmt_soc_dff_A[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END mgmt_soc_dff_A[0]
  PIN mgmt_soc_dff_A[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.680 4.000 322.280 ;
    END
  END mgmt_soc_dff_A[1]
  PIN mgmt_soc_dff_A[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.200 4.000 331.800 ;
    END
  END mgmt_soc_dff_A[2]
  PIN mgmt_soc_dff_A[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END mgmt_soc_dff_A[3]
  PIN mgmt_soc_dff_A[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END mgmt_soc_dff_A[4]
  PIN mgmt_soc_dff_A[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.760 4.000 360.360 ;
    END
  END mgmt_soc_dff_A[5]
  PIN mgmt_soc_dff_A[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.280 4.000 369.880 ;
    END
  END mgmt_soc_dff_A[6]
  PIN mgmt_soc_dff_A[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END mgmt_soc_dff_A[7]
  PIN mgmt_soc_dff_Di[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.800 4.000 5.400 ;
    END
  END mgmt_soc_dff_Di[0]
  PIN mgmt_soc_dff_Di[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END mgmt_soc_dff_Di[10]
  PIN mgmt_soc_dff_Di[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END mgmt_soc_dff_Di[11]
  PIN mgmt_soc_dff_Di[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END mgmt_soc_dff_Di[12]
  PIN mgmt_soc_dff_Di[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END mgmt_soc_dff_Di[13]
  PIN mgmt_soc_dff_Di[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END mgmt_soc_dff_Di[14]
  PIN mgmt_soc_dff_Di[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.280 4.000 148.880 ;
    END
  END mgmt_soc_dff_Di[15]
  PIN mgmt_soc_dff_Di[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END mgmt_soc_dff_Di[16]
  PIN mgmt_soc_dff_Di[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END mgmt_soc_dff_Di[17]
  PIN mgmt_soc_dff_Di[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.520 4.000 178.120 ;
    END
  END mgmt_soc_dff_Di[18]
  PIN mgmt_soc_dff_Di[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END mgmt_soc_dff_Di[19]
  PIN mgmt_soc_dff_Di[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 14.320 4.000 14.920 ;
    END
  END mgmt_soc_dff_Di[1]
  PIN mgmt_soc_dff_Di[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END mgmt_soc_dff_Di[20]
  PIN mgmt_soc_dff_Di[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.080 4.000 206.680 ;
    END
  END mgmt_soc_dff_Di[21]
  PIN mgmt_soc_dff_Di[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 215.600 4.000 216.200 ;
    END
  END mgmt_soc_dff_Di[22]
  PIN mgmt_soc_dff_Di[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END mgmt_soc_dff_Di[23]
  PIN mgmt_soc_dff_Di[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END mgmt_soc_dff_Di[24]
  PIN mgmt_soc_dff_Di[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END mgmt_soc_dff_Di[25]
  PIN mgmt_soc_dff_Di[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END mgmt_soc_dff_Di[26]
  PIN mgmt_soc_dff_Di[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 263.880 4.000 264.480 ;
    END
  END mgmt_soc_dff_Di[27]
  PIN mgmt_soc_dff_Di[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 273.400 4.000 274.000 ;
    END
  END mgmt_soc_dff_Di[28]
  PIN mgmt_soc_dff_Di[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.920 4.000 283.520 ;
    END
  END mgmt_soc_dff_Di[29]
  PIN mgmt_soc_dff_Di[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END mgmt_soc_dff_Di[2]
  PIN mgmt_soc_dff_Di[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END mgmt_soc_dff_Di[30]
  PIN mgmt_soc_dff_Di[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END mgmt_soc_dff_Di[31]
  PIN mgmt_soc_dff_Di[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END mgmt_soc_dff_Di[3]
  PIN mgmt_soc_dff_Di[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END mgmt_soc_dff_Di[4]
  PIN mgmt_soc_dff_Di[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END mgmt_soc_dff_Di[5]
  PIN mgmt_soc_dff_Di[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END mgmt_soc_dff_Di[6]
  PIN mgmt_soc_dff_Di[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END mgmt_soc_dff_Di[7]
  PIN mgmt_soc_dff_Di[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END mgmt_soc_dff_Di[8]
  PIN mgmt_soc_dff_Di[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END mgmt_soc_dff_Di[9]
  PIN mgmt_soc_dff_Do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END mgmt_soc_dff_Do[0]
  PIN mgmt_soc_dff_Do[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.160 4.000 533.760 ;
    END
  END mgmt_soc_dff_Do[10]
  PIN mgmt_soc_dff_Do[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 4.000 543.280 ;
    END
  END mgmt_soc_dff_Do[11]
  PIN mgmt_soc_dff_Do[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END mgmt_soc_dff_Do[12]
  PIN mgmt_soc_dff_Do[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 561.720 4.000 562.320 ;
    END
  END mgmt_soc_dff_Do[13]
  PIN mgmt_soc_dff_Do[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END mgmt_soc_dff_Do[14]
  PIN mgmt_soc_dff_Do[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 580.760 4.000 581.360 ;
    END
  END mgmt_soc_dff_Do[15]
  PIN mgmt_soc_dff_Do[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 590.280 4.000 590.880 ;
    END
  END mgmt_soc_dff_Do[16]
  PIN mgmt_soc_dff_Do[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 600.480 4.000 601.080 ;
    END
  END mgmt_soc_dff_Do[17]
  PIN mgmt_soc_dff_Do[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.000 4.000 610.600 ;
    END
  END mgmt_soc_dff_Do[18]
  PIN mgmt_soc_dff_Do[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 619.520 4.000 620.120 ;
    END
  END mgmt_soc_dff_Do[19]
  PIN mgmt_soc_dff_Do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.120 4.000 446.720 ;
    END
  END mgmt_soc_dff_Do[1]
  PIN mgmt_soc_dff_Do[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 629.040 4.000 629.640 ;
    END
  END mgmt_soc_dff_Do[20]
  PIN mgmt_soc_dff_Do[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 638.560 4.000 639.160 ;
    END
  END mgmt_soc_dff_Do[21]
  PIN mgmt_soc_dff_Do[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.080 4.000 648.680 ;
    END
  END mgmt_soc_dff_Do[22]
  PIN mgmt_soc_dff_Do[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 657.600 4.000 658.200 ;
    END
  END mgmt_soc_dff_Do[23]
  PIN mgmt_soc_dff_Do[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.120 4.000 667.720 ;
    END
  END mgmt_soc_dff_Do[24]
  PIN mgmt_soc_dff_Do[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 677.320 4.000 677.920 ;
    END
  END mgmt_soc_dff_Do[25]
  PIN mgmt_soc_dff_Do[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.840 4.000 687.440 ;
    END
  END mgmt_soc_dff_Do[26]
  PIN mgmt_soc_dff_Do[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 696.360 4.000 696.960 ;
    END
  END mgmt_soc_dff_Do[27]
  PIN mgmt_soc_dff_Do[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 4.000 706.480 ;
    END
  END mgmt_soc_dff_Do[28]
  PIN mgmt_soc_dff_Do[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 715.400 4.000 716.000 ;
    END
  END mgmt_soc_dff_Do[29]
  PIN mgmt_soc_dff_Do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 456.320 4.000 456.920 ;
    END
  END mgmt_soc_dff_Do[2]
  PIN mgmt_soc_dff_Do[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 724.920 4.000 725.520 ;
    END
  END mgmt_soc_dff_Do[30]
  PIN mgmt_soc_dff_Do[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END mgmt_soc_dff_Do[31]
  PIN mgmt_soc_dff_Do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END mgmt_soc_dff_Do[3]
  PIN mgmt_soc_dff_Do[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 475.360 4.000 475.960 ;
    END
  END mgmt_soc_dff_Do[4]
  PIN mgmt_soc_dff_Do[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.880 4.000 485.480 ;
    END
  END mgmt_soc_dff_Do[5]
  PIN mgmt_soc_dff_Do[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 494.400 4.000 495.000 ;
    END
  END mgmt_soc_dff_Do[6]
  PIN mgmt_soc_dff_Do[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.920 4.000 504.520 ;
    END
  END mgmt_soc_dff_Do[7]
  PIN mgmt_soc_dff_Do[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 4.000 514.040 ;
    END
  END mgmt_soc_dff_Do[8]
  PIN mgmt_soc_dff_Do[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END mgmt_soc_dff_Do[9]
  PIN mgmt_soc_dff_EN
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END mgmt_soc_dff_EN
  PIN mgmt_soc_dff_WE[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END mgmt_soc_dff_WE[0]
  PIN mgmt_soc_dff_WE[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 398.520 4.000 399.120 ;
    END
  END mgmt_soc_dff_WE[1]
  PIN mgmt_soc_dff_WE[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.040 4.000 408.640 ;
    END
  END mgmt_soc_dff_WE[2]
  PIN mgmt_soc_dff_WE[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END mgmt_soc_dff_WE[3]
  PIN mprj_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.050 736.000 1645.330 740.000 ;
    END
  END mprj_ack_i
  PIN mprj_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.150 736.000 1661.430 740.000 ;
    END
  END mprj_adr_o[0]
  PIN mprj_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.170 736.000 1770.450 740.000 ;
    END
  END mprj_adr_o[10]
  PIN mprj_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1779.830 736.000 1780.110 740.000 ;
    END
  END mprj_adr_o[11]
  PIN mprj_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1789.490 736.000 1789.770 740.000 ;
    END
  END mprj_adr_o[12]
  PIN mprj_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.150 736.000 1799.430 740.000 ;
    END
  END mprj_adr_o[13]
  PIN mprj_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1808.810 736.000 1809.090 740.000 ;
    END
  END mprj_adr_o[14]
  PIN mprj_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1818.470 736.000 1818.750 740.000 ;
    END
  END mprj_adr_o[15]
  PIN mprj_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.130 736.000 1828.410 740.000 ;
    END
  END mprj_adr_o[16]
  PIN mprj_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1837.790 736.000 1838.070 740.000 ;
    END
  END mprj_adr_o[17]
  PIN mprj_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1847.450 736.000 1847.730 740.000 ;
    END
  END mprj_adr_o[18]
  PIN mprj_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1856.650 736.000 1856.930 740.000 ;
    END
  END mprj_adr_o[19]
  PIN mprj_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.030 736.000 1674.310 740.000 ;
    END
  END mprj_adr_o[1]
  PIN mprj_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1866.310 736.000 1866.590 740.000 ;
    END
  END mprj_adr_o[20]
  PIN mprj_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1875.970 736.000 1876.250 740.000 ;
    END
  END mprj_adr_o[21]
  PIN mprj_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1885.630 736.000 1885.910 740.000 ;
    END
  END mprj_adr_o[22]
  PIN mprj_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1895.290 736.000 1895.570 740.000 ;
    END
  END mprj_adr_o[23]
  PIN mprj_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.950 736.000 1905.230 740.000 ;
    END
  END mprj_adr_o[24]
  PIN mprj_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1914.610 736.000 1914.890 740.000 ;
    END
  END mprj_adr_o[25]
  PIN mprj_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1924.270 736.000 1924.550 740.000 ;
    END
  END mprj_adr_o[26]
  PIN mprj_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1933.930 736.000 1934.210 740.000 ;
    END
  END mprj_adr_o[27]
  PIN mprj_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1943.590 736.000 1943.870 740.000 ;
    END
  END mprj_adr_o[28]
  PIN mprj_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.250 736.000 1953.530 740.000 ;
    END
  END mprj_adr_o[29]
  PIN mprj_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1686.910 736.000 1687.190 740.000 ;
    END
  END mprj_adr_o[2]
  PIN mprj_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1962.910 736.000 1963.190 740.000 ;
    END
  END mprj_adr_o[30]
  PIN mprj_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1972.570 736.000 1972.850 740.000 ;
    END
  END mprj_adr_o[31]
  PIN mprj_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.330 736.000 1699.610 740.000 ;
    END
  END mprj_adr_o[3]
  PIN mprj_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1712.210 736.000 1712.490 740.000 ;
    END
  END mprj_adr_o[4]
  PIN mprj_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.870 736.000 1722.150 740.000 ;
    END
  END mprj_adr_o[5]
  PIN mprj_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1731.530 736.000 1731.810 740.000 ;
    END
  END mprj_adr_o[6]
  PIN mprj_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1741.190 736.000 1741.470 740.000 ;
    END
  END mprj_adr_o[7]
  PIN mprj_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1750.850 736.000 1751.130 740.000 ;
    END
  END mprj_adr_o[8]
  PIN mprj_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.510 736.000 1760.790 740.000 ;
    END
  END mprj_adr_o[9]
  PIN mprj_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1648.270 736.000 1648.550 740.000 ;
    END
  END mprj_cyc_o
  PIN mprj_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1664.370 736.000 1664.650 740.000 ;
    END
  END mprj_dat_i[0]
  PIN mprj_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1773.390 736.000 1773.670 740.000 ;
    END
  END mprj_dat_i[10]
  PIN mprj_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.050 736.000 1783.330 740.000 ;
    END
  END mprj_dat_i[11]
  PIN mprj_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1792.710 736.000 1792.990 740.000 ;
    END
  END mprj_dat_i[12]
  PIN mprj_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1802.370 736.000 1802.650 740.000 ;
    END
  END mprj_dat_i[13]
  PIN mprj_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1812.030 736.000 1812.310 740.000 ;
    END
  END mprj_dat_i[14]
  PIN mprj_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1821.690 736.000 1821.970 740.000 ;
    END
  END mprj_dat_i[15]
  PIN mprj_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1831.350 736.000 1831.630 740.000 ;
    END
  END mprj_dat_i[16]
  PIN mprj_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.010 736.000 1841.290 740.000 ;
    END
  END mprj_dat_i[17]
  PIN mprj_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1850.210 736.000 1850.490 740.000 ;
    END
  END mprj_dat_i[18]
  PIN mprj_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1859.870 736.000 1860.150 740.000 ;
    END
  END mprj_dat_i[19]
  PIN mprj_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1677.250 736.000 1677.530 740.000 ;
    END
  END mprj_dat_i[1]
  PIN mprj_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1869.530 736.000 1869.810 740.000 ;
    END
  END mprj_dat_i[20]
  PIN mprj_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1879.190 736.000 1879.470 740.000 ;
    END
  END mprj_dat_i[21]
  PIN mprj_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.850 736.000 1889.130 740.000 ;
    END
  END mprj_dat_i[22]
  PIN mprj_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1898.510 736.000 1898.790 740.000 ;
    END
  END mprj_dat_i[23]
  PIN mprj_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1908.170 736.000 1908.450 740.000 ;
    END
  END mprj_dat_i[24]
  PIN mprj_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.830 736.000 1918.110 740.000 ;
    END
  END mprj_dat_i[25]
  PIN mprj_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1927.490 736.000 1927.770 740.000 ;
    END
  END mprj_dat_i[26]
  PIN mprj_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1937.150 736.000 1937.430 740.000 ;
    END
  END mprj_dat_i[27]
  PIN mprj_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1946.810 736.000 1947.090 740.000 ;
    END
  END mprj_dat_i[28]
  PIN mprj_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1956.470 736.000 1956.750 740.000 ;
    END
  END mprj_dat_i[29]
  PIN mprj_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1690.130 736.000 1690.410 740.000 ;
    END
  END mprj_dat_i[2]
  PIN mprj_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1966.130 736.000 1966.410 740.000 ;
    END
  END mprj_dat_i[30]
  PIN mprj_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1975.790 736.000 1976.070 740.000 ;
    END
  END mprj_dat_i[31]
  PIN mprj_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1702.550 736.000 1702.830 740.000 ;
    END
  END mprj_dat_i[3]
  PIN mprj_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.430 736.000 1715.710 740.000 ;
    END
  END mprj_dat_i[4]
  PIN mprj_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1725.090 736.000 1725.370 740.000 ;
    END
  END mprj_dat_i[5]
  PIN mprj_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.750 736.000 1735.030 740.000 ;
    END
  END mprj_dat_i[6]
  PIN mprj_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1744.410 736.000 1744.690 740.000 ;
    END
  END mprj_dat_i[7]
  PIN mprj_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.070 736.000 1754.350 740.000 ;
    END
  END mprj_dat_i[8]
  PIN mprj_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1763.730 736.000 1764.010 740.000 ;
    END
  END mprj_dat_i[9]
  PIN mprj_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1667.590 736.000 1667.870 740.000 ;
    END
  END mprj_dat_o[0]
  PIN mprj_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.610 736.000 1776.890 740.000 ;
    END
  END mprj_dat_o[10]
  PIN mprj_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1786.270 736.000 1786.550 740.000 ;
    END
  END mprj_dat_o[11]
  PIN mprj_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1795.930 736.000 1796.210 740.000 ;
    END
  END mprj_dat_o[12]
  PIN mprj_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.590 736.000 1805.870 740.000 ;
    END
  END mprj_dat_o[13]
  PIN mprj_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1815.250 736.000 1815.530 740.000 ;
    END
  END mprj_dat_o[14]
  PIN mprj_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.910 736.000 1825.190 740.000 ;
    END
  END mprj_dat_o[15]
  PIN mprj_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.570 736.000 1834.850 740.000 ;
    END
  END mprj_dat_o[16]
  PIN mprj_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1844.230 736.000 1844.510 740.000 ;
    END
  END mprj_dat_o[17]
  PIN mprj_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1853.430 736.000 1853.710 740.000 ;
    END
  END mprj_dat_o[18]
  PIN mprj_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1863.090 736.000 1863.370 740.000 ;
    END
  END mprj_dat_o[19]
  PIN mprj_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.470 736.000 1680.750 740.000 ;
    END
  END mprj_dat_o[1]
  PIN mprj_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1872.750 736.000 1873.030 740.000 ;
    END
  END mprj_dat_o[20]
  PIN mprj_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.410 736.000 1882.690 740.000 ;
    END
  END mprj_dat_o[21]
  PIN mprj_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1892.070 736.000 1892.350 740.000 ;
    END
  END mprj_dat_o[22]
  PIN mprj_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1901.730 736.000 1902.010 740.000 ;
    END
  END mprj_dat_o[23]
  PIN mprj_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.390 736.000 1911.670 740.000 ;
    END
  END mprj_dat_o[24]
  PIN mprj_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1921.050 736.000 1921.330 740.000 ;
    END
  END mprj_dat_o[25]
  PIN mprj_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1930.710 736.000 1930.990 740.000 ;
    END
  END mprj_dat_o[26]
  PIN mprj_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1940.370 736.000 1940.650 740.000 ;
    END
  END mprj_dat_o[27]
  PIN mprj_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1950.030 736.000 1950.310 740.000 ;
    END
  END mprj_dat_o[28]
  PIN mprj_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.690 736.000 1959.970 740.000 ;
    END
  END mprj_dat_o[29]
  PIN mprj_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.350 736.000 1693.630 740.000 ;
    END
  END mprj_dat_o[2]
  PIN mprj_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1969.350 736.000 1969.630 740.000 ;
    END
  END mprj_dat_o[30]
  PIN mprj_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1979.010 736.000 1979.290 740.000 ;
    END
  END mprj_dat_o[31]
  PIN mprj_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1705.770 736.000 1706.050 740.000 ;
    END
  END mprj_dat_o[3]
  PIN mprj_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1718.650 736.000 1718.930 740.000 ;
    END
  END mprj_dat_o[4]
  PIN mprj_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.310 736.000 1728.590 740.000 ;
    END
  END mprj_dat_o[5]
  PIN mprj_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1737.970 736.000 1738.250 740.000 ;
    END
  END mprj_dat_o[6]
  PIN mprj_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1747.630 736.000 1747.910 740.000 ;
    END
  END mprj_dat_o[7]
  PIN mprj_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1757.290 736.000 1757.570 740.000 ;
    END
  END mprj_dat_o[8]
  PIN mprj_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1766.950 736.000 1767.230 740.000 ;
    END
  END mprj_dat_o[9]
  PIN mprj_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1670.810 736.000 1671.090 740.000 ;
    END
  END mprj_sel_o[0]
  PIN mprj_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1683.690 736.000 1683.970 740.000 ;
    END
  END mprj_sel_o[1]
  PIN mprj_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1696.110 736.000 1696.390 740.000 ;
    END
  END mprj_sel_o[2]
  PIN mprj_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1708.990 736.000 1709.270 740.000 ;
    END
  END mprj_sel_o[3]
  PIN mprj_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.490 736.000 1651.770 740.000 ;
    END
  END mprj_stb_o
  PIN mprj_wb_iena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1654.710 736.000 1654.990 740.000 ;
    END
  END mprj_wb_iena
  PIN mprj_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.930 736.000 1658.210 740.000 ;
    END
  END mprj_we_o
  PIN qspi_enabled
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 402.600 2000.000 403.200 ;
    END
  END qspi_enabled
  PIN serial_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 375.400 2000.000 376.000 ;
    END
  END serial_rx
  PIN serial_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 382.200 2000.000 382.800 ;
    END
  END serial_tx
  PIN spi_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 355.680 2000.000 356.280 ;
    END
  END spi_clk
  PIN spi_cs_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 362.480 2000.000 363.080 ;
    END
  END spi_cs_n
  PIN spi_enabled
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 389.000 2000.000 389.600 ;
    END
  END spi_enabled
  PIN spi_miso
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 369.280 2000.000 369.880 ;
    END
  END spi_miso
  PIN spi_mosi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 348.880 2000.000 349.480 ;
    END
  END spi_mosi
  PIN spi_sdoenb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 342.080 2000.000 342.680 ;
    END
  END spi_sdoenb
  PIN sram_ro_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 8.880 2000.000 9.480 ;
    END
  END sram_ro_addr[0]
  PIN sram_ro_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 15.680 2000.000 16.280 ;
    END
  END sram_ro_addr[1]
  PIN sram_ro_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 22.480 2000.000 23.080 ;
    END
  END sram_ro_addr[2]
  PIN sram_ro_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 29.280 2000.000 29.880 ;
    END
  END sram_ro_addr[3]
  PIN sram_ro_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 36.080 2000.000 36.680 ;
    END
  END sram_ro_addr[4]
  PIN sram_ro_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 42.880 2000.000 43.480 ;
    END
  END sram_ro_addr[5]
  PIN sram_ro_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 49.680 2000.000 50.280 ;
    END
  END sram_ro_addr[6]
  PIN sram_ro_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 56.480 2000.000 57.080 ;
    END
  END sram_ro_addr[7]
  PIN sram_ro_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 63.280 2000.000 63.880 ;
    END
  END sram_ro_clk
  PIN sram_ro_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 2.760 2000.000 3.360 ;
    END
  END sram_ro_csb
  PIN sram_ro_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 70.080 2000.000 70.680 ;
    END
  END sram_ro_data[0]
  PIN sram_ro_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 138.080 2000.000 138.680 ;
    END
  END sram_ro_data[10]
  PIN sram_ro_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 144.880 2000.000 145.480 ;
    END
  END sram_ro_data[11]
  PIN sram_ro_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 151.680 2000.000 152.280 ;
    END
  END sram_ro_data[12]
  PIN sram_ro_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 158.480 2000.000 159.080 ;
    END
  END sram_ro_data[13]
  PIN sram_ro_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 165.280 2000.000 165.880 ;
    END
  END sram_ro_data[14]
  PIN sram_ro_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 172.080 2000.000 172.680 ;
    END
  END sram_ro_data[15]
  PIN sram_ro_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 178.880 2000.000 179.480 ;
    END
  END sram_ro_data[16]
  PIN sram_ro_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 185.680 2000.000 186.280 ;
    END
  END sram_ro_data[17]
  PIN sram_ro_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 192.480 2000.000 193.080 ;
    END
  END sram_ro_data[18]
  PIN sram_ro_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 199.280 2000.000 199.880 ;
    END
  END sram_ro_data[19]
  PIN sram_ro_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 76.880 2000.000 77.480 ;
    END
  END sram_ro_data[1]
  PIN sram_ro_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 206.080 2000.000 206.680 ;
    END
  END sram_ro_data[20]
  PIN sram_ro_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 212.880 2000.000 213.480 ;
    END
  END sram_ro_data[21]
  PIN sram_ro_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 219.680 2000.000 220.280 ;
    END
  END sram_ro_data[22]
  PIN sram_ro_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 226.480 2000.000 227.080 ;
    END
  END sram_ro_data[23]
  PIN sram_ro_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 233.280 2000.000 233.880 ;
    END
  END sram_ro_data[24]
  PIN sram_ro_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 240.080 2000.000 240.680 ;
    END
  END sram_ro_data[25]
  PIN sram_ro_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 246.880 2000.000 247.480 ;
    END
  END sram_ro_data[26]
  PIN sram_ro_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 253.680 2000.000 254.280 ;
    END
  END sram_ro_data[27]
  PIN sram_ro_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 260.480 2000.000 261.080 ;
    END
  END sram_ro_data[28]
  PIN sram_ro_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 267.280 2000.000 267.880 ;
    END
  END sram_ro_data[29]
  PIN sram_ro_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 83.680 2000.000 84.280 ;
    END
  END sram_ro_data[2]
  PIN sram_ro_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 274.080 2000.000 274.680 ;
    END
  END sram_ro_data[30]
  PIN sram_ro_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 280.880 2000.000 281.480 ;
    END
  END sram_ro_data[31]
  PIN sram_ro_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 90.480 2000.000 91.080 ;
    END
  END sram_ro_data[3]
  PIN sram_ro_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 97.280 2000.000 97.880 ;
    END
  END sram_ro_data[4]
  PIN sram_ro_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 104.080 2000.000 104.680 ;
    END
  END sram_ro_data[5]
  PIN sram_ro_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 110.880 2000.000 111.480 ;
    END
  END sram_ro_data[6]
  PIN sram_ro_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 117.680 2000.000 118.280 ;
    END
  END sram_ro_data[7]
  PIN sram_ro_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 124.480 2000.000 125.080 ;
    END
  END sram_ro_data[8]
  PIN sram_ro_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 131.280 2000.000 131.880 ;
    END
  END sram_ro_data[9]
  PIN trap
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 314.880 2000.000 315.480 ;
    END
  END trap
  PIN uart_enabled
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 395.800 2000.000 396.400 ;
    END
  END uart_enabled
  PIN user_irq[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1991.890 736.000 1992.170 740.000 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1995.110 736.000 1995.390 740.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1998.330 736.000 1998.610 740.000 ;
    END
  END user_irq[2]
  PIN user_irq[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 335.280 2000.000 335.880 ;
    END
  END user_irq[3]
  PIN user_irq[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 328.480 2000.000 329.080 ;
    END
  END user_irq[4]
  PIN user_irq[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 321.680 2000.000 322.280 ;
    END
  END user_irq[5]
  PIN user_irq_ena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1982.230 736.000 1982.510 740.000 ;
    END
  END user_irq_ena[0]
  PIN user_irq_ena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1985.450 736.000 1985.730 740.000 ;
    END
  END user_irq_ena[1]
  PIN user_irq_ena[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.670 736.000 1988.950 740.000 ;
    END
  END user_irq_ena[2]
  OBS
      LAYER li1 ;
        RECT 10.120 10.795 1989.500 729.045 ;
      LAYER met1 ;
        RECT 1.450 7.860 1998.630 734.020 ;
      LAYER met2 ;
        RECT 2.030 735.720 3.950 736.285 ;
        RECT 4.790 735.720 7.170 736.285 ;
        RECT 8.010 735.720 10.390 736.285 ;
        RECT 11.230 735.720 13.610 736.285 ;
        RECT 14.450 735.720 16.830 736.285 ;
        RECT 17.670 735.720 20.050 736.285 ;
        RECT 20.890 735.720 23.270 736.285 ;
        RECT 24.110 735.720 26.490 736.285 ;
        RECT 27.330 735.720 29.710 736.285 ;
        RECT 30.550 735.720 32.930 736.285 ;
        RECT 33.770 735.720 36.150 736.285 ;
        RECT 36.990 735.720 39.370 736.285 ;
        RECT 40.210 735.720 42.590 736.285 ;
        RECT 43.430 735.720 45.810 736.285 ;
        RECT 46.650 735.720 49.030 736.285 ;
        RECT 49.870 735.720 52.250 736.285 ;
        RECT 53.090 735.720 55.470 736.285 ;
        RECT 56.310 735.720 58.690 736.285 ;
        RECT 59.530 735.720 61.910 736.285 ;
        RECT 62.750 735.720 65.130 736.285 ;
        RECT 65.970 735.720 68.350 736.285 ;
        RECT 69.190 735.720 71.570 736.285 ;
        RECT 72.410 735.720 74.790 736.285 ;
        RECT 75.630 735.720 78.010 736.285 ;
        RECT 78.850 735.720 81.230 736.285 ;
        RECT 82.070 735.720 84.450 736.285 ;
        RECT 85.290 735.720 87.670 736.285 ;
        RECT 88.510 735.720 90.890 736.285 ;
        RECT 91.730 735.720 94.110 736.285 ;
        RECT 94.950 735.720 97.330 736.285 ;
        RECT 98.170 735.720 100.550 736.285 ;
        RECT 101.390 735.720 103.770 736.285 ;
        RECT 104.610 735.720 106.990 736.285 ;
        RECT 107.830 735.720 110.210 736.285 ;
        RECT 111.050 735.720 113.430 736.285 ;
        RECT 114.270 735.720 116.650 736.285 ;
        RECT 117.490 735.720 119.870 736.285 ;
        RECT 120.710 735.720 123.090 736.285 ;
        RECT 123.930 735.720 126.310 736.285 ;
        RECT 127.150 735.720 129.530 736.285 ;
        RECT 130.370 735.720 132.750 736.285 ;
        RECT 133.590 735.720 135.970 736.285 ;
        RECT 136.810 735.720 139.190 736.285 ;
        RECT 140.030 735.720 142.410 736.285 ;
        RECT 143.250 735.720 145.630 736.285 ;
        RECT 146.470 735.720 148.850 736.285 ;
        RECT 149.690 735.720 152.070 736.285 ;
        RECT 152.910 735.720 154.830 736.285 ;
        RECT 155.670 735.720 158.050 736.285 ;
        RECT 158.890 735.720 161.270 736.285 ;
        RECT 162.110 735.720 164.490 736.285 ;
        RECT 165.330 735.720 167.710 736.285 ;
        RECT 168.550 735.720 170.930 736.285 ;
        RECT 171.770 735.720 174.150 736.285 ;
        RECT 174.990 735.720 177.370 736.285 ;
        RECT 178.210 735.720 180.590 736.285 ;
        RECT 181.430 735.720 183.810 736.285 ;
        RECT 184.650 735.720 187.030 736.285 ;
        RECT 187.870 735.720 190.250 736.285 ;
        RECT 191.090 735.720 193.470 736.285 ;
        RECT 194.310 735.720 196.690 736.285 ;
        RECT 197.530 735.720 199.910 736.285 ;
        RECT 200.750 735.720 203.130 736.285 ;
        RECT 203.970 735.720 206.350 736.285 ;
        RECT 207.190 735.720 209.570 736.285 ;
        RECT 210.410 735.720 212.790 736.285 ;
        RECT 213.630 735.720 216.010 736.285 ;
        RECT 216.850 735.720 219.230 736.285 ;
        RECT 220.070 735.720 222.450 736.285 ;
        RECT 223.290 735.720 225.670 736.285 ;
        RECT 226.510 735.720 228.890 736.285 ;
        RECT 229.730 735.720 232.110 736.285 ;
        RECT 232.950 735.720 235.330 736.285 ;
        RECT 236.170 735.720 238.550 736.285 ;
        RECT 239.390 735.720 241.770 736.285 ;
        RECT 242.610 735.720 244.990 736.285 ;
        RECT 245.830 735.720 248.210 736.285 ;
        RECT 249.050 735.720 251.430 736.285 ;
        RECT 252.270 735.720 254.650 736.285 ;
        RECT 255.490 735.720 257.870 736.285 ;
        RECT 258.710 735.720 261.090 736.285 ;
        RECT 261.930 735.720 264.310 736.285 ;
        RECT 265.150 735.720 267.530 736.285 ;
        RECT 268.370 735.720 270.750 736.285 ;
        RECT 271.590 735.720 273.970 736.285 ;
        RECT 274.810 735.720 277.190 736.285 ;
        RECT 278.030 735.720 280.410 736.285 ;
        RECT 281.250 735.720 283.630 736.285 ;
        RECT 284.470 735.720 286.850 736.285 ;
        RECT 287.690 735.720 290.070 736.285 ;
        RECT 290.910 735.720 293.290 736.285 ;
        RECT 294.130 735.720 296.510 736.285 ;
        RECT 297.350 735.720 299.730 736.285 ;
        RECT 300.570 735.720 302.950 736.285 ;
        RECT 303.790 735.720 306.170 736.285 ;
        RECT 307.010 735.720 308.930 736.285 ;
        RECT 309.770 735.720 312.150 736.285 ;
        RECT 312.990 735.720 315.370 736.285 ;
        RECT 316.210 735.720 318.590 736.285 ;
        RECT 319.430 735.720 321.810 736.285 ;
        RECT 322.650 735.720 325.030 736.285 ;
        RECT 325.870 735.720 328.250 736.285 ;
        RECT 329.090 735.720 331.470 736.285 ;
        RECT 332.310 735.720 334.690 736.285 ;
        RECT 335.530 735.720 337.910 736.285 ;
        RECT 338.750 735.720 341.130 736.285 ;
        RECT 341.970 735.720 344.350 736.285 ;
        RECT 345.190 735.720 347.570 736.285 ;
        RECT 348.410 735.720 350.790 736.285 ;
        RECT 351.630 735.720 354.010 736.285 ;
        RECT 354.850 735.720 357.230 736.285 ;
        RECT 358.070 735.720 360.450 736.285 ;
        RECT 361.290 735.720 363.670 736.285 ;
        RECT 364.510 735.720 366.890 736.285 ;
        RECT 367.730 735.720 370.110 736.285 ;
        RECT 370.950 735.720 373.330 736.285 ;
        RECT 374.170 735.720 376.550 736.285 ;
        RECT 377.390 735.720 379.770 736.285 ;
        RECT 380.610 735.720 382.990 736.285 ;
        RECT 383.830 735.720 386.210 736.285 ;
        RECT 387.050 735.720 389.430 736.285 ;
        RECT 390.270 735.720 392.650 736.285 ;
        RECT 393.490 735.720 395.870 736.285 ;
        RECT 396.710 735.720 399.090 736.285 ;
        RECT 399.930 735.720 402.310 736.285 ;
        RECT 403.150 735.720 405.530 736.285 ;
        RECT 406.370 735.720 408.750 736.285 ;
        RECT 409.590 735.720 411.970 736.285 ;
        RECT 412.810 735.720 415.190 736.285 ;
        RECT 416.030 735.720 418.410 736.285 ;
        RECT 419.250 735.720 421.630 736.285 ;
        RECT 422.470 735.720 424.850 736.285 ;
        RECT 425.690 735.720 428.070 736.285 ;
        RECT 428.910 735.720 431.290 736.285 ;
        RECT 432.130 735.720 434.510 736.285 ;
        RECT 435.350 735.720 437.730 736.285 ;
        RECT 438.570 735.720 440.950 736.285 ;
        RECT 441.790 735.720 444.170 736.285 ;
        RECT 445.010 735.720 447.390 736.285 ;
        RECT 448.230 735.720 450.610 736.285 ;
        RECT 451.450 735.720 453.830 736.285 ;
        RECT 454.670 735.720 457.050 736.285 ;
        RECT 457.890 735.720 460.270 736.285 ;
        RECT 461.110 735.720 463.030 736.285 ;
        RECT 463.870 735.720 466.250 736.285 ;
        RECT 467.090 735.720 469.470 736.285 ;
        RECT 470.310 735.720 472.690 736.285 ;
        RECT 473.530 735.720 475.910 736.285 ;
        RECT 476.750 735.720 479.130 736.285 ;
        RECT 479.970 735.720 482.350 736.285 ;
        RECT 483.190 735.720 485.570 736.285 ;
        RECT 486.410 735.720 488.790 736.285 ;
        RECT 489.630 735.720 492.010 736.285 ;
        RECT 492.850 735.720 495.230 736.285 ;
        RECT 496.070 735.720 498.450 736.285 ;
        RECT 499.290 735.720 501.670 736.285 ;
        RECT 502.510 735.720 504.890 736.285 ;
        RECT 505.730 735.720 508.110 736.285 ;
        RECT 508.950 735.720 511.330 736.285 ;
        RECT 512.170 735.720 514.550 736.285 ;
        RECT 515.390 735.720 517.770 736.285 ;
        RECT 518.610 735.720 520.990 736.285 ;
        RECT 521.830 735.720 524.210 736.285 ;
        RECT 525.050 735.720 527.430 736.285 ;
        RECT 528.270 735.720 530.650 736.285 ;
        RECT 531.490 735.720 533.870 736.285 ;
        RECT 534.710 735.720 537.090 736.285 ;
        RECT 537.930 735.720 540.310 736.285 ;
        RECT 541.150 735.720 543.530 736.285 ;
        RECT 544.370 735.720 546.750 736.285 ;
        RECT 547.590 735.720 549.970 736.285 ;
        RECT 550.810 735.720 553.190 736.285 ;
        RECT 554.030 735.720 556.410 736.285 ;
        RECT 557.250 735.720 559.630 736.285 ;
        RECT 560.470 735.720 562.850 736.285 ;
        RECT 563.690 735.720 566.070 736.285 ;
        RECT 566.910 735.720 569.290 736.285 ;
        RECT 570.130 735.720 572.510 736.285 ;
        RECT 573.350 735.720 575.730 736.285 ;
        RECT 576.570 735.720 578.950 736.285 ;
        RECT 579.790 735.720 582.170 736.285 ;
        RECT 583.010 735.720 585.390 736.285 ;
        RECT 586.230 735.720 588.610 736.285 ;
        RECT 589.450 735.720 591.830 736.285 ;
        RECT 592.670 735.720 595.050 736.285 ;
        RECT 595.890 735.720 598.270 736.285 ;
        RECT 599.110 735.720 601.490 736.285 ;
        RECT 602.330 735.720 604.710 736.285 ;
        RECT 605.550 735.720 607.930 736.285 ;
        RECT 608.770 735.720 611.150 736.285 ;
        RECT 611.990 735.720 614.370 736.285 ;
        RECT 615.210 735.720 617.130 736.285 ;
        RECT 617.970 735.720 620.350 736.285 ;
        RECT 621.190 735.720 623.570 736.285 ;
        RECT 624.410 735.720 626.790 736.285 ;
        RECT 627.630 735.720 630.010 736.285 ;
        RECT 630.850 735.720 633.230 736.285 ;
        RECT 634.070 735.720 636.450 736.285 ;
        RECT 637.290 735.720 639.670 736.285 ;
        RECT 640.510 735.720 642.890 736.285 ;
        RECT 643.730 735.720 646.110 736.285 ;
        RECT 646.950 735.720 649.330 736.285 ;
        RECT 650.170 735.720 652.550 736.285 ;
        RECT 653.390 735.720 655.770 736.285 ;
        RECT 656.610 735.720 658.990 736.285 ;
        RECT 659.830 735.720 662.210 736.285 ;
        RECT 663.050 735.720 665.430 736.285 ;
        RECT 666.270 735.720 668.650 736.285 ;
        RECT 669.490 735.720 671.870 736.285 ;
        RECT 672.710 735.720 675.090 736.285 ;
        RECT 675.930 735.720 678.310 736.285 ;
        RECT 679.150 735.720 681.530 736.285 ;
        RECT 682.370 735.720 684.750 736.285 ;
        RECT 685.590 735.720 687.970 736.285 ;
        RECT 688.810 735.720 691.190 736.285 ;
        RECT 692.030 735.720 694.410 736.285 ;
        RECT 695.250 735.720 697.630 736.285 ;
        RECT 698.470 735.720 700.850 736.285 ;
        RECT 701.690 735.720 704.070 736.285 ;
        RECT 704.910 735.720 707.290 736.285 ;
        RECT 708.130 735.720 710.510 736.285 ;
        RECT 711.350 735.720 713.730 736.285 ;
        RECT 714.570 735.720 716.950 736.285 ;
        RECT 717.790 735.720 720.170 736.285 ;
        RECT 721.010 735.720 723.390 736.285 ;
        RECT 724.230 735.720 726.610 736.285 ;
        RECT 727.450 735.720 729.830 736.285 ;
        RECT 730.670 735.720 733.050 736.285 ;
        RECT 733.890 735.720 736.270 736.285 ;
        RECT 737.110 735.720 739.490 736.285 ;
        RECT 740.330 735.720 742.710 736.285 ;
        RECT 743.550 735.720 745.930 736.285 ;
        RECT 746.770 735.720 749.150 736.285 ;
        RECT 749.990 735.720 752.370 736.285 ;
        RECT 753.210 735.720 755.590 736.285 ;
        RECT 756.430 735.720 758.810 736.285 ;
        RECT 759.650 735.720 762.030 736.285 ;
        RECT 762.870 735.720 765.250 736.285 ;
        RECT 766.090 735.720 768.470 736.285 ;
        RECT 769.310 735.720 771.230 736.285 ;
        RECT 772.070 735.720 774.450 736.285 ;
        RECT 775.290 735.720 777.670 736.285 ;
        RECT 778.510 735.720 780.890 736.285 ;
        RECT 781.730 735.720 784.110 736.285 ;
        RECT 784.950 735.720 787.330 736.285 ;
        RECT 788.170 735.720 790.550 736.285 ;
        RECT 791.390 735.720 793.770 736.285 ;
        RECT 794.610 735.720 796.990 736.285 ;
        RECT 797.830 735.720 800.210 736.285 ;
        RECT 801.050 735.720 803.430 736.285 ;
        RECT 804.270 735.720 806.650 736.285 ;
        RECT 807.490 735.720 809.870 736.285 ;
        RECT 810.710 735.720 813.090 736.285 ;
        RECT 813.930 735.720 816.310 736.285 ;
        RECT 817.150 735.720 819.530 736.285 ;
        RECT 820.370 735.720 822.750 736.285 ;
        RECT 823.590 735.720 825.970 736.285 ;
        RECT 826.810 735.720 829.190 736.285 ;
        RECT 830.030 735.720 832.410 736.285 ;
        RECT 833.250 735.720 835.630 736.285 ;
        RECT 836.470 735.720 838.850 736.285 ;
        RECT 839.690 735.720 842.070 736.285 ;
        RECT 842.910 735.720 845.290 736.285 ;
        RECT 846.130 735.720 848.510 736.285 ;
        RECT 849.350 735.720 851.730 736.285 ;
        RECT 852.570 735.720 854.950 736.285 ;
        RECT 855.790 735.720 858.170 736.285 ;
        RECT 859.010 735.720 861.390 736.285 ;
        RECT 862.230 735.720 864.610 736.285 ;
        RECT 865.450 735.720 867.830 736.285 ;
        RECT 868.670 735.720 871.050 736.285 ;
        RECT 871.890 735.720 874.270 736.285 ;
        RECT 875.110 735.720 877.490 736.285 ;
        RECT 878.330 735.720 880.710 736.285 ;
        RECT 881.550 735.720 883.930 736.285 ;
        RECT 884.770 735.720 887.150 736.285 ;
        RECT 887.990 735.720 890.370 736.285 ;
        RECT 891.210 735.720 893.590 736.285 ;
        RECT 894.430 735.720 896.810 736.285 ;
        RECT 897.650 735.720 900.030 736.285 ;
        RECT 900.870 735.720 903.250 736.285 ;
        RECT 904.090 735.720 906.470 736.285 ;
        RECT 907.310 735.720 909.690 736.285 ;
        RECT 910.530 735.720 912.910 736.285 ;
        RECT 913.750 735.720 916.130 736.285 ;
        RECT 916.970 735.720 919.350 736.285 ;
        RECT 920.190 735.720 922.570 736.285 ;
        RECT 923.410 735.720 925.330 736.285 ;
        RECT 926.170 735.720 928.550 736.285 ;
        RECT 929.390 735.720 931.770 736.285 ;
        RECT 932.610 735.720 934.990 736.285 ;
        RECT 935.830 735.720 938.210 736.285 ;
        RECT 939.050 735.720 941.430 736.285 ;
        RECT 942.270 735.720 944.650 736.285 ;
        RECT 945.490 735.720 947.870 736.285 ;
        RECT 948.710 735.720 951.090 736.285 ;
        RECT 951.930 735.720 954.310 736.285 ;
        RECT 955.150 735.720 957.530 736.285 ;
        RECT 958.370 735.720 960.750 736.285 ;
        RECT 961.590 735.720 963.970 736.285 ;
        RECT 964.810 735.720 967.190 736.285 ;
        RECT 968.030 735.720 970.410 736.285 ;
        RECT 971.250 735.720 973.630 736.285 ;
        RECT 974.470 735.720 976.850 736.285 ;
        RECT 977.690 735.720 980.070 736.285 ;
        RECT 980.910 735.720 983.290 736.285 ;
        RECT 984.130 735.720 986.510 736.285 ;
        RECT 987.350 735.720 989.730 736.285 ;
        RECT 990.570 735.720 992.950 736.285 ;
        RECT 993.790 735.720 996.170 736.285 ;
        RECT 997.010 735.720 999.390 736.285 ;
        RECT 1000.230 735.720 1002.610 736.285 ;
        RECT 1003.450 735.720 1005.830 736.285 ;
        RECT 1006.670 735.720 1009.050 736.285 ;
        RECT 1009.890 735.720 1012.270 736.285 ;
        RECT 1013.110 735.720 1015.490 736.285 ;
        RECT 1016.330 735.720 1018.710 736.285 ;
        RECT 1019.550 735.720 1021.930 736.285 ;
        RECT 1022.770 735.720 1025.150 736.285 ;
        RECT 1025.990 735.720 1028.370 736.285 ;
        RECT 1029.210 735.720 1031.590 736.285 ;
        RECT 1032.430 735.720 1034.810 736.285 ;
        RECT 1035.650 735.720 1038.030 736.285 ;
        RECT 1038.870 735.720 1041.250 736.285 ;
        RECT 1042.090 735.720 1044.470 736.285 ;
        RECT 1045.310 735.720 1047.690 736.285 ;
        RECT 1048.530 735.720 1050.910 736.285 ;
        RECT 1051.750 735.720 1054.130 736.285 ;
        RECT 1054.970 735.720 1057.350 736.285 ;
        RECT 1058.190 735.720 1060.570 736.285 ;
        RECT 1061.410 735.720 1063.790 736.285 ;
        RECT 1064.630 735.720 1067.010 736.285 ;
        RECT 1067.850 735.720 1070.230 736.285 ;
        RECT 1071.070 735.720 1073.450 736.285 ;
        RECT 1074.290 735.720 1076.670 736.285 ;
        RECT 1077.510 735.720 1079.430 736.285 ;
        RECT 1080.270 735.720 1082.650 736.285 ;
        RECT 1083.490 735.720 1085.870 736.285 ;
        RECT 1086.710 735.720 1089.090 736.285 ;
        RECT 1089.930 735.720 1092.310 736.285 ;
        RECT 1093.150 735.720 1095.530 736.285 ;
        RECT 1096.370 735.720 1098.750 736.285 ;
        RECT 1099.590 735.720 1101.970 736.285 ;
        RECT 1102.810 735.720 1105.190 736.285 ;
        RECT 1106.030 735.720 1108.410 736.285 ;
        RECT 1109.250 735.720 1111.630 736.285 ;
        RECT 1112.470 735.720 1114.850 736.285 ;
        RECT 1115.690 735.720 1118.070 736.285 ;
        RECT 1118.910 735.720 1121.290 736.285 ;
        RECT 1122.130 735.720 1124.510 736.285 ;
        RECT 1125.350 735.720 1127.730 736.285 ;
        RECT 1128.570 735.720 1130.950 736.285 ;
        RECT 1131.790 735.720 1134.170 736.285 ;
        RECT 1135.010 735.720 1137.390 736.285 ;
        RECT 1138.230 735.720 1140.610 736.285 ;
        RECT 1141.450 735.720 1143.830 736.285 ;
        RECT 1144.670 735.720 1147.050 736.285 ;
        RECT 1147.890 735.720 1150.270 736.285 ;
        RECT 1151.110 735.720 1153.490 736.285 ;
        RECT 1154.330 735.720 1156.710 736.285 ;
        RECT 1157.550 735.720 1159.930 736.285 ;
        RECT 1160.770 735.720 1163.150 736.285 ;
        RECT 1163.990 735.720 1166.370 736.285 ;
        RECT 1167.210 735.720 1169.590 736.285 ;
        RECT 1170.430 735.720 1172.810 736.285 ;
        RECT 1173.650 735.720 1176.030 736.285 ;
        RECT 1176.870 735.720 1179.250 736.285 ;
        RECT 1180.090 735.720 1182.470 736.285 ;
        RECT 1183.310 735.720 1185.690 736.285 ;
        RECT 1186.530 735.720 1188.910 736.285 ;
        RECT 1189.750 735.720 1192.130 736.285 ;
        RECT 1192.970 735.720 1195.350 736.285 ;
        RECT 1196.190 735.720 1198.570 736.285 ;
        RECT 1199.410 735.720 1201.790 736.285 ;
        RECT 1202.630 735.720 1205.010 736.285 ;
        RECT 1205.850 735.720 1208.230 736.285 ;
        RECT 1209.070 735.720 1211.450 736.285 ;
        RECT 1212.290 735.720 1214.670 736.285 ;
        RECT 1215.510 735.720 1217.890 736.285 ;
        RECT 1218.730 735.720 1221.110 736.285 ;
        RECT 1221.950 735.720 1224.330 736.285 ;
        RECT 1225.170 735.720 1227.550 736.285 ;
        RECT 1228.390 735.720 1230.770 736.285 ;
        RECT 1231.610 735.720 1233.530 736.285 ;
        RECT 1234.370 735.720 1236.750 736.285 ;
        RECT 1237.590 735.720 1239.970 736.285 ;
        RECT 1240.810 735.720 1243.190 736.285 ;
        RECT 1244.030 735.720 1246.410 736.285 ;
        RECT 1247.250 735.720 1249.630 736.285 ;
        RECT 1250.470 735.720 1252.850 736.285 ;
        RECT 1253.690 735.720 1256.070 736.285 ;
        RECT 1256.910 735.720 1259.290 736.285 ;
        RECT 1260.130 735.720 1262.510 736.285 ;
        RECT 1263.350 735.720 1265.730 736.285 ;
        RECT 1266.570 735.720 1268.950 736.285 ;
        RECT 1269.790 735.720 1272.170 736.285 ;
        RECT 1273.010 735.720 1275.390 736.285 ;
        RECT 1276.230 735.720 1278.610 736.285 ;
        RECT 1279.450 735.720 1281.830 736.285 ;
        RECT 1282.670 735.720 1285.050 736.285 ;
        RECT 1285.890 735.720 1288.270 736.285 ;
        RECT 1289.110 735.720 1291.490 736.285 ;
        RECT 1292.330 735.720 1294.710 736.285 ;
        RECT 1295.550 735.720 1297.930 736.285 ;
        RECT 1298.770 735.720 1301.150 736.285 ;
        RECT 1301.990 735.720 1304.370 736.285 ;
        RECT 1305.210 735.720 1307.590 736.285 ;
        RECT 1308.430 735.720 1310.810 736.285 ;
        RECT 1311.650 735.720 1314.030 736.285 ;
        RECT 1314.870 735.720 1317.250 736.285 ;
        RECT 1318.090 735.720 1320.470 736.285 ;
        RECT 1321.310 735.720 1323.690 736.285 ;
        RECT 1324.530 735.720 1326.910 736.285 ;
        RECT 1327.750 735.720 1330.130 736.285 ;
        RECT 1330.970 735.720 1333.350 736.285 ;
        RECT 1334.190 735.720 1336.570 736.285 ;
        RECT 1337.410 735.720 1339.790 736.285 ;
        RECT 1340.630 735.720 1343.010 736.285 ;
        RECT 1343.850 735.720 1346.230 736.285 ;
        RECT 1347.070 735.720 1349.450 736.285 ;
        RECT 1350.290 735.720 1352.670 736.285 ;
        RECT 1353.510 735.720 1355.890 736.285 ;
        RECT 1356.730 735.720 1359.110 736.285 ;
        RECT 1359.950 735.720 1362.330 736.285 ;
        RECT 1363.170 735.720 1365.550 736.285 ;
        RECT 1366.390 735.720 1368.770 736.285 ;
        RECT 1369.610 735.720 1371.990 736.285 ;
        RECT 1372.830 735.720 1375.210 736.285 ;
        RECT 1376.050 735.720 1378.430 736.285 ;
        RECT 1379.270 735.720 1381.650 736.285 ;
        RECT 1382.490 735.720 1384.870 736.285 ;
        RECT 1385.710 735.720 1387.630 736.285 ;
        RECT 1388.470 735.720 1390.850 736.285 ;
        RECT 1391.690 735.720 1394.070 736.285 ;
        RECT 1394.910 735.720 1397.290 736.285 ;
        RECT 1398.130 735.720 1400.510 736.285 ;
        RECT 1401.350 735.720 1403.730 736.285 ;
        RECT 1404.570 735.720 1406.950 736.285 ;
        RECT 1407.790 735.720 1410.170 736.285 ;
        RECT 1411.010 735.720 1413.390 736.285 ;
        RECT 1414.230 735.720 1416.610 736.285 ;
        RECT 1417.450 735.720 1419.830 736.285 ;
        RECT 1420.670 735.720 1423.050 736.285 ;
        RECT 1423.890 735.720 1426.270 736.285 ;
        RECT 1427.110 735.720 1429.490 736.285 ;
        RECT 1430.330 735.720 1432.710 736.285 ;
        RECT 1433.550 735.720 1435.930 736.285 ;
        RECT 1436.770 735.720 1439.150 736.285 ;
        RECT 1439.990 735.720 1442.370 736.285 ;
        RECT 1443.210 735.720 1445.590 736.285 ;
        RECT 1446.430 735.720 1448.810 736.285 ;
        RECT 1449.650 735.720 1452.030 736.285 ;
        RECT 1452.870 735.720 1455.250 736.285 ;
        RECT 1456.090 735.720 1458.470 736.285 ;
        RECT 1459.310 735.720 1461.690 736.285 ;
        RECT 1462.530 735.720 1464.910 736.285 ;
        RECT 1465.750 735.720 1468.130 736.285 ;
        RECT 1468.970 735.720 1471.350 736.285 ;
        RECT 1472.190 735.720 1474.570 736.285 ;
        RECT 1475.410 735.720 1477.790 736.285 ;
        RECT 1478.630 735.720 1481.010 736.285 ;
        RECT 1481.850 735.720 1484.230 736.285 ;
        RECT 1485.070 735.720 1487.450 736.285 ;
        RECT 1488.290 735.720 1490.670 736.285 ;
        RECT 1491.510 735.720 1493.890 736.285 ;
        RECT 1494.730 735.720 1497.110 736.285 ;
        RECT 1497.950 735.720 1500.330 736.285 ;
        RECT 1501.170 735.720 1503.550 736.285 ;
        RECT 1504.390 735.720 1506.770 736.285 ;
        RECT 1507.610 735.720 1509.990 736.285 ;
        RECT 1510.830 735.720 1513.210 736.285 ;
        RECT 1514.050 735.720 1516.430 736.285 ;
        RECT 1517.270 735.720 1519.650 736.285 ;
        RECT 1520.490 735.720 1522.870 736.285 ;
        RECT 1523.710 735.720 1526.090 736.285 ;
        RECT 1526.930 735.720 1529.310 736.285 ;
        RECT 1530.150 735.720 1532.530 736.285 ;
        RECT 1533.370 735.720 1535.750 736.285 ;
        RECT 1536.590 735.720 1538.970 736.285 ;
        RECT 1539.810 735.720 1541.730 736.285 ;
        RECT 1542.570 735.720 1544.950 736.285 ;
        RECT 1545.790 735.720 1548.170 736.285 ;
        RECT 1549.010 735.720 1551.390 736.285 ;
        RECT 1552.230 735.720 1554.610 736.285 ;
        RECT 1555.450 735.720 1557.830 736.285 ;
        RECT 1558.670 735.720 1561.050 736.285 ;
        RECT 1561.890 735.720 1564.270 736.285 ;
        RECT 1565.110 735.720 1567.490 736.285 ;
        RECT 1568.330 735.720 1570.710 736.285 ;
        RECT 1571.550 735.720 1573.930 736.285 ;
        RECT 1574.770 735.720 1577.150 736.285 ;
        RECT 1577.990 735.720 1580.370 736.285 ;
        RECT 1581.210 735.720 1583.590 736.285 ;
        RECT 1584.430 735.720 1586.810 736.285 ;
        RECT 1587.650 735.720 1590.030 736.285 ;
        RECT 1590.870 735.720 1593.250 736.285 ;
        RECT 1594.090 735.720 1596.470 736.285 ;
        RECT 1597.310 735.720 1599.690 736.285 ;
        RECT 1600.530 735.720 1602.910 736.285 ;
        RECT 1603.750 735.720 1606.130 736.285 ;
        RECT 1606.970 735.720 1609.350 736.285 ;
        RECT 1610.190 735.720 1612.570 736.285 ;
        RECT 1613.410 735.720 1615.790 736.285 ;
        RECT 1616.630 735.720 1619.010 736.285 ;
        RECT 1619.850 735.720 1622.230 736.285 ;
        RECT 1623.070 735.720 1625.450 736.285 ;
        RECT 1626.290 735.720 1628.670 736.285 ;
        RECT 1629.510 735.720 1631.890 736.285 ;
        RECT 1632.730 735.720 1635.110 736.285 ;
        RECT 1635.950 735.720 1638.330 736.285 ;
        RECT 1639.170 735.720 1641.550 736.285 ;
        RECT 1642.390 735.720 1644.770 736.285 ;
        RECT 1645.610 735.720 1647.990 736.285 ;
        RECT 1648.830 735.720 1651.210 736.285 ;
        RECT 1652.050 735.720 1654.430 736.285 ;
        RECT 1655.270 735.720 1657.650 736.285 ;
        RECT 1658.490 735.720 1660.870 736.285 ;
        RECT 1661.710 735.720 1664.090 736.285 ;
        RECT 1664.930 735.720 1667.310 736.285 ;
        RECT 1668.150 735.720 1670.530 736.285 ;
        RECT 1671.370 735.720 1673.750 736.285 ;
        RECT 1674.590 735.720 1676.970 736.285 ;
        RECT 1677.810 735.720 1680.190 736.285 ;
        RECT 1681.030 735.720 1683.410 736.285 ;
        RECT 1684.250 735.720 1686.630 736.285 ;
        RECT 1687.470 735.720 1689.850 736.285 ;
        RECT 1690.690 735.720 1693.070 736.285 ;
        RECT 1693.910 735.720 1695.830 736.285 ;
        RECT 1696.670 735.720 1699.050 736.285 ;
        RECT 1699.890 735.720 1702.270 736.285 ;
        RECT 1703.110 735.720 1705.490 736.285 ;
        RECT 1706.330 735.720 1708.710 736.285 ;
        RECT 1709.550 735.720 1711.930 736.285 ;
        RECT 1712.770 735.720 1715.150 736.285 ;
        RECT 1715.990 735.720 1718.370 736.285 ;
        RECT 1719.210 735.720 1721.590 736.285 ;
        RECT 1722.430 735.720 1724.810 736.285 ;
        RECT 1725.650 735.720 1728.030 736.285 ;
        RECT 1728.870 735.720 1731.250 736.285 ;
        RECT 1732.090 735.720 1734.470 736.285 ;
        RECT 1735.310 735.720 1737.690 736.285 ;
        RECT 1738.530 735.720 1740.910 736.285 ;
        RECT 1741.750 735.720 1744.130 736.285 ;
        RECT 1744.970 735.720 1747.350 736.285 ;
        RECT 1748.190 735.720 1750.570 736.285 ;
        RECT 1751.410 735.720 1753.790 736.285 ;
        RECT 1754.630 735.720 1757.010 736.285 ;
        RECT 1757.850 735.720 1760.230 736.285 ;
        RECT 1761.070 735.720 1763.450 736.285 ;
        RECT 1764.290 735.720 1766.670 736.285 ;
        RECT 1767.510 735.720 1769.890 736.285 ;
        RECT 1770.730 735.720 1773.110 736.285 ;
        RECT 1773.950 735.720 1776.330 736.285 ;
        RECT 1777.170 735.720 1779.550 736.285 ;
        RECT 1780.390 735.720 1782.770 736.285 ;
        RECT 1783.610 735.720 1785.990 736.285 ;
        RECT 1786.830 735.720 1789.210 736.285 ;
        RECT 1790.050 735.720 1792.430 736.285 ;
        RECT 1793.270 735.720 1795.650 736.285 ;
        RECT 1796.490 735.720 1798.870 736.285 ;
        RECT 1799.710 735.720 1802.090 736.285 ;
        RECT 1802.930 735.720 1805.310 736.285 ;
        RECT 1806.150 735.720 1808.530 736.285 ;
        RECT 1809.370 735.720 1811.750 736.285 ;
        RECT 1812.590 735.720 1814.970 736.285 ;
        RECT 1815.810 735.720 1818.190 736.285 ;
        RECT 1819.030 735.720 1821.410 736.285 ;
        RECT 1822.250 735.720 1824.630 736.285 ;
        RECT 1825.470 735.720 1827.850 736.285 ;
        RECT 1828.690 735.720 1831.070 736.285 ;
        RECT 1831.910 735.720 1834.290 736.285 ;
        RECT 1835.130 735.720 1837.510 736.285 ;
        RECT 1838.350 735.720 1840.730 736.285 ;
        RECT 1841.570 735.720 1843.950 736.285 ;
        RECT 1844.790 735.720 1847.170 736.285 ;
        RECT 1848.010 735.720 1849.930 736.285 ;
        RECT 1850.770 735.720 1853.150 736.285 ;
        RECT 1853.990 735.720 1856.370 736.285 ;
        RECT 1857.210 735.720 1859.590 736.285 ;
        RECT 1860.430 735.720 1862.810 736.285 ;
        RECT 1863.650 735.720 1866.030 736.285 ;
        RECT 1866.870 735.720 1869.250 736.285 ;
        RECT 1870.090 735.720 1872.470 736.285 ;
        RECT 1873.310 735.720 1875.690 736.285 ;
        RECT 1876.530 735.720 1878.910 736.285 ;
        RECT 1879.750 735.720 1882.130 736.285 ;
        RECT 1882.970 735.720 1885.350 736.285 ;
        RECT 1886.190 735.720 1888.570 736.285 ;
        RECT 1889.410 735.720 1891.790 736.285 ;
        RECT 1892.630 735.720 1895.010 736.285 ;
        RECT 1895.850 735.720 1898.230 736.285 ;
        RECT 1899.070 735.720 1901.450 736.285 ;
        RECT 1902.290 735.720 1904.670 736.285 ;
        RECT 1905.510 735.720 1907.890 736.285 ;
        RECT 1908.730 735.720 1911.110 736.285 ;
        RECT 1911.950 735.720 1914.330 736.285 ;
        RECT 1915.170 735.720 1917.550 736.285 ;
        RECT 1918.390 735.720 1920.770 736.285 ;
        RECT 1921.610 735.720 1923.990 736.285 ;
        RECT 1924.830 735.720 1927.210 736.285 ;
        RECT 1928.050 735.720 1930.430 736.285 ;
        RECT 1931.270 735.720 1933.650 736.285 ;
        RECT 1934.490 735.720 1936.870 736.285 ;
        RECT 1937.710 735.720 1940.090 736.285 ;
        RECT 1940.930 735.720 1943.310 736.285 ;
        RECT 1944.150 735.720 1946.530 736.285 ;
        RECT 1947.370 735.720 1949.750 736.285 ;
        RECT 1950.590 735.720 1952.970 736.285 ;
        RECT 1953.810 735.720 1956.190 736.285 ;
        RECT 1957.030 735.720 1959.410 736.285 ;
        RECT 1960.250 735.720 1962.630 736.285 ;
        RECT 1963.470 735.720 1965.850 736.285 ;
        RECT 1966.690 735.720 1969.070 736.285 ;
        RECT 1969.910 735.720 1972.290 736.285 ;
        RECT 1973.130 735.720 1975.510 736.285 ;
        RECT 1976.350 735.720 1978.730 736.285 ;
        RECT 1979.570 735.720 1981.950 736.285 ;
        RECT 1982.790 735.720 1985.170 736.285 ;
        RECT 1986.010 735.720 1988.390 736.285 ;
        RECT 1989.230 735.720 1991.610 736.285 ;
        RECT 1992.450 735.720 1994.830 736.285 ;
        RECT 1995.670 735.720 1998.050 736.285 ;
        RECT 1.480 4.280 1998.600 735.720 ;
        RECT 1.480 2.875 124.470 4.280 ;
        RECT 125.310 2.875 374.250 4.280 ;
        RECT 375.090 2.875 624.490 4.280 ;
        RECT 625.330 2.875 874.270 4.280 ;
        RECT 875.110 2.875 1124.510 4.280 ;
        RECT 1125.350 2.875 1374.290 4.280 ;
        RECT 1375.130 2.875 1624.530 4.280 ;
        RECT 1625.370 2.875 1874.310 4.280 ;
        RECT 1875.150 2.875 1998.600 4.280 ;
      LAYER met3 ;
        RECT 4.000 735.440 1995.600 736.265 ;
        RECT 4.400 735.400 1995.600 735.440 ;
        RECT 4.400 734.040 1996.000 735.400 ;
        RECT 4.000 730.000 1996.000 734.040 ;
        RECT 4.000 728.600 1995.600 730.000 ;
        RECT 4.000 725.920 1996.000 728.600 ;
        RECT 4.400 724.520 1996.000 725.920 ;
        RECT 4.000 723.200 1996.000 724.520 ;
        RECT 4.000 721.800 1995.600 723.200 ;
        RECT 4.000 716.400 1996.000 721.800 ;
        RECT 4.400 715.000 1995.600 716.400 ;
        RECT 4.000 709.600 1996.000 715.000 ;
        RECT 4.000 708.200 1995.600 709.600 ;
        RECT 4.000 706.880 1996.000 708.200 ;
        RECT 4.400 705.480 1996.000 706.880 ;
        RECT 4.000 702.800 1996.000 705.480 ;
        RECT 4.000 701.400 1995.600 702.800 ;
        RECT 4.000 697.360 1996.000 701.400 ;
        RECT 4.400 696.000 1996.000 697.360 ;
        RECT 4.400 695.960 1995.600 696.000 ;
        RECT 4.000 694.600 1995.600 695.960 ;
        RECT 4.000 689.200 1996.000 694.600 ;
        RECT 4.000 687.840 1995.600 689.200 ;
        RECT 4.400 687.800 1995.600 687.840 ;
        RECT 4.400 686.440 1996.000 687.800 ;
        RECT 4.000 682.400 1996.000 686.440 ;
        RECT 4.000 681.000 1995.600 682.400 ;
        RECT 4.000 678.320 1996.000 681.000 ;
        RECT 4.400 676.920 1996.000 678.320 ;
        RECT 4.000 675.600 1996.000 676.920 ;
        RECT 4.000 674.200 1995.600 675.600 ;
        RECT 4.000 668.800 1996.000 674.200 ;
        RECT 4.000 668.120 1995.600 668.800 ;
        RECT 4.400 667.400 1995.600 668.120 ;
        RECT 4.400 666.720 1996.000 667.400 ;
        RECT 4.000 662.000 1996.000 666.720 ;
        RECT 4.000 660.600 1995.600 662.000 ;
        RECT 4.000 658.600 1996.000 660.600 ;
        RECT 4.400 657.200 1996.000 658.600 ;
        RECT 4.000 655.200 1996.000 657.200 ;
        RECT 4.000 653.800 1995.600 655.200 ;
        RECT 4.000 649.080 1996.000 653.800 ;
        RECT 4.400 648.400 1996.000 649.080 ;
        RECT 4.400 647.680 1995.600 648.400 ;
        RECT 4.000 647.000 1995.600 647.680 ;
        RECT 4.000 641.600 1996.000 647.000 ;
        RECT 4.000 640.200 1995.600 641.600 ;
        RECT 4.000 639.560 1996.000 640.200 ;
        RECT 4.400 638.160 1996.000 639.560 ;
        RECT 4.000 634.800 1996.000 638.160 ;
        RECT 4.000 633.400 1995.600 634.800 ;
        RECT 4.000 630.040 1996.000 633.400 ;
        RECT 4.400 628.640 1996.000 630.040 ;
        RECT 4.000 628.000 1996.000 628.640 ;
        RECT 4.000 626.600 1995.600 628.000 ;
        RECT 4.000 621.200 1996.000 626.600 ;
        RECT 4.000 620.520 1995.600 621.200 ;
        RECT 4.400 619.800 1995.600 620.520 ;
        RECT 4.400 619.120 1996.000 619.800 ;
        RECT 4.000 614.400 1996.000 619.120 ;
        RECT 4.000 613.000 1995.600 614.400 ;
        RECT 4.000 611.000 1996.000 613.000 ;
        RECT 4.400 609.600 1996.000 611.000 ;
        RECT 4.000 607.600 1996.000 609.600 ;
        RECT 4.000 606.200 1995.600 607.600 ;
        RECT 4.000 601.480 1996.000 606.200 ;
        RECT 4.400 600.800 1996.000 601.480 ;
        RECT 4.400 600.080 1995.600 600.800 ;
        RECT 4.000 599.400 1995.600 600.080 ;
        RECT 4.000 594.000 1996.000 599.400 ;
        RECT 4.000 592.600 1995.600 594.000 ;
        RECT 4.000 591.280 1996.000 592.600 ;
        RECT 4.400 589.880 1996.000 591.280 ;
        RECT 4.000 587.200 1996.000 589.880 ;
        RECT 4.000 585.800 1995.600 587.200 ;
        RECT 4.000 581.760 1996.000 585.800 ;
        RECT 4.400 580.400 1996.000 581.760 ;
        RECT 4.400 580.360 1995.600 580.400 ;
        RECT 4.000 579.000 1995.600 580.360 ;
        RECT 4.000 573.600 1996.000 579.000 ;
        RECT 4.000 572.240 1995.600 573.600 ;
        RECT 4.400 572.200 1995.600 572.240 ;
        RECT 4.400 570.840 1996.000 572.200 ;
        RECT 4.000 566.800 1996.000 570.840 ;
        RECT 4.000 565.400 1995.600 566.800 ;
        RECT 4.000 562.720 1996.000 565.400 ;
        RECT 4.400 561.320 1996.000 562.720 ;
        RECT 4.000 560.000 1996.000 561.320 ;
        RECT 4.000 558.600 1995.600 560.000 ;
        RECT 4.000 553.200 1996.000 558.600 ;
        RECT 4.400 551.800 1995.600 553.200 ;
        RECT 4.000 546.400 1996.000 551.800 ;
        RECT 4.000 545.000 1995.600 546.400 ;
        RECT 4.000 543.680 1996.000 545.000 ;
        RECT 4.400 542.280 1996.000 543.680 ;
        RECT 4.000 539.600 1996.000 542.280 ;
        RECT 4.000 538.200 1995.600 539.600 ;
        RECT 4.000 534.160 1996.000 538.200 ;
        RECT 4.400 532.800 1996.000 534.160 ;
        RECT 4.400 532.760 1995.600 532.800 ;
        RECT 4.000 531.400 1995.600 532.760 ;
        RECT 4.000 526.000 1996.000 531.400 ;
        RECT 4.000 524.640 1995.600 526.000 ;
        RECT 4.400 524.600 1995.600 524.640 ;
        RECT 4.400 523.240 1996.000 524.600 ;
        RECT 4.000 519.200 1996.000 523.240 ;
        RECT 4.000 517.800 1995.600 519.200 ;
        RECT 4.000 514.440 1996.000 517.800 ;
        RECT 4.400 513.040 1996.000 514.440 ;
        RECT 4.000 512.400 1996.000 513.040 ;
        RECT 4.000 511.000 1995.600 512.400 ;
        RECT 4.000 505.600 1996.000 511.000 ;
        RECT 4.000 504.920 1995.600 505.600 ;
        RECT 4.400 504.200 1995.600 504.920 ;
        RECT 4.400 503.520 1996.000 504.200 ;
        RECT 4.000 498.800 1996.000 503.520 ;
        RECT 4.000 497.400 1995.600 498.800 ;
        RECT 4.000 495.400 1996.000 497.400 ;
        RECT 4.400 494.000 1996.000 495.400 ;
        RECT 4.000 492.000 1996.000 494.000 ;
        RECT 4.000 490.600 1995.600 492.000 ;
        RECT 4.000 485.880 1996.000 490.600 ;
        RECT 4.400 485.200 1996.000 485.880 ;
        RECT 4.400 484.480 1995.600 485.200 ;
        RECT 4.000 483.800 1995.600 484.480 ;
        RECT 4.000 478.400 1996.000 483.800 ;
        RECT 4.000 477.000 1995.600 478.400 ;
        RECT 4.000 476.360 1996.000 477.000 ;
        RECT 4.400 474.960 1996.000 476.360 ;
        RECT 4.000 471.600 1996.000 474.960 ;
        RECT 4.000 470.200 1995.600 471.600 ;
        RECT 4.000 466.840 1996.000 470.200 ;
        RECT 4.400 465.440 1996.000 466.840 ;
        RECT 4.000 464.800 1996.000 465.440 ;
        RECT 4.000 463.400 1995.600 464.800 ;
        RECT 4.000 458.000 1996.000 463.400 ;
        RECT 4.000 457.320 1995.600 458.000 ;
        RECT 4.400 456.600 1995.600 457.320 ;
        RECT 4.400 455.920 1996.000 456.600 ;
        RECT 4.000 451.200 1996.000 455.920 ;
        RECT 4.000 449.800 1995.600 451.200 ;
        RECT 4.000 447.120 1996.000 449.800 ;
        RECT 4.400 445.720 1996.000 447.120 ;
        RECT 4.000 444.400 1996.000 445.720 ;
        RECT 4.000 443.000 1995.600 444.400 ;
        RECT 4.000 437.600 1996.000 443.000 ;
        RECT 4.400 436.200 1995.600 437.600 ;
        RECT 4.000 430.800 1996.000 436.200 ;
        RECT 4.000 429.400 1995.600 430.800 ;
        RECT 4.000 428.080 1996.000 429.400 ;
        RECT 4.400 426.680 1996.000 428.080 ;
        RECT 4.000 424.000 1996.000 426.680 ;
        RECT 4.000 422.600 1995.600 424.000 ;
        RECT 4.000 418.560 1996.000 422.600 ;
        RECT 4.400 417.200 1996.000 418.560 ;
        RECT 4.400 417.160 1995.600 417.200 ;
        RECT 4.000 415.800 1995.600 417.160 ;
        RECT 4.000 410.400 1996.000 415.800 ;
        RECT 4.000 409.040 1995.600 410.400 ;
        RECT 4.400 409.000 1995.600 409.040 ;
        RECT 4.400 407.640 1996.000 409.000 ;
        RECT 4.000 403.600 1996.000 407.640 ;
        RECT 4.000 402.200 1995.600 403.600 ;
        RECT 4.000 399.520 1996.000 402.200 ;
        RECT 4.400 398.120 1996.000 399.520 ;
        RECT 4.000 396.800 1996.000 398.120 ;
        RECT 4.000 395.400 1995.600 396.800 ;
        RECT 4.000 390.000 1996.000 395.400 ;
        RECT 4.400 388.600 1995.600 390.000 ;
        RECT 4.000 383.200 1996.000 388.600 ;
        RECT 4.000 381.800 1995.600 383.200 ;
        RECT 4.000 380.480 1996.000 381.800 ;
        RECT 4.400 379.080 1996.000 380.480 ;
        RECT 4.000 376.400 1996.000 379.080 ;
        RECT 4.000 375.000 1995.600 376.400 ;
        RECT 4.000 370.280 1996.000 375.000 ;
        RECT 4.400 368.880 1995.600 370.280 ;
        RECT 4.000 363.480 1996.000 368.880 ;
        RECT 4.000 362.080 1995.600 363.480 ;
        RECT 4.000 360.760 1996.000 362.080 ;
        RECT 4.400 359.360 1996.000 360.760 ;
        RECT 4.000 356.680 1996.000 359.360 ;
        RECT 4.000 355.280 1995.600 356.680 ;
        RECT 4.000 351.240 1996.000 355.280 ;
        RECT 4.400 349.880 1996.000 351.240 ;
        RECT 4.400 349.840 1995.600 349.880 ;
        RECT 4.000 348.480 1995.600 349.840 ;
        RECT 4.000 343.080 1996.000 348.480 ;
        RECT 4.000 341.720 1995.600 343.080 ;
        RECT 4.400 341.680 1995.600 341.720 ;
        RECT 4.400 340.320 1996.000 341.680 ;
        RECT 4.000 336.280 1996.000 340.320 ;
        RECT 4.000 334.880 1995.600 336.280 ;
        RECT 4.000 332.200 1996.000 334.880 ;
        RECT 4.400 330.800 1996.000 332.200 ;
        RECT 4.000 329.480 1996.000 330.800 ;
        RECT 4.000 328.080 1995.600 329.480 ;
        RECT 4.000 322.680 1996.000 328.080 ;
        RECT 4.400 321.280 1995.600 322.680 ;
        RECT 4.000 315.880 1996.000 321.280 ;
        RECT 4.000 314.480 1995.600 315.880 ;
        RECT 4.000 313.160 1996.000 314.480 ;
        RECT 4.400 311.760 1996.000 313.160 ;
        RECT 4.000 309.080 1996.000 311.760 ;
        RECT 4.000 307.680 1995.600 309.080 ;
        RECT 4.000 303.640 1996.000 307.680 ;
        RECT 4.400 302.280 1996.000 303.640 ;
        RECT 4.400 302.240 1995.600 302.280 ;
        RECT 4.000 300.880 1995.600 302.240 ;
        RECT 4.000 295.480 1996.000 300.880 ;
        RECT 4.000 294.080 1995.600 295.480 ;
        RECT 4.000 293.440 1996.000 294.080 ;
        RECT 4.400 292.040 1996.000 293.440 ;
        RECT 4.000 288.680 1996.000 292.040 ;
        RECT 4.000 287.280 1995.600 288.680 ;
        RECT 4.000 283.920 1996.000 287.280 ;
        RECT 4.400 282.520 1996.000 283.920 ;
        RECT 4.000 281.880 1996.000 282.520 ;
        RECT 4.000 280.480 1995.600 281.880 ;
        RECT 4.000 275.080 1996.000 280.480 ;
        RECT 4.000 274.400 1995.600 275.080 ;
        RECT 4.400 273.680 1995.600 274.400 ;
        RECT 4.400 273.000 1996.000 273.680 ;
        RECT 4.000 268.280 1996.000 273.000 ;
        RECT 4.000 266.880 1995.600 268.280 ;
        RECT 4.000 264.880 1996.000 266.880 ;
        RECT 4.400 263.480 1996.000 264.880 ;
        RECT 4.000 261.480 1996.000 263.480 ;
        RECT 4.000 260.080 1995.600 261.480 ;
        RECT 4.000 255.360 1996.000 260.080 ;
        RECT 4.400 254.680 1996.000 255.360 ;
        RECT 4.400 253.960 1995.600 254.680 ;
        RECT 4.000 253.280 1995.600 253.960 ;
        RECT 4.000 247.880 1996.000 253.280 ;
        RECT 4.000 246.480 1995.600 247.880 ;
        RECT 4.000 245.840 1996.000 246.480 ;
        RECT 4.400 244.440 1996.000 245.840 ;
        RECT 4.000 241.080 1996.000 244.440 ;
        RECT 4.000 239.680 1995.600 241.080 ;
        RECT 4.000 236.320 1996.000 239.680 ;
        RECT 4.400 234.920 1996.000 236.320 ;
        RECT 4.000 234.280 1996.000 234.920 ;
        RECT 4.000 232.880 1995.600 234.280 ;
        RECT 4.000 227.480 1996.000 232.880 ;
        RECT 4.000 226.120 1995.600 227.480 ;
        RECT 4.400 226.080 1995.600 226.120 ;
        RECT 4.400 224.720 1996.000 226.080 ;
        RECT 4.000 220.680 1996.000 224.720 ;
        RECT 4.000 219.280 1995.600 220.680 ;
        RECT 4.000 216.600 1996.000 219.280 ;
        RECT 4.400 215.200 1996.000 216.600 ;
        RECT 4.000 213.880 1996.000 215.200 ;
        RECT 4.000 212.480 1995.600 213.880 ;
        RECT 4.000 207.080 1996.000 212.480 ;
        RECT 4.400 205.680 1995.600 207.080 ;
        RECT 4.000 200.280 1996.000 205.680 ;
        RECT 4.000 198.880 1995.600 200.280 ;
        RECT 4.000 197.560 1996.000 198.880 ;
        RECT 4.400 196.160 1996.000 197.560 ;
        RECT 4.000 193.480 1996.000 196.160 ;
        RECT 4.000 192.080 1995.600 193.480 ;
        RECT 4.000 188.040 1996.000 192.080 ;
        RECT 4.400 186.680 1996.000 188.040 ;
        RECT 4.400 186.640 1995.600 186.680 ;
        RECT 4.000 185.280 1995.600 186.640 ;
        RECT 4.000 179.880 1996.000 185.280 ;
        RECT 4.000 178.520 1995.600 179.880 ;
        RECT 4.400 178.480 1995.600 178.520 ;
        RECT 4.400 177.120 1996.000 178.480 ;
        RECT 4.000 173.080 1996.000 177.120 ;
        RECT 4.000 171.680 1995.600 173.080 ;
        RECT 4.000 169.000 1996.000 171.680 ;
        RECT 4.400 167.600 1996.000 169.000 ;
        RECT 4.000 166.280 1996.000 167.600 ;
        RECT 4.000 164.880 1995.600 166.280 ;
        RECT 4.000 159.480 1996.000 164.880 ;
        RECT 4.400 158.080 1995.600 159.480 ;
        RECT 4.000 152.680 1996.000 158.080 ;
        RECT 4.000 151.280 1995.600 152.680 ;
        RECT 4.000 149.280 1996.000 151.280 ;
        RECT 4.400 147.880 1996.000 149.280 ;
        RECT 4.000 145.880 1996.000 147.880 ;
        RECT 4.000 144.480 1995.600 145.880 ;
        RECT 4.000 139.760 1996.000 144.480 ;
        RECT 4.400 139.080 1996.000 139.760 ;
        RECT 4.400 138.360 1995.600 139.080 ;
        RECT 4.000 137.680 1995.600 138.360 ;
        RECT 4.000 132.280 1996.000 137.680 ;
        RECT 4.000 130.880 1995.600 132.280 ;
        RECT 4.000 130.240 1996.000 130.880 ;
        RECT 4.400 128.840 1996.000 130.240 ;
        RECT 4.000 125.480 1996.000 128.840 ;
        RECT 4.000 124.080 1995.600 125.480 ;
        RECT 4.000 120.720 1996.000 124.080 ;
        RECT 4.400 119.320 1996.000 120.720 ;
        RECT 4.000 118.680 1996.000 119.320 ;
        RECT 4.000 117.280 1995.600 118.680 ;
        RECT 4.000 111.880 1996.000 117.280 ;
        RECT 4.000 111.200 1995.600 111.880 ;
        RECT 4.400 110.480 1995.600 111.200 ;
        RECT 4.400 109.800 1996.000 110.480 ;
        RECT 4.000 105.080 1996.000 109.800 ;
        RECT 4.000 103.680 1995.600 105.080 ;
        RECT 4.000 101.680 1996.000 103.680 ;
        RECT 4.400 100.280 1996.000 101.680 ;
        RECT 4.000 98.280 1996.000 100.280 ;
        RECT 4.000 96.880 1995.600 98.280 ;
        RECT 4.000 92.160 1996.000 96.880 ;
        RECT 4.400 91.480 1996.000 92.160 ;
        RECT 4.400 90.760 1995.600 91.480 ;
        RECT 4.000 90.080 1995.600 90.760 ;
        RECT 4.000 84.680 1996.000 90.080 ;
        RECT 4.000 83.280 1995.600 84.680 ;
        RECT 4.000 82.640 1996.000 83.280 ;
        RECT 4.400 81.240 1996.000 82.640 ;
        RECT 4.000 77.880 1996.000 81.240 ;
        RECT 4.000 76.480 1995.600 77.880 ;
        RECT 4.000 72.440 1996.000 76.480 ;
        RECT 4.400 71.080 1996.000 72.440 ;
        RECT 4.400 71.040 1995.600 71.080 ;
        RECT 4.000 69.680 1995.600 71.040 ;
        RECT 4.000 64.280 1996.000 69.680 ;
        RECT 4.000 62.920 1995.600 64.280 ;
        RECT 4.400 62.880 1995.600 62.920 ;
        RECT 4.400 61.520 1996.000 62.880 ;
        RECT 4.000 57.480 1996.000 61.520 ;
        RECT 4.000 56.080 1995.600 57.480 ;
        RECT 4.000 53.400 1996.000 56.080 ;
        RECT 4.400 52.000 1996.000 53.400 ;
        RECT 4.000 50.680 1996.000 52.000 ;
        RECT 4.000 49.280 1995.600 50.680 ;
        RECT 4.000 43.880 1996.000 49.280 ;
        RECT 4.400 42.480 1995.600 43.880 ;
        RECT 4.000 37.080 1996.000 42.480 ;
        RECT 4.000 35.680 1995.600 37.080 ;
        RECT 4.000 34.360 1996.000 35.680 ;
        RECT 4.400 32.960 1996.000 34.360 ;
        RECT 4.000 30.280 1996.000 32.960 ;
        RECT 4.000 28.880 1995.600 30.280 ;
        RECT 4.000 24.840 1996.000 28.880 ;
        RECT 4.400 23.480 1996.000 24.840 ;
        RECT 4.400 23.440 1995.600 23.480 ;
        RECT 4.000 22.080 1995.600 23.440 ;
        RECT 4.000 16.680 1996.000 22.080 ;
        RECT 4.000 15.320 1995.600 16.680 ;
        RECT 4.400 15.280 1995.600 15.320 ;
        RECT 4.400 13.920 1996.000 15.280 ;
        RECT 4.000 9.880 1996.000 13.920 ;
        RECT 4.000 8.480 1995.600 9.880 ;
        RECT 4.000 5.800 1996.000 8.480 ;
        RECT 4.400 4.400 1996.000 5.800 ;
        RECT 4.000 3.760 1996.000 4.400 ;
        RECT 4.000 2.895 1995.600 3.760 ;
      LAYER met4 ;
        RECT 13.670 70.895 25.240 726.065 ;
        RECT 27.640 70.895 50.240 726.065 ;
        RECT 52.640 70.895 75.240 726.065 ;
        RECT 77.640 536.900 100.240 726.065 ;
        RECT 102.640 536.900 125.240 726.065 ;
        RECT 127.640 536.900 150.240 726.065 ;
        RECT 152.640 536.900 175.240 726.065 ;
        RECT 177.640 536.900 200.240 726.065 ;
        RECT 202.640 536.900 225.240 726.065 ;
        RECT 227.640 536.900 250.240 726.065 ;
        RECT 252.640 536.900 275.240 726.065 ;
        RECT 277.640 536.900 300.240 726.065 ;
        RECT 302.640 536.900 325.240 726.065 ;
        RECT 327.640 536.900 350.240 726.065 ;
        RECT 352.640 536.900 375.240 726.065 ;
        RECT 377.640 536.900 400.240 726.065 ;
        RECT 402.640 536.900 425.240 726.065 ;
        RECT 427.640 536.900 450.240 726.065 ;
        RECT 452.640 536.900 475.240 726.065 ;
        RECT 477.640 536.900 500.240 726.065 ;
        RECT 502.640 536.900 525.240 726.065 ;
        RECT 527.640 536.900 550.240 726.065 ;
        RECT 552.640 536.900 575.240 726.065 ;
        RECT 577.640 536.900 600.240 726.065 ;
        RECT 602.640 536.900 625.240 726.065 ;
        RECT 627.640 536.900 650.240 726.065 ;
        RECT 652.640 536.900 675.240 726.065 ;
        RECT 677.640 536.900 700.240 726.065 ;
        RECT 702.640 536.900 725.240 726.065 ;
        RECT 727.640 536.900 750.240 726.065 ;
        RECT 752.640 536.900 775.240 726.065 ;
        RECT 777.640 536.900 800.240 726.065 ;
        RECT 77.640 101.640 800.240 536.900 ;
        RECT 77.640 70.895 100.240 101.640 ;
        RECT 102.640 70.895 125.240 101.640 ;
        RECT 127.640 70.895 150.240 101.640 ;
        RECT 152.640 70.895 175.240 101.640 ;
        RECT 177.640 70.895 200.240 101.640 ;
        RECT 202.640 70.895 225.240 101.640 ;
        RECT 227.640 70.895 250.240 101.640 ;
        RECT 252.640 70.895 275.240 101.640 ;
        RECT 277.640 70.895 300.240 101.640 ;
        RECT 302.640 70.895 325.240 101.640 ;
        RECT 327.640 70.895 350.240 101.640 ;
        RECT 352.640 70.895 375.240 101.640 ;
        RECT 377.640 70.895 400.240 101.640 ;
        RECT 402.640 70.895 425.240 101.640 ;
        RECT 427.640 70.895 450.240 101.640 ;
        RECT 452.640 70.895 475.240 101.640 ;
        RECT 477.640 70.895 500.240 101.640 ;
        RECT 502.640 70.895 525.240 101.640 ;
        RECT 527.640 70.895 550.240 101.640 ;
        RECT 552.640 70.895 575.240 101.640 ;
        RECT 577.640 70.895 600.240 101.640 ;
        RECT 602.640 70.895 625.240 101.640 ;
        RECT 627.640 70.895 650.240 101.640 ;
        RECT 652.640 70.895 675.240 101.640 ;
        RECT 677.640 70.895 700.240 101.640 ;
        RECT 702.640 70.895 725.240 101.640 ;
        RECT 727.640 70.895 750.240 101.640 ;
        RECT 752.640 70.895 775.240 101.640 ;
        RECT 777.640 70.895 800.240 101.640 ;
        RECT 802.640 70.895 825.240 726.065 ;
        RECT 827.640 70.895 850.240 726.065 ;
        RECT 852.640 70.895 875.240 726.065 ;
        RECT 877.640 70.895 900.240 726.065 ;
        RECT 902.640 70.895 925.240 726.065 ;
        RECT 927.640 70.895 950.240 726.065 ;
        RECT 952.640 70.895 975.240 726.065 ;
        RECT 977.640 70.895 1000.240 726.065 ;
        RECT 1002.640 70.895 1025.240 726.065 ;
        RECT 1027.640 70.895 1050.240 726.065 ;
        RECT 1052.640 70.895 1075.240 726.065 ;
        RECT 1077.640 70.895 1100.240 726.065 ;
        RECT 1102.640 70.895 1125.240 726.065 ;
        RECT 1127.640 70.895 1150.240 726.065 ;
        RECT 1152.640 70.895 1175.240 726.065 ;
        RECT 1177.640 70.895 1200.240 726.065 ;
        RECT 1202.640 70.895 1225.240 726.065 ;
        RECT 1227.640 70.895 1250.240 726.065 ;
        RECT 1252.640 70.895 1275.240 726.065 ;
        RECT 1277.640 70.895 1300.240 726.065 ;
        RECT 1302.640 70.895 1325.240 726.065 ;
        RECT 1327.640 70.895 1350.240 726.065 ;
        RECT 1352.640 70.895 1375.240 726.065 ;
        RECT 1377.640 70.895 1400.240 726.065 ;
        RECT 1402.640 70.895 1425.240 726.065 ;
        RECT 1427.640 70.895 1450.240 726.065 ;
        RECT 1452.640 70.895 1475.240 726.065 ;
        RECT 1477.640 70.895 1500.240 726.065 ;
        RECT 1502.640 70.895 1525.240 726.065 ;
        RECT 1527.640 70.895 1550.240 726.065 ;
        RECT 1552.640 70.895 1575.240 726.065 ;
        RECT 1577.640 70.895 1600.240 726.065 ;
        RECT 1602.640 70.895 1625.240 726.065 ;
        RECT 1627.640 70.895 1650.240 726.065 ;
        RECT 1652.640 70.895 1675.240 726.065 ;
        RECT 1677.640 70.895 1700.240 726.065 ;
        RECT 1702.640 70.895 1725.240 726.065 ;
        RECT 1727.640 70.895 1748.625 726.065 ;
      LAYER met5 ;
        RECT 13.460 679.690 1679.340 682.500 ;
        RECT 13.460 614.690 1679.340 674.890 ;
        RECT 13.460 549.690 1679.340 609.890 ;
        RECT 13.460 484.690 1679.340 544.890 ;
        RECT 13.460 419.690 1679.340 479.890 ;
        RECT 13.460 354.690 1679.340 414.890 ;
        RECT 13.460 289.690 1679.340 349.890 ;
        RECT 13.460 235.500 1679.340 284.890 ;
  END
END mgmt_core
END LIBRARY

