VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO RAM128
  CLASS BLOCK ;
  FOREIGN RAM128 ;
  ORIGIN 0.000 0.000 ;
  SIZE 480.000 BY 450.000 ;
  PIN A0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 15.000 480.000 15.600 ;
    END
  END A0[0]
  PIN A0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 24.520 480.000 25.120 ;
    END
  END A0[1]
  PIN A0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 34.040 480.000 34.640 ;
    END
  END A0[2]
  PIN A0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 43.560 480.000 44.160 ;
    END
  END A0[3]
  PIN A0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 53.080 480.000 53.680 ;
    END
  END A0[4]
  PIN A0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 62.600 480.000 63.200 ;
    END
  END A0[5]
  PIN A0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 72.120 480.000 72.720 ;
    END
  END A0[6]
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 281.560 480.000 282.160 ;
    END
  END CLK
  PIN Di0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 129.240 480.000 129.840 ;
    END
  END Di0[0]
  PIN Di0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 224.440 480.000 225.040 ;
    END
  END Di0[10]
  PIN Di0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 233.960 480.000 234.560 ;
    END
  END Di0[11]
  PIN Di0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 243.480 480.000 244.080 ;
    END
  END Di0[12]
  PIN Di0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 253.000 480.000 253.600 ;
    END
  END Di0[13]
  PIN Di0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 262.520 480.000 263.120 ;
    END
  END Di0[14]
  PIN Di0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 272.040 480.000 272.640 ;
    END
  END Di0[15]
  PIN Di0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 291.080 480.000 291.680 ;
    END
  END Di0[16]
  PIN Di0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 300.600 480.000 301.200 ;
    END
  END Di0[17]
  PIN Di0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 310.120 480.000 310.720 ;
    END
  END Di0[18]
  PIN Di0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 319.640 480.000 320.240 ;
    END
  END Di0[19]
  PIN Di0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 138.760 480.000 139.360 ;
    END
  END Di0[1]
  PIN Di0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 329.160 480.000 329.760 ;
    END
  END Di0[20]
  PIN Di0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 338.680 480.000 339.280 ;
    END
  END Di0[21]
  PIN Di0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 348.200 480.000 348.800 ;
    END
  END Di0[22]
  PIN Di0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 357.720 480.000 358.320 ;
    END
  END Di0[23]
  PIN Di0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 367.240 480.000 367.840 ;
    END
  END Di0[24]
  PIN Di0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 376.760 480.000 377.360 ;
    END
  END Di0[25]
  PIN Di0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 386.280 480.000 386.880 ;
    END
  END Di0[26]
  PIN Di0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 395.800 480.000 396.400 ;
    END
  END Di0[27]
  PIN Di0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 405.320 480.000 405.920 ;
    END
  END Di0[28]
  PIN Di0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 414.840 480.000 415.440 ;
    END
  END Di0[29]
  PIN Di0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 148.280 480.000 148.880 ;
    END
  END Di0[2]
  PIN Di0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 424.360 480.000 424.960 ;
    END
  END Di0[30]
  PIN Di0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 433.880 480.000 434.480 ;
    END
  END Di0[31]
  PIN Di0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 157.800 480.000 158.400 ;
    END
  END Di0[3]
  PIN Di0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 167.320 480.000 167.920 ;
    END
  END Di0[4]
  PIN Di0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 176.840 480.000 177.440 ;
    END
  END Di0[5]
  PIN Di0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 186.360 480.000 186.960 ;
    END
  END Di0[6]
  PIN Di0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 195.880 480.000 196.480 ;
    END
  END Di0[7]
  PIN Di0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 205.400 480.000 206.000 ;
    END
  END Di0[8]
  PIN Di0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 214.920 480.000 215.520 ;
    END
  END Di0[9]
  PIN Do0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 446.000 11.870 450.000 ;
    END
  END Do0[0]
  PIN Do0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 446.000 159.070 450.000 ;
    END
  END Do0[10]
  PIN Do0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 446.000 173.790 450.000 ;
    END
  END Do0[11]
  PIN Do0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 446.000 188.510 450.000 ;
    END
  END Do0[12]
  PIN Do0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 446.000 203.230 450.000 ;
    END
  END Do0[13]
  PIN Do0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 446.000 217.950 450.000 ;
    END
  END Do0[14]
  PIN Do0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.390 446.000 232.670 450.000 ;
    END
  END Do0[15]
  PIN Do0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.110 446.000 247.390 450.000 ;
    END
  END Do0[16]
  PIN Do0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.830 446.000 262.110 450.000 ;
    END
  END Do0[17]
  PIN Do0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 446.000 276.830 450.000 ;
    END
  END Do0[18]
  PIN Do0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 446.000 291.550 450.000 ;
    END
  END Do0[19]
  PIN Do0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 446.000 26.590 450.000 ;
    END
  END Do0[1]
  PIN Do0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.990 446.000 306.270 450.000 ;
    END
  END Do0[20]
  PIN Do0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.710 446.000 320.990 450.000 ;
    END
  END Do0[21]
  PIN Do0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 446.000 335.710 450.000 ;
    END
  END Do0[22]
  PIN Do0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.150 446.000 350.430 450.000 ;
    END
  END Do0[23]
  PIN Do0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.870 446.000 365.150 450.000 ;
    END
  END Do0[24]
  PIN Do0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 446.000 379.870 450.000 ;
    END
  END Do0[25]
  PIN Do0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 446.000 394.590 450.000 ;
    END
  END Do0[26]
  PIN Do0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 446.000 409.310 450.000 ;
    END
  END Do0[27]
  PIN Do0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 446.000 424.030 450.000 ;
    END
  END Do0[28]
  PIN Do0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.470 446.000 438.750 450.000 ;
    END
  END Do0[29]
  PIN Do0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.030 446.000 41.310 450.000 ;
    END
  END Do0[2]
  PIN Do0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 446.000 453.470 450.000 ;
    END
  END Do0[30]
  PIN Do0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 467.910 446.000 468.190 450.000 ;
    END
  END Do0[31]
  PIN Do0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 446.000 56.030 450.000 ;
    END
  END Do0[3]
  PIN Do0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 446.000 70.750 450.000 ;
    END
  END Do0[4]
  PIN Do0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 446.000 85.470 450.000 ;
    END
  END Do0[5]
  PIN Do0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 446.000 100.190 450.000 ;
    END
  END Do0[6]
  PIN Do0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 446.000 114.910 450.000 ;
    END
  END Do0[7]
  PIN Do0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 446.000 129.630 450.000 ;
    END
  END Do0[8]
  PIN Do0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 446.000 144.350 450.000 ;
    END
  END Do0[9]
  PIN EN0
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 119.720 480.000 120.320 ;
    END
  END EN0
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.920 10.640 98.520 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 250.520 10.640 252.120 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 404.120 10.640 405.720 438.160 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.120 10.640 21.720 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 173.720 10.640 175.320 438.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 327.320 10.640 328.920 438.160 ;
    END
  END VPWR
  PIN WE0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 81.640 480.000 82.240 ;
    END
  END WE0[0]
  PIN WE0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 91.160 480.000 91.760 ;
    END
  END WE0[1]
  PIN WE0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 100.680 480.000 101.280 ;
    END
  END WE0[2]
  PIN WE0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 476.000 110.200 480.000 110.800 ;
    END
  END WE0[3]
  OBS
      LAYER nwell ;
        RECT 4.410 436.505 475.370 438.110 ;
        RECT 4.410 431.065 475.370 433.895 ;
        RECT 4.410 425.675 475.370 428.455 ;
        RECT 4.410 425.625 73.280 425.675 ;
        RECT 4.410 422.965 13.940 423.015 ;
        RECT 4.410 420.235 475.370 422.965 ;
        RECT 4.410 420.185 88.920 420.235 ;
        RECT 4.410 417.525 39.240 417.575 ;
        RECT 4.410 414.795 475.370 417.525 ;
        RECT 4.410 414.745 10.655 414.795 ;
        RECT 4.410 412.085 176.255 412.135 ;
        RECT 4.410 409.355 475.370 412.085 ;
        RECT 4.410 409.305 97.595 409.355 ;
        RECT 4.410 406.645 109.095 406.695 ;
        RECT 4.410 403.915 475.370 406.645 ;
        RECT 4.410 403.865 46.535 403.915 ;
        RECT 4.410 401.205 24.915 401.255 ;
        RECT 4.410 398.475 475.370 401.205 ;
        RECT 4.410 398.425 99.040 398.475 ;
        RECT 4.410 393.035 475.370 395.815 ;
        RECT 4.410 392.985 12.100 393.035 ;
        RECT 4.410 390.325 27.740 390.375 ;
        RECT 4.410 387.595 475.370 390.325 ;
        RECT 4.410 387.545 11.115 387.595 ;
        RECT 4.410 384.885 102.195 384.935 ;
        RECT 4.410 382.155 475.370 384.885 ;
        RECT 4.410 382.105 186.835 382.155 ;
        RECT 4.410 379.445 58.035 379.495 ;
        RECT 4.410 376.715 475.370 379.445 ;
        RECT 4.410 376.665 92.140 376.715 ;
        RECT 4.410 374.005 31.815 374.055 ;
        RECT 4.410 371.275 475.370 374.005 ;
        RECT 4.410 371.225 321.155 371.275 ;
        RECT 4.410 368.565 128.940 368.615 ;
        RECT 4.410 365.835 475.370 368.565 ;
        RECT 4.410 365.785 49.755 365.835 ;
        RECT 4.410 363.125 19.460 363.175 ;
        RECT 4.410 360.395 475.370 363.125 ;
        RECT 4.410 360.345 23.995 360.395 ;
        RECT 4.410 354.955 475.370 357.735 ;
        RECT 4.410 354.905 49.295 354.955 ;
        RECT 4.410 352.245 169.355 352.295 ;
        RECT 4.410 349.515 475.370 352.245 ;
        RECT 4.410 349.465 26.360 349.515 ;
        RECT 4.410 346.805 164.755 346.855 ;
        RECT 4.410 344.075 475.370 346.805 ;
        RECT 4.410 344.025 85.635 344.075 ;
        RECT 4.410 341.365 167.580 341.415 ;
        RECT 4.410 338.635 475.370 341.365 ;
        RECT 4.410 338.585 29.580 338.635 ;
        RECT 4.410 335.925 138.600 335.975 ;
        RECT 4.410 333.195 475.370 335.925 ;
        RECT 4.410 333.145 253.995 333.195 ;
        RECT 4.410 330.485 134.855 330.535 ;
        RECT 4.410 327.755 475.370 330.485 ;
        RECT 4.410 327.705 74.660 327.755 ;
        RECT 4.410 325.045 23.075 325.095 ;
        RECT 4.410 322.315 475.370 325.045 ;
        RECT 4.410 322.265 32.735 322.315 ;
        RECT 4.410 319.605 99.895 319.655 ;
        RECT 4.410 316.875 475.370 319.605 ;
        RECT 4.410 316.825 158.775 316.875 ;
        RECT 4.410 314.165 96.215 314.215 ;
        RECT 4.410 311.435 475.370 314.165 ;
        RECT 4.410 311.385 23.075 311.435 ;
        RECT 4.410 308.725 21.300 308.775 ;
        RECT 4.410 305.995 475.370 308.725 ;
        RECT 4.410 305.945 33.195 305.995 ;
        RECT 4.410 303.285 109.095 303.335 ;
        RECT 4.410 300.555 475.370 303.285 ;
        RECT 4.410 300.505 305.120 300.555 ;
        RECT 4.410 297.845 57.575 297.895 ;
        RECT 4.410 295.115 475.370 297.845 ;
        RECT 4.410 295.065 23.600 295.115 ;
        RECT 4.410 292.405 144.055 292.455 ;
        RECT 4.410 289.675 475.370 292.405 ;
        RECT 4.410 289.625 70.455 289.675 ;
        RECT 4.410 286.965 53.500 287.015 ;
        RECT 4.410 284.235 475.370 286.965 ;
        RECT 4.410 284.185 176.320 284.235 ;
        RECT 4.410 281.525 289.415 281.575 ;
        RECT 4.410 278.795 475.370 281.525 ;
        RECT 4.410 278.745 21.760 278.795 ;
        RECT 4.410 276.085 70.915 276.135 ;
        RECT 4.410 273.355 475.370 276.085 ;
        RECT 4.410 273.305 21.760 273.355 ;
        RECT 4.410 270.645 50.675 270.695 ;
        RECT 4.410 267.915 475.370 270.645 ;
        RECT 4.410 267.865 176.320 267.915 ;
        RECT 4.410 265.205 31.815 265.255 ;
        RECT 4.410 262.475 475.370 265.205 ;
        RECT 4.410 262.425 180.855 262.475 ;
        RECT 4.410 259.765 307.420 259.815 ;
        RECT 4.410 257.035 475.370 259.765 ;
        RECT 4.410 256.985 23.140 257.035 ;
        RECT 4.410 254.325 45.615 254.375 ;
        RECT 4.410 251.595 475.370 254.325 ;
        RECT 4.410 251.545 449.100 251.595 ;
        RECT 4.410 248.885 443.975 248.935 ;
        RECT 4.410 246.155 475.370 248.885 ;
        RECT 4.410 246.105 279.360 246.155 ;
        RECT 4.410 243.445 289.415 243.495 ;
        RECT 4.410 240.715 475.370 243.445 ;
        RECT 4.410 240.665 380.035 240.715 ;
        RECT 4.410 235.275 475.370 238.055 ;
        RECT 4.410 235.225 303.675 235.275 ;
        RECT 4.410 232.565 394.755 232.615 ;
        RECT 4.410 229.835 475.370 232.565 ;
        RECT 4.410 229.785 334.495 229.835 ;
        RECT 4.410 227.125 292.240 227.175 ;
        RECT 4.410 224.395 475.370 227.125 ;
        RECT 4.410 224.345 10.260 224.395 ;
        RECT 4.410 221.685 24.455 221.735 ;
        RECT 4.410 218.955 475.370 221.685 ;
        RECT 4.410 218.905 48.835 218.955 ;
        RECT 4.410 216.245 147.275 216.295 ;
        RECT 4.410 213.515 475.370 216.245 ;
        RECT 4.410 213.465 103.640 213.515 ;
        RECT 4.410 210.805 27.740 210.855 ;
        RECT 4.410 208.075 475.370 210.805 ;
        RECT 4.410 208.025 10.260 208.075 ;
        RECT 4.410 205.365 145.895 205.415 ;
        RECT 4.410 202.635 475.370 205.365 ;
        RECT 4.410 202.585 58.495 202.635 ;
        RECT 4.410 199.925 126.640 199.975 ;
        RECT 4.410 197.145 475.370 199.925 ;
        RECT 4.410 191.705 475.370 194.535 ;
        RECT 4.410 189.045 325.295 189.095 ;
        RECT 4.410 186.315 475.370 189.045 ;
        RECT 4.410 186.265 21.760 186.315 ;
        RECT 4.410 183.605 43.840 183.655 ;
        RECT 4.410 180.875 475.370 183.605 ;
        RECT 4.410 180.825 108.175 180.875 ;
        RECT 4.410 178.165 96.740 178.215 ;
        RECT 4.410 175.435 475.370 178.165 ;
        RECT 4.410 175.385 353.815 175.435 ;
        RECT 4.410 172.725 61.715 172.775 ;
        RECT 4.410 169.995 475.370 172.725 ;
        RECT 4.410 169.945 312.020 169.995 ;
        RECT 4.410 167.285 21.300 167.335 ;
        RECT 4.410 164.555 475.370 167.285 ;
        RECT 4.410 164.505 23.075 164.555 ;
        RECT 4.410 161.845 110.475 161.895 ;
        RECT 4.410 159.115 475.370 161.845 ;
        RECT 4.410 159.065 80.115 159.115 ;
        RECT 4.410 156.405 42.855 156.455 ;
        RECT 4.410 153.675 475.370 156.405 ;
        RECT 4.410 153.625 383.715 153.675 ;
        RECT 4.410 150.965 23.140 151.015 ;
        RECT 4.410 148.235 475.370 150.965 ;
        RECT 4.410 148.185 27.280 148.235 ;
        RECT 4.410 145.525 186.375 145.575 ;
        RECT 4.410 142.795 475.370 145.525 ;
        RECT 4.410 142.745 73.280 142.795 ;
        RECT 4.410 140.085 34.640 140.135 ;
        RECT 4.410 137.355 475.370 140.085 ;
        RECT 4.410 137.305 53.435 137.355 ;
        RECT 4.410 134.645 38.715 134.695 ;
        RECT 4.410 131.915 475.370 134.645 ;
        RECT 4.410 131.865 30.040 131.915 ;
        RECT 4.410 129.205 36.940 129.255 ;
        RECT 4.410 126.475 475.370 129.205 ;
        RECT 4.410 126.425 345.995 126.475 ;
        RECT 4.410 123.765 268.320 123.815 ;
        RECT 4.410 121.035 475.370 123.765 ;
        RECT 4.410 120.985 173.495 121.035 ;
        RECT 4.410 118.325 237.895 118.375 ;
        RECT 4.410 115.595 475.370 118.325 ;
        RECT 4.410 115.545 154.635 115.595 ;
        RECT 4.410 112.885 121.515 112.935 ;
        RECT 4.410 110.155 475.370 112.885 ;
        RECT 4.410 110.105 165.675 110.155 ;
        RECT 4.410 107.445 69.535 107.495 ;
        RECT 4.410 104.715 475.370 107.445 ;
        RECT 4.410 104.665 18.935 104.715 ;
        RECT 4.410 102.005 167.975 102.055 ;
        RECT 4.410 99.275 475.370 102.005 ;
        RECT 4.410 99.225 100.420 99.275 ;
        RECT 4.410 96.565 224.095 96.615 ;
        RECT 4.410 93.835 475.370 96.565 ;
        RECT 4.410 93.785 126.180 93.835 ;
        RECT 4.410 91.125 188.675 91.175 ;
        RECT 4.410 88.395 475.370 91.125 ;
        RECT 4.410 88.345 63.620 88.395 ;
        RECT 4.410 85.685 134.855 85.735 ;
        RECT 4.410 82.955 475.370 85.685 ;
        RECT 4.410 82.905 10.260 82.955 ;
        RECT 4.410 80.245 23.075 80.295 ;
        RECT 4.410 77.515 475.370 80.245 ;
        RECT 4.410 77.465 45.155 77.515 ;
        RECT 4.410 74.805 192.815 74.855 ;
        RECT 4.410 72.075 475.370 74.805 ;
        RECT 4.410 72.025 88.395 72.075 ;
        RECT 4.410 69.365 255.835 69.415 ;
        RECT 4.410 66.635 475.370 69.365 ;
        RECT 4.410 66.585 234.280 66.635 ;
        RECT 4.410 63.925 19.920 63.975 ;
        RECT 4.410 61.195 475.370 63.925 ;
        RECT 4.410 61.145 443.055 61.195 ;
        RECT 4.410 58.485 89.380 58.535 ;
        RECT 4.410 55.755 475.370 58.485 ;
        RECT 4.410 55.705 21.760 55.755 ;
        RECT 4.410 53.045 99.895 53.095 ;
        RECT 4.410 50.315 475.370 53.045 ;
        RECT 4.410 50.265 44.695 50.315 ;
        RECT 4.410 47.605 237.895 47.655 ;
        RECT 4.410 44.875 475.370 47.605 ;
        RECT 4.410 44.825 137.615 44.875 ;
        RECT 4.410 42.165 115.140 42.215 ;
        RECT 4.410 39.385 475.370 42.165 ;
        RECT 4.410 36.725 48.440 36.775 ;
        RECT 4.410 33.995 475.370 36.725 ;
        RECT 4.410 33.945 10.720 33.995 ;
        RECT 4.410 31.285 23.535 31.335 ;
        RECT 4.410 28.555 475.370 31.285 ;
        RECT 4.410 28.505 87.935 28.555 ;
        RECT 4.410 25.845 113.760 25.895 ;
        RECT 4.410 23.115 475.370 25.845 ;
        RECT 4.410 23.065 70.455 23.115 ;
        RECT 4.410 17.625 475.370 20.455 ;
        RECT 4.410 12.185 475.370 15.015 ;
      LAYER li1 ;
        RECT 4.600 10.795 475.180 438.005 ;
      LAYER met1 ;
        RECT 4.600 9.560 475.480 439.920 ;
      LAYER met2 ;
        RECT 6.080 445.720 11.310 446.490 ;
        RECT 12.150 445.720 26.030 446.490 ;
        RECT 26.870 445.720 40.750 446.490 ;
        RECT 41.590 445.720 55.470 446.490 ;
        RECT 56.310 445.720 70.190 446.490 ;
        RECT 71.030 445.720 84.910 446.490 ;
        RECT 85.750 445.720 99.630 446.490 ;
        RECT 100.470 445.720 114.350 446.490 ;
        RECT 115.190 445.720 129.070 446.490 ;
        RECT 129.910 445.720 143.790 446.490 ;
        RECT 144.630 445.720 158.510 446.490 ;
        RECT 159.350 445.720 173.230 446.490 ;
        RECT 174.070 445.720 187.950 446.490 ;
        RECT 188.790 445.720 202.670 446.490 ;
        RECT 203.510 445.720 217.390 446.490 ;
        RECT 218.230 445.720 232.110 446.490 ;
        RECT 232.950 445.720 246.830 446.490 ;
        RECT 247.670 445.720 261.550 446.490 ;
        RECT 262.390 445.720 276.270 446.490 ;
        RECT 277.110 445.720 290.990 446.490 ;
        RECT 291.830 445.720 305.710 446.490 ;
        RECT 306.550 445.720 320.430 446.490 ;
        RECT 321.270 445.720 335.150 446.490 ;
        RECT 335.990 445.720 349.870 446.490 ;
        RECT 350.710 445.720 364.590 446.490 ;
        RECT 365.430 445.720 379.310 446.490 ;
        RECT 380.150 445.720 394.030 446.490 ;
        RECT 394.870 445.720 408.750 446.490 ;
        RECT 409.590 445.720 423.470 446.490 ;
        RECT 424.310 445.720 438.190 446.490 ;
        RECT 439.030 445.720 452.910 446.490 ;
        RECT 453.750 445.720 467.630 446.490 ;
        RECT 468.470 445.720 475.090 446.490 ;
        RECT 6.080 9.530 475.090 445.720 ;
      LAYER met3 ;
        RECT 7.885 434.880 476.000 438.085 ;
        RECT 7.885 433.480 475.600 434.880 ;
        RECT 7.885 425.360 476.000 433.480 ;
        RECT 7.885 423.960 475.600 425.360 ;
        RECT 7.885 415.840 476.000 423.960 ;
        RECT 7.885 414.440 475.600 415.840 ;
        RECT 7.885 406.320 476.000 414.440 ;
        RECT 7.885 404.920 475.600 406.320 ;
        RECT 7.885 396.800 476.000 404.920 ;
        RECT 7.885 395.400 475.600 396.800 ;
        RECT 7.885 387.280 476.000 395.400 ;
        RECT 7.885 385.880 475.600 387.280 ;
        RECT 7.885 377.760 476.000 385.880 ;
        RECT 7.885 376.360 475.600 377.760 ;
        RECT 7.885 368.240 476.000 376.360 ;
        RECT 7.885 366.840 475.600 368.240 ;
        RECT 7.885 358.720 476.000 366.840 ;
        RECT 7.885 357.320 475.600 358.720 ;
        RECT 7.885 349.200 476.000 357.320 ;
        RECT 7.885 347.800 475.600 349.200 ;
        RECT 7.885 339.680 476.000 347.800 ;
        RECT 7.885 338.280 475.600 339.680 ;
        RECT 7.885 330.160 476.000 338.280 ;
        RECT 7.885 328.760 475.600 330.160 ;
        RECT 7.885 320.640 476.000 328.760 ;
        RECT 7.885 319.240 475.600 320.640 ;
        RECT 7.885 311.120 476.000 319.240 ;
        RECT 7.885 309.720 475.600 311.120 ;
        RECT 7.885 301.600 476.000 309.720 ;
        RECT 7.885 300.200 475.600 301.600 ;
        RECT 7.885 292.080 476.000 300.200 ;
        RECT 7.885 290.680 475.600 292.080 ;
        RECT 7.885 282.560 476.000 290.680 ;
        RECT 7.885 281.160 475.600 282.560 ;
        RECT 7.885 273.040 476.000 281.160 ;
        RECT 7.885 271.640 475.600 273.040 ;
        RECT 7.885 263.520 476.000 271.640 ;
        RECT 7.885 262.120 475.600 263.520 ;
        RECT 7.885 254.000 476.000 262.120 ;
        RECT 7.885 252.600 475.600 254.000 ;
        RECT 7.885 244.480 476.000 252.600 ;
        RECT 7.885 243.080 475.600 244.480 ;
        RECT 7.885 234.960 476.000 243.080 ;
        RECT 7.885 233.560 475.600 234.960 ;
        RECT 7.885 225.440 476.000 233.560 ;
        RECT 7.885 224.040 475.600 225.440 ;
        RECT 7.885 215.920 476.000 224.040 ;
        RECT 7.885 214.520 475.600 215.920 ;
        RECT 7.885 206.400 476.000 214.520 ;
        RECT 7.885 205.000 475.600 206.400 ;
        RECT 7.885 196.880 476.000 205.000 ;
        RECT 7.885 195.480 475.600 196.880 ;
        RECT 7.885 187.360 476.000 195.480 ;
        RECT 7.885 185.960 475.600 187.360 ;
        RECT 7.885 177.840 476.000 185.960 ;
        RECT 7.885 176.440 475.600 177.840 ;
        RECT 7.885 168.320 476.000 176.440 ;
        RECT 7.885 166.920 475.600 168.320 ;
        RECT 7.885 158.800 476.000 166.920 ;
        RECT 7.885 157.400 475.600 158.800 ;
        RECT 7.885 149.280 476.000 157.400 ;
        RECT 7.885 147.880 475.600 149.280 ;
        RECT 7.885 139.760 476.000 147.880 ;
        RECT 7.885 138.360 475.600 139.760 ;
        RECT 7.885 130.240 476.000 138.360 ;
        RECT 7.885 128.840 475.600 130.240 ;
        RECT 7.885 120.720 476.000 128.840 ;
        RECT 7.885 119.320 475.600 120.720 ;
        RECT 7.885 111.200 476.000 119.320 ;
        RECT 7.885 109.800 475.600 111.200 ;
        RECT 7.885 101.680 476.000 109.800 ;
        RECT 7.885 100.280 475.600 101.680 ;
        RECT 7.885 92.160 476.000 100.280 ;
        RECT 7.885 90.760 475.600 92.160 ;
        RECT 7.885 82.640 476.000 90.760 ;
        RECT 7.885 81.240 475.600 82.640 ;
        RECT 7.885 73.120 476.000 81.240 ;
        RECT 7.885 71.720 475.600 73.120 ;
        RECT 7.885 63.600 476.000 71.720 ;
        RECT 7.885 62.200 475.600 63.600 ;
        RECT 7.885 54.080 476.000 62.200 ;
        RECT 7.885 52.680 475.600 54.080 ;
        RECT 7.885 44.560 476.000 52.680 ;
        RECT 7.885 43.160 475.600 44.560 ;
        RECT 7.885 35.040 476.000 43.160 ;
        RECT 7.885 33.640 475.600 35.040 ;
        RECT 7.885 25.520 476.000 33.640 ;
        RECT 7.885 24.120 475.600 25.520 ;
        RECT 7.885 16.000 476.000 24.120 ;
        RECT 7.885 14.600 475.600 16.000 ;
        RECT 7.885 10.715 476.000 14.600 ;
      LAYER met4 ;
        RECT 18.695 11.735 19.720 433.665 ;
        RECT 22.120 11.735 96.520 433.665 ;
        RECT 98.920 11.735 173.320 433.665 ;
        RECT 175.720 11.735 250.120 433.665 ;
        RECT 252.520 11.735 326.920 433.665 ;
        RECT 329.320 11.735 403.720 433.665 ;
        RECT 406.120 11.735 467.065 433.665 ;
  END
END RAM128
END LIBRARY

