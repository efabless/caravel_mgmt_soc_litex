VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_core_wrapper
  CLASS BLOCK ;
  FOREIGN mgmt_core_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2620.000 BY 820.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -0.780 2.700 0.820 816.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 2.700 2620.480 4.300 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 814.420 2620.480 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.880 2.700 2620.480 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 37.240 2.700 38.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 87.240 2.700 88.840 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 87.240 658.605 88.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 137.240 2.700 138.840 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 137.240 658.605 138.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 187.240 2.700 188.840 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 187.240 658.605 188.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.240 2.700 238.840 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 237.240 658.605 238.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 287.240 2.700 288.840 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 287.240 658.605 288.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 337.240 2.700 338.840 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 337.240 658.605 338.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.240 2.700 388.840 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 387.240 658.605 388.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 437.240 2.700 438.840 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 437.240 658.605 438.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 487.240 2.700 488.840 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 487.240 658.605 488.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 537.240 2.700 538.840 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 537.240 658.605 538.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 587.240 2.700 588.840 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 587.240 658.605 588.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 637.240 2.700 638.840 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 637.240 658.605 638.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 687.240 2.700 688.840 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 687.240 658.605 688.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 737.240 2.700 738.840 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 737.240 658.605 738.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 787.240 2.700 788.840 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 787.240 658.605 788.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.240 2.700 838.840 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 837.240 660.380 838.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 887.240 2.700 888.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 937.240 2.700 938.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 987.240 2.700 988.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1037.240 2.700 1038.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1087.240 2.700 1088.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1137.240 2.700 1138.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1187.240 2.700 1188.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1237.240 2.700 1238.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1287.240 2.700 1288.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1337.240 2.700 1338.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1387.240 2.700 1388.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1437.240 2.700 1438.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1487.240 2.700 1488.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1537.240 2.700 1538.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1587.240 2.700 1588.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1637.240 2.700 1638.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1687.240 2.700 1688.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.240 2.700 1738.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.240 2.700 1788.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1837.240 2.700 1838.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1887.240 2.700 1888.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1937.240 2.700 1938.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1987.240 2.700 1988.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2037.240 2.700 2038.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2087.240 2.700 2088.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2137.240 2.700 2138.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.240 2.700 2188.840 242.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2187.240 652.220 2188.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2237.240 2.700 2238.840 258.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 2237.240 654.525 2238.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2287.240 2.700 2288.840 258.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 2287.240 654.525 2288.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2337.240 2.700 2338.840 258.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 2337.240 654.525 2338.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2387.240 2.700 2388.840 258.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 2387.240 654.525 2388.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.240 2.700 2438.840 258.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.240 654.525 2438.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2487.240 2.700 2488.840 258.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 2487.240 654.525 2488.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2537.240 2.700 2538.840 258.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 2537.240 654.525 2538.840 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2587.240 2.700 2588.840 816.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 41.050 2620.480 42.650 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 91.050 2620.480 92.650 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 141.050 2620.480 142.650 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 191.050 2620.480 192.650 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 241.050 2620.480 242.650 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 291.050 2620.480 292.650 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 341.050 2620.480 342.650 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 391.050 2620.480 392.650 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 441.050 2620.480 442.650 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 491.050 2620.480 492.650 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 541.050 2620.480 542.650 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 591.050 2620.480 592.650 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 641.050 2620.480 642.650 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 691.050 2620.480 692.650 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 741.050 2620.480 742.650 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 791.050 2620.480 792.650 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2.520 6.000 4.120 812.720 ;
    END
    PORT
      LAYER met5 ;
        RECT 2.520 6.000 2617.180 7.600 ;
    END
    PORT
      LAYER met5 ;
        RECT 2.520 811.120 2617.180 812.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 2615.580 6.000 2617.180 812.720 ;
    END
    PORT
      LAYER met4 ;
        RECT 25.640 2.700 27.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 75.640 2.700 77.240 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 75.640 658.605 77.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.640 2.700 127.240 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.640 658.605 127.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 175.640 2.700 177.240 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 175.640 658.605 177.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 225.640 2.700 227.240 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 225.640 658.605 227.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 275.640 2.700 277.240 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 275.640 658.605 277.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.640 2.700 327.240 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.640 658.605 327.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 375.640 2.700 377.240 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 375.640 660.380 377.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 425.640 2.700 427.240 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 425.640 658.605 427.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 475.640 2.700 477.240 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 475.640 658.605 477.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 525.640 2.700 527.240 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 525.640 658.605 527.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.640 2.700 577.240 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.640 658.605 577.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 625.640 2.700 627.240 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 625.640 658.605 627.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.640 2.700 677.240 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.640 658.605 677.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 725.640 2.700 727.240 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 725.640 658.605 727.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 775.640 2.700 777.240 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 775.640 658.605 777.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 825.640 2.700 827.240 239.875 ;
    END
    PORT
      LAYER met4 ;
        RECT 825.640 658.605 827.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 875.640 2.700 877.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 925.640 2.700 927.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 975.640 2.700 977.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.640 2.700 1027.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1075.640 2.700 1077.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1125.640 2.700 1127.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1175.640 2.700 1177.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1225.640 2.700 1227.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.640 2.700 1277.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1325.640 2.700 1327.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1375.640 2.700 1377.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1425.640 2.700 1427.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.640 2.700 1477.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1525.640 2.700 1527.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1575.640 2.700 1577.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1625.640 2.700 1627.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1675.640 2.700 1677.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1725.640 2.700 1727.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1775.640 2.700 1777.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1825.640 2.700 1827.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1875.640 2.700 1877.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1925.640 2.700 1927.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 1975.640 2.700 1977.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2025.640 2.700 2027.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2075.640 2.700 2077.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2125.640 2.700 2127.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2175.640 2.700 2177.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2225.640 2.700 2227.240 258.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 2225.640 654.525 2227.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2275.640 2.700 2277.240 258.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 2275.640 654.525 2277.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.640 2.700 2327.240 258.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.640 654.525 2327.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2375.640 2.700 2377.240 258.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 2375.640 654.525 2377.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2425.640 2.700 2427.240 258.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 2425.640 654.525 2427.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2475.640 2.700 2477.240 258.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 2475.640 654.525 2477.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2525.640 2.700 2527.240 258.235 ;
    END
    PORT
      LAYER met4 ;
        RECT 2525.640 654.525 2527.240 816.020 ;
    END
    PORT
      LAYER met4 ;
        RECT 2575.640 2.700 2577.240 816.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 29.450 2620.480 31.050 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 79.450 2620.480 81.050 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 129.450 2620.480 131.050 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 179.450 2620.480 181.050 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 229.450 2620.480 231.050 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 279.450 2620.480 281.050 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 329.450 2620.480 331.050 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 379.450 2620.480 381.050 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 429.450 2620.480 431.050 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 479.450 2620.480 481.050 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 529.450 2620.480 531.050 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 579.450 2620.480 581.050 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 629.450 2620.480 631.050 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 679.450 2620.480 681.050 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 729.450 2620.480 731.050 ;
    END
    PORT
      LAYER met5 ;
        RECT -0.780 779.450 2620.480 781.050 ;
    END
    PORT
      LAYER met4 ;
        RECT 2594.980 239.120 2596.580 658.480 ;
    END
  END VPWR
  PIN clk_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1309.860 0.000 1310.140 4.000 ;
    END
  END clk_in
  PIN clk_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1193.790 816.000 1194.070 820.000 ;
    END
  END clk_out
  PIN core_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1299.860 0.000 1300.140 4.000 ;
    END
  END core_clk
  PIN core_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1319.860 0.000 1320.140 4.000 ;
    END
  END core_rstn
  PIN debug_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 88.440 2620.000 89.040 ;
    END
  END debug_in
  PIN debug_mode
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 99.320 2620.000 99.920 ;
    END
  END debug_mode
  PIN debug_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 110.200 2620.000 110.800 ;
    END
  END debug_oeb
  PIN debug_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 121.080 2620.000 121.680 ;
    END
  END debug_out
  PIN flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 675.960 2620.000 676.560 ;
    END
  END flash_clk
  PIN flash_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 665.080 2620.000 665.680 ;
    END
  END flash_csb
  PIN flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 686.840 2620.000 687.440 ;
    END
  END flash_io0_di
  PIN flash_io0_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 697.720 2620.000 698.320 ;
    END
  END flash_io0_do
  PIN flash_io0_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 708.600 2620.000 709.200 ;
    END
  END flash_io0_oeb
  PIN flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 719.480 2620.000 720.080 ;
    END
  END flash_io1_di
  PIN flash_io1_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 730.360 2620.000 730.960 ;
    END
  END flash_io1_do
  PIN flash_io1_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 741.240 2620.000 741.840 ;
    END
  END flash_io1_oeb
  PIN flash_io2_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 752.120 2620.000 752.720 ;
    END
  END flash_io2_di
  PIN flash_io2_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 763.000 2620.000 763.600 ;
    END
  END flash_io2_do
  PIN flash_io2_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 773.880 2620.000 774.480 ;
    END
  END flash_io2_oeb
  PIN flash_io3_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 784.760 2620.000 785.360 ;
    END
  END flash_io3_di
  PIN flash_io3_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 795.640 2620.000 796.240 ;
    END
  END flash_io3_do
  PIN flash_io3_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 806.520 2620.000 807.120 ;
    END
  END flash_io3_oeb
  PIN gpio_in_pad
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2459.860 0.000 2460.140 4.000 ;
    END
  END gpio_in_pad
  PIN gpio_inenb_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2469.860 0.000 2470.140 4.000 ;
    END
  END gpio_inenb_pad
  PIN gpio_mode0_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2479.860 0.000 2480.140 4.000 ;
    END
  END gpio_mode0_pad
  PIN gpio_mode1_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2489.860 0.000 2490.140 4.000 ;
    END
  END gpio_mode1_pad
  PIN gpio_out_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2499.860 0.000 2500.140 4.000 ;
    END
  END gpio_out_pad
  PIN gpio_outenb_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2509.860 0.000 2510.140 4.000 ;
    END
  END gpio_outenb_pad
  PIN hk_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 284.280 2620.000 284.880 ;
    END
  END hk_ack_i
  PIN hk_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 306.040 2620.000 306.640 ;
    END
  END hk_cyc_o
  PIN hk_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 316.920 2620.000 317.520 ;
    END
  END hk_dat_i[0]
  PIN hk_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 425.720 2620.000 426.320 ;
    END
  END hk_dat_i[10]
  PIN hk_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 436.600 2620.000 437.200 ;
    END
  END hk_dat_i[11]
  PIN hk_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 447.480 2620.000 448.080 ;
    END
  END hk_dat_i[12]
  PIN hk_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 458.360 2620.000 458.960 ;
    END
  END hk_dat_i[13]
  PIN hk_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 469.240 2620.000 469.840 ;
    END
  END hk_dat_i[14]
  PIN hk_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 480.120 2620.000 480.720 ;
    END
  END hk_dat_i[15]
  PIN hk_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 491.000 2620.000 491.600 ;
    END
  END hk_dat_i[16]
  PIN hk_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 501.880 2620.000 502.480 ;
    END
  END hk_dat_i[17]
  PIN hk_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 512.760 2620.000 513.360 ;
    END
  END hk_dat_i[18]
  PIN hk_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 523.640 2620.000 524.240 ;
    END
  END hk_dat_i[19]
  PIN hk_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 327.800 2620.000 328.400 ;
    END
  END hk_dat_i[1]
  PIN hk_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 534.520 2620.000 535.120 ;
    END
  END hk_dat_i[20]
  PIN hk_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 545.400 2620.000 546.000 ;
    END
  END hk_dat_i[21]
  PIN hk_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 556.280 2620.000 556.880 ;
    END
  END hk_dat_i[22]
  PIN hk_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 567.160 2620.000 567.760 ;
    END
  END hk_dat_i[23]
  PIN hk_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 578.040 2620.000 578.640 ;
    END
  END hk_dat_i[24]
  PIN hk_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 588.920 2620.000 589.520 ;
    END
  END hk_dat_i[25]
  PIN hk_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 599.800 2620.000 600.400 ;
    END
  END hk_dat_i[26]
  PIN hk_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 610.680 2620.000 611.280 ;
    END
  END hk_dat_i[27]
  PIN hk_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 621.560 2620.000 622.160 ;
    END
  END hk_dat_i[28]
  PIN hk_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 632.440 2620.000 633.040 ;
    END
  END hk_dat_i[29]
  PIN hk_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 338.680 2620.000 339.280 ;
    END
  END hk_dat_i[2]
  PIN hk_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 643.320 2620.000 643.920 ;
    END
  END hk_dat_i[30]
  PIN hk_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 654.200 2620.000 654.800 ;
    END
  END hk_dat_i[31]
  PIN hk_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 349.560 2620.000 350.160 ;
    END
  END hk_dat_i[3]
  PIN hk_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 360.440 2620.000 361.040 ;
    END
  END hk_dat_i[4]
  PIN hk_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 371.320 2620.000 371.920 ;
    END
  END hk_dat_i[5]
  PIN hk_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 382.200 2620.000 382.800 ;
    END
  END hk_dat_i[6]
  PIN hk_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 393.080 2620.000 393.680 ;
    END
  END hk_dat_i[7]
  PIN hk_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 403.960 2620.000 404.560 ;
    END
  END hk_dat_i[8]
  PIN hk_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 414.840 2620.000 415.440 ;
    END
  END hk_dat_i[9]
  PIN hk_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 295.160 2620.000 295.760 ;
    END
  END hk_stb_o
  PIN irq[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2593.110 816.000 2593.390 820.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2597.250 816.000 2597.530 820.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2601.390 816.000 2601.670 820.000 ;
    END
  END irq[2]
  PIN irq[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 164.600 2620.000 165.200 ;
    END
  END irq[3]
  PIN irq[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 153.720 2620.000 154.320 ;
    END
  END irq[4]
  PIN irq[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 142.840 2620.000 143.440 ;
    END
  END irq[5]
  PIN la_iena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 816.000 18.310 820.000 ;
    END
  END la_iena[0]
  PIN la_iena[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1682.310 816.000 1682.590 820.000 ;
    END
  END la_iena[100]
  PIN la_iena[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1698.870 816.000 1699.150 820.000 ;
    END
  END la_iena[101]
  PIN la_iena[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.430 816.000 1715.710 820.000 ;
    END
  END la_iena[102]
  PIN la_iena[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1731.990 816.000 1732.270 820.000 ;
    END
  END la_iena[103]
  PIN la_iena[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1748.550 816.000 1748.830 820.000 ;
    END
  END la_iena[104]
  PIN la_iena[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1765.110 816.000 1765.390 820.000 ;
    END
  END la_iena[105]
  PIN la_iena[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.670 816.000 1781.950 820.000 ;
    END
  END la_iena[106]
  PIN la_iena[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1798.230 816.000 1798.510 820.000 ;
    END
  END la_iena[107]
  PIN la_iena[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1814.790 816.000 1815.070 820.000 ;
    END
  END la_iena[108]
  PIN la_iena[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1831.350 816.000 1831.630 820.000 ;
    END
  END la_iena[109]
  PIN la_iena[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 816.000 183.910 820.000 ;
    END
  END la_iena[10]
  PIN la_iena[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1847.910 816.000 1848.190 820.000 ;
    END
  END la_iena[110]
  PIN la_iena[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.470 816.000 1864.750 820.000 ;
    END
  END la_iena[111]
  PIN la_iena[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.030 816.000 1881.310 820.000 ;
    END
  END la_iena[112]
  PIN la_iena[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1897.590 816.000 1897.870 820.000 ;
    END
  END la_iena[113]
  PIN la_iena[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1914.150 816.000 1914.430 820.000 ;
    END
  END la_iena[114]
  PIN la_iena[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1930.710 816.000 1930.990 820.000 ;
    END
  END la_iena[115]
  PIN la_iena[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.270 816.000 1947.550 820.000 ;
    END
  END la_iena[116]
  PIN la_iena[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1963.830 816.000 1964.110 820.000 ;
    END
  END la_iena[117]
  PIN la_iena[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1980.390 816.000 1980.670 820.000 ;
    END
  END la_iena[118]
  PIN la_iena[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1996.950 816.000 1997.230 820.000 ;
    END
  END la_iena[119]
  PIN la_iena[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.190 816.000 200.470 820.000 ;
    END
  END la_iena[11]
  PIN la_iena[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2013.510 816.000 2013.790 820.000 ;
    END
  END la_iena[120]
  PIN la_iena[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.070 816.000 2030.350 820.000 ;
    END
  END la_iena[121]
  PIN la_iena[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2046.630 816.000 2046.910 820.000 ;
    END
  END la_iena[122]
  PIN la_iena[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2063.190 816.000 2063.470 820.000 ;
    END
  END la_iena[123]
  PIN la_iena[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2079.750 816.000 2080.030 820.000 ;
    END
  END la_iena[124]
  PIN la_iena[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2096.310 816.000 2096.590 820.000 ;
    END
  END la_iena[125]
  PIN la_iena[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.870 816.000 2113.150 820.000 ;
    END
  END la_iena[126]
  PIN la_iena[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2129.430 816.000 2129.710 820.000 ;
    END
  END la_iena[127]
  PIN la_iena[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 816.000 217.030 820.000 ;
    END
  END la_iena[12]
  PIN la_iena[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 816.000 233.590 820.000 ;
    END
  END la_iena[13]
  PIN la_iena[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.870 816.000 250.150 820.000 ;
    END
  END la_iena[14]
  PIN la_iena[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.430 816.000 266.710 820.000 ;
    END
  END la_iena[15]
  PIN la_iena[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.990 816.000 283.270 820.000 ;
    END
  END la_iena[16]
  PIN la_iena[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 816.000 299.830 820.000 ;
    END
  END la_iena[17]
  PIN la_iena[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.110 816.000 316.390 820.000 ;
    END
  END la_iena[18]
  PIN la_iena[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.670 816.000 332.950 820.000 ;
    END
  END la_iena[19]
  PIN la_iena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.590 816.000 34.870 820.000 ;
    END
  END la_iena[1]
  PIN la_iena[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 816.000 349.510 820.000 ;
    END
  END la_iena[20]
  PIN la_iena[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 816.000 366.070 820.000 ;
    END
  END la_iena[21]
  PIN la_iena[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.350 816.000 382.630 820.000 ;
    END
  END la_iena[22]
  PIN la_iena[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.910 816.000 399.190 820.000 ;
    END
  END la_iena[23]
  PIN la_iena[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 816.000 415.750 820.000 ;
    END
  END la_iena[24]
  PIN la_iena[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.030 816.000 432.310 820.000 ;
    END
  END la_iena[25]
  PIN la_iena[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.590 816.000 448.870 820.000 ;
    END
  END la_iena[26]
  PIN la_iena[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.150 816.000 465.430 820.000 ;
    END
  END la_iena[27]
  PIN la_iena[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.710 816.000 481.990 820.000 ;
    END
  END la_iena[28]
  PIN la_iena[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.270 816.000 498.550 820.000 ;
    END
  END la_iena[29]
  PIN la_iena[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 816.000 51.430 820.000 ;
    END
  END la_iena[2]
  PIN la_iena[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 514.830 816.000 515.110 820.000 ;
    END
  END la_iena[30]
  PIN la_iena[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 816.000 531.670 820.000 ;
    END
  END la_iena[31]
  PIN la_iena[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.950 816.000 548.230 820.000 ;
    END
  END la_iena[32]
  PIN la_iena[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 816.000 564.790 820.000 ;
    END
  END la_iena[33]
  PIN la_iena[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 816.000 581.350 820.000 ;
    END
  END la_iena[34]
  PIN la_iena[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 816.000 597.910 820.000 ;
    END
  END la_iena[35]
  PIN la_iena[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.190 816.000 614.470 820.000 ;
    END
  END la_iena[36]
  PIN la_iena[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.750 816.000 631.030 820.000 ;
    END
  END la_iena[37]
  PIN la_iena[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.310 816.000 647.590 820.000 ;
    END
  END la_iena[38]
  PIN la_iena[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.870 816.000 664.150 820.000 ;
    END
  END la_iena[39]
  PIN la_iena[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 816.000 67.990 820.000 ;
    END
  END la_iena[3]
  PIN la_iena[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 816.000 680.710 820.000 ;
    END
  END la_iena[40]
  PIN la_iena[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.990 816.000 697.270 820.000 ;
    END
  END la_iena[41]
  PIN la_iena[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.550 816.000 713.830 820.000 ;
    END
  END la_iena[42]
  PIN la_iena[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 816.000 730.390 820.000 ;
    END
  END la_iena[43]
  PIN la_iena[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.670 816.000 746.950 820.000 ;
    END
  END la_iena[44]
  PIN la_iena[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 816.000 763.510 820.000 ;
    END
  END la_iena[45]
  PIN la_iena[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.790 816.000 780.070 820.000 ;
    END
  END la_iena[46]
  PIN la_iena[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.350 816.000 796.630 820.000 ;
    END
  END la_iena[47]
  PIN la_iena[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.910 816.000 813.190 820.000 ;
    END
  END la_iena[48]
  PIN la_iena[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.470 816.000 829.750 820.000 ;
    END
  END la_iena[49]
  PIN la_iena[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.270 816.000 84.550 820.000 ;
    END
  END la_iena[4]
  PIN la_iena[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.030 816.000 846.310 820.000 ;
    END
  END la_iena[50]
  PIN la_iena[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.590 816.000 862.870 820.000 ;
    END
  END la_iena[51]
  PIN la_iena[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 816.000 879.430 820.000 ;
    END
  END la_iena[52]
  PIN la_iena[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.710 816.000 895.990 820.000 ;
    END
  END la_iena[53]
  PIN la_iena[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.270 816.000 912.550 820.000 ;
    END
  END la_iena[54]
  PIN la_iena[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 928.830 816.000 929.110 820.000 ;
    END
  END la_iena[55]
  PIN la_iena[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.390 816.000 945.670 820.000 ;
    END
  END la_iena[56]
  PIN la_iena[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 961.950 816.000 962.230 820.000 ;
    END
  END la_iena[57]
  PIN la_iena[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.510 816.000 978.790 820.000 ;
    END
  END la_iena[58]
  PIN la_iena[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.070 816.000 995.350 820.000 ;
    END
  END la_iena[59]
  PIN la_iena[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 100.830 816.000 101.110 820.000 ;
    END
  END la_iena[5]
  PIN la_iena[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.630 816.000 1011.910 820.000 ;
    END
  END la_iena[60]
  PIN la_iena[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1028.190 816.000 1028.470 820.000 ;
    END
  END la_iena[61]
  PIN la_iena[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1044.750 816.000 1045.030 820.000 ;
    END
  END la_iena[62]
  PIN la_iena[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.310 816.000 1061.590 820.000 ;
    END
  END la_iena[63]
  PIN la_iena[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1077.870 816.000 1078.150 820.000 ;
    END
  END la_iena[64]
  PIN la_iena[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.430 816.000 1094.710 820.000 ;
    END
  END la_iena[65]
  PIN la_iena[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.990 816.000 1111.270 820.000 ;
    END
  END la_iena[66]
  PIN la_iena[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.550 816.000 1127.830 820.000 ;
    END
  END la_iena[67]
  PIN la_iena[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1144.110 816.000 1144.390 820.000 ;
    END
  END la_iena[68]
  PIN la_iena[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.670 816.000 1160.950 820.000 ;
    END
  END la_iena[69]
  PIN la_iena[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.390 816.000 117.670 820.000 ;
    END
  END la_iena[6]
  PIN la_iena[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.230 816.000 1177.510 820.000 ;
    END
  END la_iena[70]
  PIN la_iena[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.070 816.000 1202.350 820.000 ;
    END
  END la_iena[71]
  PIN la_iena[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.630 816.000 1218.910 820.000 ;
    END
  END la_iena[72]
  PIN la_iena[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1235.190 816.000 1235.470 820.000 ;
    END
  END la_iena[73]
  PIN la_iena[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1251.750 816.000 1252.030 820.000 ;
    END
  END la_iena[74]
  PIN la_iena[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.310 816.000 1268.590 820.000 ;
    END
  END la_iena[75]
  PIN la_iena[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1284.870 816.000 1285.150 820.000 ;
    END
  END la_iena[76]
  PIN la_iena[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.430 816.000 1301.710 820.000 ;
    END
  END la_iena[77]
  PIN la_iena[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1317.990 816.000 1318.270 820.000 ;
    END
  END la_iena[78]
  PIN la_iena[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1334.550 816.000 1334.830 820.000 ;
    END
  END la_iena[79]
  PIN la_iena[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 816.000 134.230 820.000 ;
    END
  END la_iena[7]
  PIN la_iena[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1351.110 816.000 1351.390 820.000 ;
    END
  END la_iena[80]
  PIN la_iena[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.670 816.000 1367.950 820.000 ;
    END
  END la_iena[81]
  PIN la_iena[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1384.230 816.000 1384.510 820.000 ;
    END
  END la_iena[82]
  PIN la_iena[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.790 816.000 1401.070 820.000 ;
    END
  END la_iena[83]
  PIN la_iena[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.350 816.000 1417.630 820.000 ;
    END
  END la_iena[84]
  PIN la_iena[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1433.910 816.000 1434.190 820.000 ;
    END
  END la_iena[85]
  PIN la_iena[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.470 816.000 1450.750 820.000 ;
    END
  END la_iena[86]
  PIN la_iena[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.030 816.000 1467.310 820.000 ;
    END
  END la_iena[87]
  PIN la_iena[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1483.590 816.000 1483.870 820.000 ;
    END
  END la_iena[88]
  PIN la_iena[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.150 816.000 1500.430 820.000 ;
    END
  END la_iena[89]
  PIN la_iena[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 816.000 150.790 820.000 ;
    END
  END la_iena[8]
  PIN la_iena[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1516.710 816.000 1516.990 820.000 ;
    END
  END la_iena[90]
  PIN la_iena[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.270 816.000 1533.550 820.000 ;
    END
  END la_iena[91]
  PIN la_iena[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1549.830 816.000 1550.110 820.000 ;
    END
  END la_iena[92]
  PIN la_iena[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1566.390 816.000 1566.670 820.000 ;
    END
  END la_iena[93]
  PIN la_iena[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1582.950 816.000 1583.230 820.000 ;
    END
  END la_iena[94]
  PIN la_iena[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1599.510 816.000 1599.790 820.000 ;
    END
  END la_iena[95]
  PIN la_iena[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.070 816.000 1616.350 820.000 ;
    END
  END la_iena[96]
  PIN la_iena[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.630 816.000 1632.910 820.000 ;
    END
  END la_iena[97]
  PIN la_iena[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1649.190 816.000 1649.470 820.000 ;
    END
  END la_iena[98]
  PIN la_iena[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1665.750 816.000 1666.030 820.000 ;
    END
  END la_iena[99]
  PIN la_iena[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 816.000 167.350 820.000 ;
    END
  END la_iena[9]
  PIN la_input[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.170 816.000 22.450 820.000 ;
    END
  END la_input[0]
  PIN la_input[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1686.450 816.000 1686.730 820.000 ;
    END
  END la_input[100]
  PIN la_input[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1703.010 816.000 1703.290 820.000 ;
    END
  END la_input[101]
  PIN la_input[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1719.570 816.000 1719.850 820.000 ;
    END
  END la_input[102]
  PIN la_input[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1736.130 816.000 1736.410 820.000 ;
    END
  END la_input[103]
  PIN la_input[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.690 816.000 1752.970 820.000 ;
    END
  END la_input[104]
  PIN la_input[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1769.250 816.000 1769.530 820.000 ;
    END
  END la_input[105]
  PIN la_input[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1785.810 816.000 1786.090 820.000 ;
    END
  END la_input[106]
  PIN la_input[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1802.370 816.000 1802.650 820.000 ;
    END
  END la_input[107]
  PIN la_input[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1818.930 816.000 1819.210 820.000 ;
    END
  END la_input[108]
  PIN la_input[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1835.490 816.000 1835.770 820.000 ;
    END
  END la_input[109]
  PIN la_input[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 816.000 188.050 820.000 ;
    END
  END la_input[10]
  PIN la_input[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.050 816.000 1852.330 820.000 ;
    END
  END la_input[110]
  PIN la_input[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1868.610 816.000 1868.890 820.000 ;
    END
  END la_input[111]
  PIN la_input[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1885.170 816.000 1885.450 820.000 ;
    END
  END la_input[112]
  PIN la_input[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1901.730 816.000 1902.010 820.000 ;
    END
  END la_input[113]
  PIN la_input[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1918.290 816.000 1918.570 820.000 ;
    END
  END la_input[114]
  PIN la_input[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1934.850 816.000 1935.130 820.000 ;
    END
  END la_input[115]
  PIN la_input[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1951.410 816.000 1951.690 820.000 ;
    END
  END la_input[116]
  PIN la_input[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1967.970 816.000 1968.250 820.000 ;
    END
  END la_input[117]
  PIN la_input[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1984.530 816.000 1984.810 820.000 ;
    END
  END la_input[118]
  PIN la_input[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2001.090 816.000 2001.370 820.000 ;
    END
  END la_input[119]
  PIN la_input[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.330 816.000 204.610 820.000 ;
    END
  END la_input[11]
  PIN la_input[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.650 816.000 2017.930 820.000 ;
    END
  END la_input[120]
  PIN la_input[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2034.210 816.000 2034.490 820.000 ;
    END
  END la_input[121]
  PIN la_input[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2050.770 816.000 2051.050 820.000 ;
    END
  END la_input[122]
  PIN la_input[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2067.330 816.000 2067.610 820.000 ;
    END
  END la_input[123]
  PIN la_input[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.890 816.000 2084.170 820.000 ;
    END
  END la_input[124]
  PIN la_input[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.450 816.000 2100.730 820.000 ;
    END
  END la_input[125]
  PIN la_input[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2117.010 816.000 2117.290 820.000 ;
    END
  END la_input[126]
  PIN la_input[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2133.570 816.000 2133.850 820.000 ;
    END
  END la_input[127]
  PIN la_input[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 816.000 221.170 820.000 ;
    END
  END la_input[12]
  PIN la_input[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 816.000 237.730 820.000 ;
    END
  END la_input[13]
  PIN la_input[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 816.000 254.290 820.000 ;
    END
  END la_input[14]
  PIN la_input[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 816.000 270.850 820.000 ;
    END
  END la_input[15]
  PIN la_input[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 816.000 287.410 820.000 ;
    END
  END la_input[16]
  PIN la_input[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 816.000 303.970 820.000 ;
    END
  END la_input[17]
  PIN la_input[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 816.000 320.530 820.000 ;
    END
  END la_input[18]
  PIN la_input[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.810 816.000 337.090 820.000 ;
    END
  END la_input[19]
  PIN la_input[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 816.000 39.010 820.000 ;
    END
  END la_input[1]
  PIN la_input[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 816.000 353.650 820.000 ;
    END
  END la_input[20]
  PIN la_input[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.930 816.000 370.210 820.000 ;
    END
  END la_input[21]
  PIN la_input[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 816.000 386.770 820.000 ;
    END
  END la_input[22]
  PIN la_input[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 816.000 403.330 820.000 ;
    END
  END la_input[23]
  PIN la_input[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.610 816.000 419.890 820.000 ;
    END
  END la_input[24]
  PIN la_input[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.170 816.000 436.450 820.000 ;
    END
  END la_input[25]
  PIN la_input[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.730 816.000 453.010 820.000 ;
    END
  END la_input[26]
  PIN la_input[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.290 816.000 469.570 820.000 ;
    END
  END la_input[27]
  PIN la_input[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 816.000 486.130 820.000 ;
    END
  END la_input[28]
  PIN la_input[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 816.000 502.690 820.000 ;
    END
  END la_input[29]
  PIN la_input[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.290 816.000 55.570 820.000 ;
    END
  END la_input[2]
  PIN la_input[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 816.000 519.250 820.000 ;
    END
  END la_input[30]
  PIN la_input[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.530 816.000 535.810 820.000 ;
    END
  END la_input[31]
  PIN la_input[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.090 816.000 552.370 820.000 ;
    END
  END la_input[32]
  PIN la_input[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.650 816.000 568.930 820.000 ;
    END
  END la_input[33]
  PIN la_input[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.210 816.000 585.490 820.000 ;
    END
  END la_input[34]
  PIN la_input[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.770 816.000 602.050 820.000 ;
    END
  END la_input[35]
  PIN la_input[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.330 816.000 618.610 820.000 ;
    END
  END la_input[36]
  PIN la_input[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.890 816.000 635.170 820.000 ;
    END
  END la_input[37]
  PIN la_input[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.450 816.000 651.730 820.000 ;
    END
  END la_input[38]
  PIN la_input[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.010 816.000 668.290 820.000 ;
    END
  END la_input[39]
  PIN la_input[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 816.000 72.130 820.000 ;
    END
  END la_input[3]
  PIN la_input[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.570 816.000 684.850 820.000 ;
    END
  END la_input[40]
  PIN la_input[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.130 816.000 701.410 820.000 ;
    END
  END la_input[41]
  PIN la_input[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.690 816.000 717.970 820.000 ;
    END
  END la_input[42]
  PIN la_input[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 816.000 734.530 820.000 ;
    END
  END la_input[43]
  PIN la_input[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.810 816.000 751.090 820.000 ;
    END
  END la_input[44]
  PIN la_input[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.370 816.000 767.650 820.000 ;
    END
  END la_input[45]
  PIN la_input[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.930 816.000 784.210 820.000 ;
    END
  END la_input[46]
  PIN la_input[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.490 816.000 800.770 820.000 ;
    END
  END la_input[47]
  PIN la_input[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.050 816.000 817.330 820.000 ;
    END
  END la_input[48]
  PIN la_input[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.610 816.000 833.890 820.000 ;
    END
  END la_input[49]
  PIN la_input[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 816.000 88.690 820.000 ;
    END
  END la_input[4]
  PIN la_input[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 816.000 850.450 820.000 ;
    END
  END la_input[50]
  PIN la_input[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.730 816.000 867.010 820.000 ;
    END
  END la_input[51]
  PIN la_input[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.290 816.000 883.570 820.000 ;
    END
  END la_input[52]
  PIN la_input[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.850 816.000 900.130 820.000 ;
    END
  END la_input[53]
  PIN la_input[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 916.410 816.000 916.690 820.000 ;
    END
  END la_input[54]
  PIN la_input[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.970 816.000 933.250 820.000 ;
    END
  END la_input[55]
  PIN la_input[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.530 816.000 949.810 820.000 ;
    END
  END la_input[56]
  PIN la_input[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 816.000 966.370 820.000 ;
    END
  END la_input[57]
  PIN la_input[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.650 816.000 982.930 820.000 ;
    END
  END la_input[58]
  PIN la_input[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.210 816.000 999.490 820.000 ;
    END
  END la_input[59]
  PIN la_input[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 816.000 105.250 820.000 ;
    END
  END la_input[5]
  PIN la_input[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.770 816.000 1016.050 820.000 ;
    END
  END la_input[60]
  PIN la_input[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1032.330 816.000 1032.610 820.000 ;
    END
  END la_input[61]
  PIN la_input[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.890 816.000 1049.170 820.000 ;
    END
  END la_input[62]
  PIN la_input[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.450 816.000 1065.730 820.000 ;
    END
  END la_input[63]
  PIN la_input[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1082.010 816.000 1082.290 820.000 ;
    END
  END la_input[64]
  PIN la_input[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1098.570 816.000 1098.850 820.000 ;
    END
  END la_input[65]
  PIN la_input[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1115.130 816.000 1115.410 820.000 ;
    END
  END la_input[66]
  PIN la_input[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.690 816.000 1131.970 820.000 ;
    END
  END la_input[67]
  PIN la_input[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1148.250 816.000 1148.530 820.000 ;
    END
  END la_input[68]
  PIN la_input[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.810 816.000 1165.090 820.000 ;
    END
  END la_input[69]
  PIN la_input[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 816.000 121.810 820.000 ;
    END
  END la_input[6]
  PIN la_input[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.370 816.000 1181.650 820.000 ;
    END
  END la_input[70]
  PIN la_input[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1206.210 816.000 1206.490 820.000 ;
    END
  END la_input[71]
  PIN la_input[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1222.770 816.000 1223.050 820.000 ;
    END
  END la_input[72]
  PIN la_input[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1239.330 816.000 1239.610 820.000 ;
    END
  END la_input[73]
  PIN la_input[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.890 816.000 1256.170 820.000 ;
    END
  END la_input[74]
  PIN la_input[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1272.450 816.000 1272.730 820.000 ;
    END
  END la_input[75]
  PIN la_input[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.010 816.000 1289.290 820.000 ;
    END
  END la_input[76]
  PIN la_input[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1305.570 816.000 1305.850 820.000 ;
    END
  END la_input[77]
  PIN la_input[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1322.130 816.000 1322.410 820.000 ;
    END
  END la_input[78]
  PIN la_input[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.690 816.000 1338.970 820.000 ;
    END
  END la_input[79]
  PIN la_input[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.090 816.000 138.370 820.000 ;
    END
  END la_input[7]
  PIN la_input[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1355.250 816.000 1355.530 820.000 ;
    END
  END la_input[80]
  PIN la_input[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.810 816.000 1372.090 820.000 ;
    END
  END la_input[81]
  PIN la_input[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1388.370 816.000 1388.650 820.000 ;
    END
  END la_input[82]
  PIN la_input[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.930 816.000 1405.210 820.000 ;
    END
  END la_input[83]
  PIN la_input[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.490 816.000 1421.770 820.000 ;
    END
  END la_input[84]
  PIN la_input[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.050 816.000 1438.330 820.000 ;
    END
  END la_input[85]
  PIN la_input[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1454.610 816.000 1454.890 820.000 ;
    END
  END la_input[86]
  PIN la_input[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.170 816.000 1471.450 820.000 ;
    END
  END la_input[87]
  PIN la_input[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1487.730 816.000 1488.010 820.000 ;
    END
  END la_input[88]
  PIN la_input[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1504.290 816.000 1504.570 820.000 ;
    END
  END la_input[89]
  PIN la_input[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 816.000 154.930 820.000 ;
    END
  END la_input[8]
  PIN la_input[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1520.850 816.000 1521.130 820.000 ;
    END
  END la_input[90]
  PIN la_input[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1537.410 816.000 1537.690 820.000 ;
    END
  END la_input[91]
  PIN la_input[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1553.970 816.000 1554.250 820.000 ;
    END
  END la_input[92]
  PIN la_input[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1570.530 816.000 1570.810 820.000 ;
    END
  END la_input[93]
  PIN la_input[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1587.090 816.000 1587.370 820.000 ;
    END
  END la_input[94]
  PIN la_input[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.650 816.000 1603.930 820.000 ;
    END
  END la_input[95]
  PIN la_input[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1620.210 816.000 1620.490 820.000 ;
    END
  END la_input[96]
  PIN la_input[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1636.770 816.000 1637.050 820.000 ;
    END
  END la_input[97]
  PIN la_input[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1653.330 816.000 1653.610 820.000 ;
    END
  END la_input[98]
  PIN la_input[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.890 816.000 1670.170 820.000 ;
    END
  END la_input[99]
  PIN la_input[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.210 816.000 171.490 820.000 ;
    END
  END la_input[9]
  PIN la_oenb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 816.000 26.590 820.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1690.590 816.000 1690.870 820.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1707.150 816.000 1707.430 820.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1723.710 816.000 1723.990 820.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.270 816.000 1740.550 820.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1756.830 816.000 1757.110 820.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1773.390 816.000 1773.670 820.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1789.950 816.000 1790.230 820.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1806.510 816.000 1806.790 820.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1823.070 816.000 1823.350 820.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1839.630 816.000 1839.910 820.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 816.000 192.190 820.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1856.190 816.000 1856.470 820.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1872.750 816.000 1873.030 820.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1889.310 816.000 1889.590 820.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.870 816.000 1906.150 820.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.430 816.000 1922.710 820.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.990 816.000 1939.270 820.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1955.550 816.000 1955.830 820.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1972.110 816.000 1972.390 820.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.670 816.000 1988.950 820.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2005.230 816.000 2005.510 820.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 816.000 208.750 820.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2021.790 816.000 2022.070 820.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2038.350 816.000 2038.630 820.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2054.910 816.000 2055.190 820.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.470 816.000 2071.750 820.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2088.030 816.000 2088.310 820.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2104.590 816.000 2104.870 820.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2121.150 816.000 2121.430 820.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2137.710 816.000 2137.990 820.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 816.000 225.310 820.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 816.000 241.870 820.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 816.000 258.430 820.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 816.000 274.990 820.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.270 816.000 291.550 820.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 816.000 308.110 820.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.390 816.000 324.670 820.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 816.000 341.230 820.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 816.000 43.150 820.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 816.000 357.790 820.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 816.000 374.350 820.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.630 816.000 390.910 820.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 816.000 407.470 820.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.750 816.000 424.030 820.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 816.000 440.590 820.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 816.000 457.150 820.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 816.000 473.710 820.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.990 816.000 490.270 820.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 816.000 506.830 820.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 816.000 59.710 820.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.110 816.000 523.390 820.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.670 816.000 539.950 820.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 816.000 556.510 820.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 816.000 573.070 820.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.350 816.000 589.630 820.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 816.000 606.190 820.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 816.000 622.750 820.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 816.000 639.310 820.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.590 816.000 655.870 820.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.150 816.000 672.430 820.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 816.000 76.270 820.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.710 816.000 688.990 820.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 816.000 705.550 820.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 721.830 816.000 722.110 820.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.390 816.000 738.670 820.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.950 816.000 755.230 820.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 816.000 771.790 820.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.070 816.000 788.350 820.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.630 816.000 804.910 820.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 816.000 821.470 820.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.750 816.000 838.030 820.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 816.000 92.830 820.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.310 816.000 854.590 820.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.870 816.000 871.150 820.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.430 816.000 887.710 820.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.990 816.000 904.270 820.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.550 816.000 920.830 820.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 816.000 937.390 820.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.670 816.000 953.950 820.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.230 816.000 970.510 820.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.790 816.000 987.070 820.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1003.350 816.000 1003.630 820.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 816.000 109.390 820.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.910 816.000 1020.190 820.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.470 816.000 1036.750 820.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.030 816.000 1053.310 820.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.590 816.000 1069.870 820.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.150 816.000 1086.430 820.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.710 816.000 1102.990 820.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.270 816.000 1119.550 820.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1135.830 816.000 1136.110 820.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.390 816.000 1152.670 820.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.950 816.000 1169.230 820.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 816.000 125.950 820.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.510 816.000 1185.790 820.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.350 816.000 1210.630 820.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1226.910 816.000 1227.190 820.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.470 816.000 1243.750 820.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.030 816.000 1260.310 820.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1276.590 816.000 1276.870 820.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.150 816.000 1293.430 820.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1309.710 816.000 1309.990 820.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.270 816.000 1326.550 820.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1342.830 816.000 1343.110 820.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 816.000 142.510 820.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1359.390 816.000 1359.670 820.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.950 816.000 1376.230 820.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1392.510 816.000 1392.790 820.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.070 816.000 1409.350 820.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1425.630 816.000 1425.910 820.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.190 816.000 1442.470 820.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.750 816.000 1459.030 820.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.310 816.000 1475.590 820.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1491.870 816.000 1492.150 820.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1508.430 816.000 1508.710 820.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 816.000 159.070 820.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1524.990 816.000 1525.270 820.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1541.550 816.000 1541.830 820.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1558.110 816.000 1558.390 820.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.670 816.000 1574.950 820.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1591.230 816.000 1591.510 820.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1607.790 816.000 1608.070 820.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1624.350 816.000 1624.630 820.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1640.910 816.000 1641.190 820.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.470 816.000 1657.750 820.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.030 816.000 1674.310 820.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 816.000 175.630 820.000 ;
    END
  END la_oenb[9]
  PIN la_output[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 816.000 30.730 820.000 ;
    END
  END la_output[0]
  PIN la_output[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1694.730 816.000 1695.010 820.000 ;
    END
  END la_output[100]
  PIN la_output[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1711.290 816.000 1711.570 820.000 ;
    END
  END la_output[101]
  PIN la_output[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.850 816.000 1728.130 820.000 ;
    END
  END la_output[102]
  PIN la_output[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1744.410 816.000 1744.690 820.000 ;
    END
  END la_output[103]
  PIN la_output[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.970 816.000 1761.250 820.000 ;
    END
  END la_output[104]
  PIN la_output[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.530 816.000 1777.810 820.000 ;
    END
  END la_output[105]
  PIN la_output[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1794.090 816.000 1794.370 820.000 ;
    END
  END la_output[106]
  PIN la_output[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.650 816.000 1810.930 820.000 ;
    END
  END la_output[107]
  PIN la_output[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1827.210 816.000 1827.490 820.000 ;
    END
  END la_output[108]
  PIN la_output[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1843.770 816.000 1844.050 820.000 ;
    END
  END la_output[109]
  PIN la_output[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 816.000 196.330 820.000 ;
    END
  END la_output[10]
  PIN la_output[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1860.330 816.000 1860.610 820.000 ;
    END
  END la_output[110]
  PIN la_output[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.890 816.000 1877.170 820.000 ;
    END
  END la_output[111]
  PIN la_output[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1893.450 816.000 1893.730 820.000 ;
    END
  END la_output[112]
  PIN la_output[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1910.010 816.000 1910.290 820.000 ;
    END
  END la_output[113]
  PIN la_output[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1926.570 816.000 1926.850 820.000 ;
    END
  END la_output[114]
  PIN la_output[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1943.130 816.000 1943.410 820.000 ;
    END
  END la_output[115]
  PIN la_output[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.690 816.000 1959.970 820.000 ;
    END
  END la_output[116]
  PIN la_output[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.250 816.000 1976.530 820.000 ;
    END
  END la_output[117]
  PIN la_output[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1992.810 816.000 1993.090 820.000 ;
    END
  END la_output[118]
  PIN la_output[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2009.370 816.000 2009.650 820.000 ;
    END
  END la_output[119]
  PIN la_output[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 816.000 212.890 820.000 ;
    END
  END la_output[11]
  PIN la_output[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2025.930 816.000 2026.210 820.000 ;
    END
  END la_output[120]
  PIN la_output[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2042.490 816.000 2042.770 820.000 ;
    END
  END la_output[121]
  PIN la_output[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.050 816.000 2059.330 820.000 ;
    END
  END la_output[122]
  PIN la_output[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2075.610 816.000 2075.890 820.000 ;
    END
  END la_output[123]
  PIN la_output[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2092.170 816.000 2092.450 820.000 ;
    END
  END la_output[124]
  PIN la_output[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2108.730 816.000 2109.010 820.000 ;
    END
  END la_output[125]
  PIN la_output[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2125.290 816.000 2125.570 820.000 ;
    END
  END la_output[126]
  PIN la_output[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2141.850 816.000 2142.130 820.000 ;
    END
  END la_output[127]
  PIN la_output[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 816.000 229.450 820.000 ;
    END
  END la_output[12]
  PIN la_output[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.730 816.000 246.010 820.000 ;
    END
  END la_output[13]
  PIN la_output[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 816.000 262.570 820.000 ;
    END
  END la_output[14]
  PIN la_output[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 816.000 279.130 820.000 ;
    END
  END la_output[15]
  PIN la_output[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 816.000 295.690 820.000 ;
    END
  END la_output[16]
  PIN la_output[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.970 816.000 312.250 820.000 ;
    END
  END la_output[17]
  PIN la_output[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 816.000 328.810 820.000 ;
    END
  END la_output[18]
  PIN la_output[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 816.000 345.370 820.000 ;
    END
  END la_output[19]
  PIN la_output[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 47.010 816.000 47.290 820.000 ;
    END
  END la_output[1]
  PIN la_output[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 816.000 361.930 820.000 ;
    END
  END la_output[20]
  PIN la_output[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 816.000 378.490 820.000 ;
    END
  END la_output[21]
  PIN la_output[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 816.000 395.050 820.000 ;
    END
  END la_output[22]
  PIN la_output[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 816.000 411.610 820.000 ;
    END
  END la_output[23]
  PIN la_output[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 816.000 428.170 820.000 ;
    END
  END la_output[24]
  PIN la_output[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 816.000 444.730 820.000 ;
    END
  END la_output[25]
  PIN la_output[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 816.000 461.290 820.000 ;
    END
  END la_output[26]
  PIN la_output[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.570 816.000 477.850 820.000 ;
    END
  END la_output[27]
  PIN la_output[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.130 816.000 494.410 820.000 ;
    END
  END la_output[28]
  PIN la_output[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.690 816.000 510.970 820.000 ;
    END
  END la_output[29]
  PIN la_output[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 816.000 63.850 820.000 ;
    END
  END la_output[2]
  PIN la_output[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.250 816.000 527.530 820.000 ;
    END
  END la_output[30]
  PIN la_output[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.810 816.000 544.090 820.000 ;
    END
  END la_output[31]
  PIN la_output[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 816.000 560.650 820.000 ;
    END
  END la_output[32]
  PIN la_output[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 816.000 577.210 820.000 ;
    END
  END la_output[33]
  PIN la_output[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 816.000 593.770 820.000 ;
    END
  END la_output[34]
  PIN la_output[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.050 816.000 610.330 820.000 ;
    END
  END la_output[35]
  PIN la_output[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.610 816.000 626.890 820.000 ;
    END
  END la_output[36]
  PIN la_output[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 816.000 643.450 820.000 ;
    END
  END la_output[37]
  PIN la_output[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.730 816.000 660.010 820.000 ;
    END
  END la_output[38]
  PIN la_output[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.290 816.000 676.570 820.000 ;
    END
  END la_output[39]
  PIN la_output[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.130 816.000 80.410 820.000 ;
    END
  END la_output[3]
  PIN la_output[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.850 816.000 693.130 820.000 ;
    END
  END la_output[40]
  PIN la_output[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 709.410 816.000 709.690 820.000 ;
    END
  END la_output[41]
  PIN la_output[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.970 816.000 726.250 820.000 ;
    END
  END la_output[42]
  PIN la_output[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.530 816.000 742.810 820.000 ;
    END
  END la_output[43]
  PIN la_output[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 816.000 759.370 820.000 ;
    END
  END la_output[44]
  PIN la_output[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.650 816.000 775.930 820.000 ;
    END
  END la_output[45]
  PIN la_output[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 816.000 792.490 820.000 ;
    END
  END la_output[46]
  PIN la_output[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.770 816.000 809.050 820.000 ;
    END
  END la_output[47]
  PIN la_output[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 825.330 816.000 825.610 820.000 ;
    END
  END la_output[48]
  PIN la_output[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.890 816.000 842.170 820.000 ;
    END
  END la_output[49]
  PIN la_output[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 816.000 96.970 820.000 ;
    END
  END la_output[4]
  PIN la_output[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 858.450 816.000 858.730 820.000 ;
    END
  END la_output[50]
  PIN la_output[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.010 816.000 875.290 820.000 ;
    END
  END la_output[51]
  PIN la_output[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 891.570 816.000 891.850 820.000 ;
    END
  END la_output[52]
  PIN la_output[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.130 816.000 908.410 820.000 ;
    END
  END la_output[53]
  PIN la_output[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.690 816.000 924.970 820.000 ;
    END
  END la_output[54]
  PIN la_output[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.250 816.000 941.530 820.000 ;
    END
  END la_output[55]
  PIN la_output[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.810 816.000 958.090 820.000 ;
    END
  END la_output[56]
  PIN la_output[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 974.370 816.000 974.650 820.000 ;
    END
  END la_output[57]
  PIN la_output[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.930 816.000 991.210 820.000 ;
    END
  END la_output[58]
  PIN la_output[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.490 816.000 1007.770 820.000 ;
    END
  END la_output[59]
  PIN la_output[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 816.000 113.530 820.000 ;
    END
  END la_output[5]
  PIN la_output[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1024.050 816.000 1024.330 820.000 ;
    END
  END la_output[60]
  PIN la_output[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.610 816.000 1040.890 820.000 ;
    END
  END la_output[61]
  PIN la_output[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1057.170 816.000 1057.450 820.000 ;
    END
  END la_output[62]
  PIN la_output[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.730 816.000 1074.010 820.000 ;
    END
  END la_output[63]
  PIN la_output[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.290 816.000 1090.570 820.000 ;
    END
  END la_output[64]
  PIN la_output[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.850 816.000 1107.130 820.000 ;
    END
  END la_output[65]
  PIN la_output[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.410 816.000 1123.690 820.000 ;
    END
  END la_output[66]
  PIN la_output[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.970 816.000 1140.250 820.000 ;
    END
  END la_output[67]
  PIN la_output[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1156.530 816.000 1156.810 820.000 ;
    END
  END la_output[68]
  PIN la_output[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1173.090 816.000 1173.370 820.000 ;
    END
  END la_output[69]
  PIN la_output[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 816.000 130.090 820.000 ;
    END
  END la_output[6]
  PIN la_output[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1189.650 816.000 1189.930 820.000 ;
    END
  END la_output[70]
  PIN la_output[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.490 816.000 1214.770 820.000 ;
    END
  END la_output[71]
  PIN la_output[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.050 816.000 1231.330 820.000 ;
    END
  END la_output[72]
  PIN la_output[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.610 816.000 1247.890 820.000 ;
    END
  END la_output[73]
  PIN la_output[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.170 816.000 1264.450 820.000 ;
    END
  END la_output[74]
  PIN la_output[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.730 816.000 1281.010 820.000 ;
    END
  END la_output[75]
  PIN la_output[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.290 816.000 1297.570 820.000 ;
    END
  END la_output[76]
  PIN la_output[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.850 816.000 1314.130 820.000 ;
    END
  END la_output[77]
  PIN la_output[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1330.410 816.000 1330.690 820.000 ;
    END
  END la_output[78]
  PIN la_output[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.970 816.000 1347.250 820.000 ;
    END
  END la_output[79]
  PIN la_output[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 146.370 816.000 146.650 820.000 ;
    END
  END la_output[7]
  PIN la_output[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.530 816.000 1363.810 820.000 ;
    END
  END la_output[80]
  PIN la_output[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.090 816.000 1380.370 820.000 ;
    END
  END la_output[81]
  PIN la_output[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.650 816.000 1396.930 820.000 ;
    END
  END la_output[82]
  PIN la_output[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1413.210 816.000 1413.490 820.000 ;
    END
  END la_output[83]
  PIN la_output[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.770 816.000 1430.050 820.000 ;
    END
  END la_output[84]
  PIN la_output[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1446.330 816.000 1446.610 820.000 ;
    END
  END la_output[85]
  PIN la_output[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.890 816.000 1463.170 820.000 ;
    END
  END la_output[86]
  PIN la_output[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1479.450 816.000 1479.730 820.000 ;
    END
  END la_output[87]
  PIN la_output[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.010 816.000 1496.290 820.000 ;
    END
  END la_output[88]
  PIN la_output[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1512.570 816.000 1512.850 820.000 ;
    END
  END la_output[89]
  PIN la_output[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 816.000 163.210 820.000 ;
    END
  END la_output[8]
  PIN la_output[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1529.130 816.000 1529.410 820.000 ;
    END
  END la_output[90]
  PIN la_output[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.690 816.000 1545.970 820.000 ;
    END
  END la_output[91]
  PIN la_output[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1562.250 816.000 1562.530 820.000 ;
    END
  END la_output[92]
  PIN la_output[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1578.810 816.000 1579.090 820.000 ;
    END
  END la_output[93]
  PIN la_output[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1595.370 816.000 1595.650 820.000 ;
    END
  END la_output[94]
  PIN la_output[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.930 816.000 1612.210 820.000 ;
    END
  END la_output[95]
  PIN la_output[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1628.490 816.000 1628.770 820.000 ;
    END
  END la_output[96]
  PIN la_output[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.050 816.000 1645.330 820.000 ;
    END
  END la_output[97]
  PIN la_output[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.610 816.000 1661.890 820.000 ;
    END
  END la_output[98]
  PIN la_output[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1678.170 816.000 1678.450 820.000 ;
    END
  END la_output[99]
  PIN la_output[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.490 816.000 179.770 820.000 ;
    END
  END la_output[9]
  PIN mprj_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2145.990 816.000 2146.270 820.000 ;
    END
  END mprj_ack_i
  PIN mprj_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2166.690 816.000 2166.970 820.000 ;
    END
  END mprj_adr_o[0]
  PIN mprj_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2307.450 816.000 2307.730 820.000 ;
    END
  END mprj_adr_o[10]
  PIN mprj_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2319.870 816.000 2320.150 820.000 ;
    END
  END mprj_adr_o[11]
  PIN mprj_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2332.290 816.000 2332.570 820.000 ;
    END
  END mprj_adr_o[12]
  PIN mprj_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2344.710 816.000 2344.990 820.000 ;
    END
  END mprj_adr_o[13]
  PIN mprj_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2357.130 816.000 2357.410 820.000 ;
    END
  END mprj_adr_o[14]
  PIN mprj_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2369.550 816.000 2369.830 820.000 ;
    END
  END mprj_adr_o[15]
  PIN mprj_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2381.970 816.000 2382.250 820.000 ;
    END
  END mprj_adr_o[16]
  PIN mprj_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2394.390 816.000 2394.670 820.000 ;
    END
  END mprj_adr_o[17]
  PIN mprj_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2406.810 816.000 2407.090 820.000 ;
    END
  END mprj_adr_o[18]
  PIN mprj_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2419.230 816.000 2419.510 820.000 ;
    END
  END mprj_adr_o[19]
  PIN mprj_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.250 816.000 2183.530 820.000 ;
    END
  END mprj_adr_o[1]
  PIN mprj_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.650 816.000 2431.930 820.000 ;
    END
  END mprj_adr_o[20]
  PIN mprj_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2444.070 816.000 2444.350 820.000 ;
    END
  END mprj_adr_o[21]
  PIN mprj_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2456.490 816.000 2456.770 820.000 ;
    END
  END mprj_adr_o[22]
  PIN mprj_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2468.910 816.000 2469.190 820.000 ;
    END
  END mprj_adr_o[23]
  PIN mprj_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2481.330 816.000 2481.610 820.000 ;
    END
  END mprj_adr_o[24]
  PIN mprj_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2493.750 816.000 2494.030 820.000 ;
    END
  END mprj_adr_o[25]
  PIN mprj_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2506.170 816.000 2506.450 820.000 ;
    END
  END mprj_adr_o[26]
  PIN mprj_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2518.590 816.000 2518.870 820.000 ;
    END
  END mprj_adr_o[27]
  PIN mprj_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2531.010 816.000 2531.290 820.000 ;
    END
  END mprj_adr_o[28]
  PIN mprj_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2543.430 816.000 2543.710 820.000 ;
    END
  END mprj_adr_o[29]
  PIN mprj_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2199.810 816.000 2200.090 820.000 ;
    END
  END mprj_adr_o[2]
  PIN mprj_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2555.850 816.000 2556.130 820.000 ;
    END
  END mprj_adr_o[30]
  PIN mprj_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2568.270 816.000 2568.550 820.000 ;
    END
  END mprj_adr_o[31]
  PIN mprj_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2216.370 816.000 2216.650 820.000 ;
    END
  END mprj_adr_o[3]
  PIN mprj_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2232.930 816.000 2233.210 820.000 ;
    END
  END mprj_adr_o[4]
  PIN mprj_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2245.350 816.000 2245.630 820.000 ;
    END
  END mprj_adr_o[5]
  PIN mprj_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2257.770 816.000 2258.050 820.000 ;
    END
  END mprj_adr_o[6]
  PIN mprj_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2270.190 816.000 2270.470 820.000 ;
    END
  END mprj_adr_o[7]
  PIN mprj_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2282.610 816.000 2282.890 820.000 ;
    END
  END mprj_adr_o[8]
  PIN mprj_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.030 816.000 2295.310 820.000 ;
    END
  END mprj_adr_o[9]
  PIN mprj_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2150.130 816.000 2150.410 820.000 ;
    END
  END mprj_cyc_o
  PIN mprj_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2170.830 816.000 2171.110 820.000 ;
    END
  END mprj_dat_i[0]
  PIN mprj_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.590 816.000 2311.870 820.000 ;
    END
  END mprj_dat_i[10]
  PIN mprj_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2324.010 816.000 2324.290 820.000 ;
    END
  END mprj_dat_i[11]
  PIN mprj_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2336.430 816.000 2336.710 820.000 ;
    END
  END mprj_dat_i[12]
  PIN mprj_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2348.850 816.000 2349.130 820.000 ;
    END
  END mprj_dat_i[13]
  PIN mprj_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.270 816.000 2361.550 820.000 ;
    END
  END mprj_dat_i[14]
  PIN mprj_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2373.690 816.000 2373.970 820.000 ;
    END
  END mprj_dat_i[15]
  PIN mprj_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2386.110 816.000 2386.390 820.000 ;
    END
  END mprj_dat_i[16]
  PIN mprj_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2398.530 816.000 2398.810 820.000 ;
    END
  END mprj_dat_i[17]
  PIN mprj_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2410.950 816.000 2411.230 820.000 ;
    END
  END mprj_dat_i[18]
  PIN mprj_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2423.370 816.000 2423.650 820.000 ;
    END
  END mprj_dat_i[19]
  PIN mprj_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2187.390 816.000 2187.670 820.000 ;
    END
  END mprj_dat_i[1]
  PIN mprj_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2435.790 816.000 2436.070 820.000 ;
    END
  END mprj_dat_i[20]
  PIN mprj_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2448.210 816.000 2448.490 820.000 ;
    END
  END mprj_dat_i[21]
  PIN mprj_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2460.630 816.000 2460.910 820.000 ;
    END
  END mprj_dat_i[22]
  PIN mprj_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.050 816.000 2473.330 820.000 ;
    END
  END mprj_dat_i[23]
  PIN mprj_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.470 816.000 2485.750 820.000 ;
    END
  END mprj_dat_i[24]
  PIN mprj_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2497.890 816.000 2498.170 820.000 ;
    END
  END mprj_dat_i[25]
  PIN mprj_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2510.310 816.000 2510.590 820.000 ;
    END
  END mprj_dat_i[26]
  PIN mprj_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2522.730 816.000 2523.010 820.000 ;
    END
  END mprj_dat_i[27]
  PIN mprj_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2535.150 816.000 2535.430 820.000 ;
    END
  END mprj_dat_i[28]
  PIN mprj_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2547.570 816.000 2547.850 820.000 ;
    END
  END mprj_dat_i[29]
  PIN mprj_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2203.950 816.000 2204.230 820.000 ;
    END
  END mprj_dat_i[2]
  PIN mprj_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2559.990 816.000 2560.270 820.000 ;
    END
  END mprj_dat_i[30]
  PIN mprj_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2572.410 816.000 2572.690 820.000 ;
    END
  END mprj_dat_i[31]
  PIN mprj_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2220.510 816.000 2220.790 820.000 ;
    END
  END mprj_dat_i[3]
  PIN mprj_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2237.070 816.000 2237.350 820.000 ;
    END
  END mprj_dat_i[4]
  PIN mprj_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2249.490 816.000 2249.770 820.000 ;
    END
  END mprj_dat_i[5]
  PIN mprj_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2261.910 816.000 2262.190 820.000 ;
    END
  END mprj_dat_i[6]
  PIN mprj_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2274.330 816.000 2274.610 820.000 ;
    END
  END mprj_dat_i[7]
  PIN mprj_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2286.750 816.000 2287.030 820.000 ;
    END
  END mprj_dat_i[8]
  PIN mprj_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2299.170 816.000 2299.450 820.000 ;
    END
  END mprj_dat_i[9]
  PIN mprj_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2174.970 816.000 2175.250 820.000 ;
    END
  END mprj_dat_o[0]
  PIN mprj_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2315.730 816.000 2316.010 820.000 ;
    END
  END mprj_dat_o[10]
  PIN mprj_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.150 816.000 2328.430 820.000 ;
    END
  END mprj_dat_o[11]
  PIN mprj_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2340.570 816.000 2340.850 820.000 ;
    END
  END mprj_dat_o[12]
  PIN mprj_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2352.990 816.000 2353.270 820.000 ;
    END
  END mprj_dat_o[13]
  PIN mprj_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2365.410 816.000 2365.690 820.000 ;
    END
  END mprj_dat_o[14]
  PIN mprj_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2377.830 816.000 2378.110 820.000 ;
    END
  END mprj_dat_o[15]
  PIN mprj_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.250 816.000 2390.530 820.000 ;
    END
  END mprj_dat_o[16]
  PIN mprj_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2402.670 816.000 2402.950 820.000 ;
    END
  END mprj_dat_o[17]
  PIN mprj_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2415.090 816.000 2415.370 820.000 ;
    END
  END mprj_dat_o[18]
  PIN mprj_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2427.510 816.000 2427.790 820.000 ;
    END
  END mprj_dat_o[19]
  PIN mprj_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2191.530 816.000 2191.810 820.000 ;
    END
  END mprj_dat_o[1]
  PIN mprj_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2439.930 816.000 2440.210 820.000 ;
    END
  END mprj_dat_o[20]
  PIN mprj_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2452.350 816.000 2452.630 820.000 ;
    END
  END mprj_dat_o[21]
  PIN mprj_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2464.770 816.000 2465.050 820.000 ;
    END
  END mprj_dat_o[22]
  PIN mprj_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2477.190 816.000 2477.470 820.000 ;
    END
  END mprj_dat_o[23]
  PIN mprj_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2489.610 816.000 2489.890 820.000 ;
    END
  END mprj_dat_o[24]
  PIN mprj_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2502.030 816.000 2502.310 820.000 ;
    END
  END mprj_dat_o[25]
  PIN mprj_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2514.450 816.000 2514.730 820.000 ;
    END
  END mprj_dat_o[26]
  PIN mprj_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2526.870 816.000 2527.150 820.000 ;
    END
  END mprj_dat_o[27]
  PIN mprj_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2539.290 816.000 2539.570 820.000 ;
    END
  END mprj_dat_o[28]
  PIN mprj_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2551.710 816.000 2551.990 820.000 ;
    END
  END mprj_dat_o[29]
  PIN mprj_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2208.090 816.000 2208.370 820.000 ;
    END
  END mprj_dat_o[2]
  PIN mprj_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2564.130 816.000 2564.410 820.000 ;
    END
  END mprj_dat_o[30]
  PIN mprj_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2576.550 816.000 2576.830 820.000 ;
    END
  END mprj_dat_o[31]
  PIN mprj_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.650 816.000 2224.930 820.000 ;
    END
  END mprj_dat_o[3]
  PIN mprj_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2241.210 816.000 2241.490 820.000 ;
    END
  END mprj_dat_o[4]
  PIN mprj_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2253.630 816.000 2253.910 820.000 ;
    END
  END mprj_dat_o[5]
  PIN mprj_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2266.050 816.000 2266.330 820.000 ;
    END
  END mprj_dat_o[6]
  PIN mprj_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2278.470 816.000 2278.750 820.000 ;
    END
  END mprj_dat_o[7]
  PIN mprj_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.890 816.000 2291.170 820.000 ;
    END
  END mprj_dat_o[8]
  PIN mprj_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2303.310 816.000 2303.590 820.000 ;
    END
  END mprj_dat_o[9]
  PIN mprj_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2179.110 816.000 2179.390 820.000 ;
    END
  END mprj_sel_o[0]
  PIN mprj_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.670 816.000 2195.950 820.000 ;
    END
  END mprj_sel_o[1]
  PIN mprj_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2212.230 816.000 2212.510 820.000 ;
    END
  END mprj_sel_o[2]
  PIN mprj_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2228.790 816.000 2229.070 820.000 ;
    END
  END mprj_sel_o[3]
  PIN mprj_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.270 816.000 2154.550 820.000 ;
    END
  END mprj_stb_o
  PIN mprj_wb_iena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2158.410 816.000 2158.690 820.000 ;
    END
  END mprj_wb_iena
  PIN mprj_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2162.550 816.000 2162.830 820.000 ;
    END
  END mprj_we_o
  PIN por_l_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 66.680 2620.000 67.280 ;
    END
  END por_l_in
  PIN por_l_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.860 0.000 1280.140 4.000 ;
    END
  END por_l_out
  PIN porb_h_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 77.560 2620.000 78.160 ;
    END
  END porb_h_in
  PIN porb_h_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.860 0.000 1290.140 4.000 ;
    END
  END porb_h_out
  PIN qspi_enabled
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 273.400 2620.000 274.000 ;
    END
  END qspi_enabled
  PIN resetn_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.860 0.000 1330.140 4.000 ;
    END
  END resetn_in
  PIN resetn_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 816.000 1198.210 820.000 ;
    END
  END resetn_out
  PIN rstb_l_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.860 0.000 1270.140 4.000 ;
    END
  END rstb_l_in
  PIN rstb_l_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 12.280 2620.000 12.880 ;
    END
  END rstb_l_out
  PIN ser_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 229.880 2620.000 230.480 ;
    END
  END ser_rx
  PIN ser_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 240.760 2620.000 241.360 ;
    END
  END ser_tx
  PIN serial_clock_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 55.800 2620.000 56.400 ;
    END
  END serial_clock_in
  PIN serial_clock_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.760 4.000 717.360 ;
    END
  END serial_clock_out
  PIN serial_data_2_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 34.040 2620.000 34.640 ;
    END
  END serial_data_2_in
  PIN serial_data_2_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 696.760 4.000 697.360 ;
    END
  END serial_data_2_out
  PIN serial_load_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 23.160 2620.000 23.760 ;
    END
  END serial_load_in
  PIN serial_load_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 686.760 4.000 687.360 ;
    END
  END serial_load_out
  PIN serial_resetn_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 44.920 2620.000 45.520 ;
    END
  END serial_resetn_in
  PIN serial_resetn_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 706.760 4.000 707.360 ;
    END
  END serial_resetn_out
  PIN spi_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 208.120 2620.000 208.720 ;
    END
  END spi_csb
  PIN spi_enabled
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 251.640 2620.000 252.240 ;
    END
  END spi_enabled
  PIN spi_sck
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 197.240 2620.000 197.840 ;
    END
  END spi_sck
  PIN spi_sdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 219.000 2620.000 219.600 ;
    END
  END spi_sdi
  PIN spi_sdo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 186.360 2620.000 186.960 ;
    END
  END spi_sdo
  PIN spi_sdoenb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 175.480 2620.000 176.080 ;
    END
  END spi_sdoenb
  PIN trap
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 131.960 2620.000 132.560 ;
    END
  END trap
  PIN uart_enabled
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2616.000 262.520 2620.000 263.120 ;
    END
  END uart_enabled
  PIN user_irq_ena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2580.690 816.000 2580.970 820.000 ;
    END
  END user_irq_ena[0]
  PIN user_irq_ena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2584.830 816.000 2585.110 820.000 ;
    END
  END user_irq_ena[1]
  PIN user_irq_ena[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2588.970 816.000 2589.250 820.000 ;
    END
  END user_irq_ena[2]
  OBS
      LAYER li1 ;
        RECT 10.120 13.515 2609.580 805.205 ;
      LAYER met1 ;
        RECT 10.120 13.360 2609.580 819.700 ;
      LAYER met2 ;
        RECT 14.350 815.720 17.750 819.730 ;
        RECT 18.590 815.720 21.890 819.730 ;
        RECT 22.730 815.720 26.030 819.730 ;
        RECT 26.870 815.720 30.170 819.730 ;
        RECT 31.010 815.720 34.310 819.730 ;
        RECT 35.150 815.720 38.450 819.730 ;
        RECT 39.290 815.720 42.590 819.730 ;
        RECT 43.430 815.720 46.730 819.730 ;
        RECT 47.570 815.720 50.870 819.730 ;
        RECT 51.710 815.720 55.010 819.730 ;
        RECT 55.850 815.720 59.150 819.730 ;
        RECT 59.990 815.720 63.290 819.730 ;
        RECT 64.130 815.720 67.430 819.730 ;
        RECT 68.270 815.720 71.570 819.730 ;
        RECT 72.410 815.720 75.710 819.730 ;
        RECT 76.550 815.720 79.850 819.730 ;
        RECT 80.690 815.720 83.990 819.730 ;
        RECT 84.830 815.720 88.130 819.730 ;
        RECT 88.970 815.720 92.270 819.730 ;
        RECT 93.110 815.720 96.410 819.730 ;
        RECT 97.250 815.720 100.550 819.730 ;
        RECT 101.390 815.720 104.690 819.730 ;
        RECT 105.530 815.720 108.830 819.730 ;
        RECT 109.670 815.720 112.970 819.730 ;
        RECT 113.810 815.720 117.110 819.730 ;
        RECT 117.950 815.720 121.250 819.730 ;
        RECT 122.090 815.720 125.390 819.730 ;
        RECT 126.230 815.720 129.530 819.730 ;
        RECT 130.370 815.720 133.670 819.730 ;
        RECT 134.510 815.720 137.810 819.730 ;
        RECT 138.650 815.720 141.950 819.730 ;
        RECT 142.790 815.720 146.090 819.730 ;
        RECT 146.930 815.720 150.230 819.730 ;
        RECT 151.070 815.720 154.370 819.730 ;
        RECT 155.210 815.720 158.510 819.730 ;
        RECT 159.350 815.720 162.650 819.730 ;
        RECT 163.490 815.720 166.790 819.730 ;
        RECT 167.630 815.720 170.930 819.730 ;
        RECT 171.770 815.720 175.070 819.730 ;
        RECT 175.910 815.720 179.210 819.730 ;
        RECT 180.050 815.720 183.350 819.730 ;
        RECT 184.190 815.720 187.490 819.730 ;
        RECT 188.330 815.720 191.630 819.730 ;
        RECT 192.470 815.720 195.770 819.730 ;
        RECT 196.610 815.720 199.910 819.730 ;
        RECT 200.750 815.720 204.050 819.730 ;
        RECT 204.890 815.720 208.190 819.730 ;
        RECT 209.030 815.720 212.330 819.730 ;
        RECT 213.170 815.720 216.470 819.730 ;
        RECT 217.310 815.720 220.610 819.730 ;
        RECT 221.450 815.720 224.750 819.730 ;
        RECT 225.590 815.720 228.890 819.730 ;
        RECT 229.730 815.720 233.030 819.730 ;
        RECT 233.870 815.720 237.170 819.730 ;
        RECT 238.010 815.720 241.310 819.730 ;
        RECT 242.150 815.720 245.450 819.730 ;
        RECT 246.290 815.720 249.590 819.730 ;
        RECT 250.430 815.720 253.730 819.730 ;
        RECT 254.570 815.720 257.870 819.730 ;
        RECT 258.710 815.720 262.010 819.730 ;
        RECT 262.850 815.720 266.150 819.730 ;
        RECT 266.990 815.720 270.290 819.730 ;
        RECT 271.130 815.720 274.430 819.730 ;
        RECT 275.270 815.720 278.570 819.730 ;
        RECT 279.410 815.720 282.710 819.730 ;
        RECT 283.550 815.720 286.850 819.730 ;
        RECT 287.690 815.720 290.990 819.730 ;
        RECT 291.830 815.720 295.130 819.730 ;
        RECT 295.970 815.720 299.270 819.730 ;
        RECT 300.110 815.720 303.410 819.730 ;
        RECT 304.250 815.720 307.550 819.730 ;
        RECT 308.390 815.720 311.690 819.730 ;
        RECT 312.530 815.720 315.830 819.730 ;
        RECT 316.670 815.720 319.970 819.730 ;
        RECT 320.810 815.720 324.110 819.730 ;
        RECT 324.950 815.720 328.250 819.730 ;
        RECT 329.090 815.720 332.390 819.730 ;
        RECT 333.230 815.720 336.530 819.730 ;
        RECT 337.370 815.720 340.670 819.730 ;
        RECT 341.510 815.720 344.810 819.730 ;
        RECT 345.650 815.720 348.950 819.730 ;
        RECT 349.790 815.720 353.090 819.730 ;
        RECT 353.930 815.720 357.230 819.730 ;
        RECT 358.070 815.720 361.370 819.730 ;
        RECT 362.210 815.720 365.510 819.730 ;
        RECT 366.350 815.720 369.650 819.730 ;
        RECT 370.490 815.720 373.790 819.730 ;
        RECT 374.630 815.720 377.930 819.730 ;
        RECT 378.770 815.720 382.070 819.730 ;
        RECT 382.910 815.720 386.210 819.730 ;
        RECT 387.050 815.720 390.350 819.730 ;
        RECT 391.190 815.720 394.490 819.730 ;
        RECT 395.330 815.720 398.630 819.730 ;
        RECT 399.470 815.720 402.770 819.730 ;
        RECT 403.610 815.720 406.910 819.730 ;
        RECT 407.750 815.720 411.050 819.730 ;
        RECT 411.890 815.720 415.190 819.730 ;
        RECT 416.030 815.720 419.330 819.730 ;
        RECT 420.170 815.720 423.470 819.730 ;
        RECT 424.310 815.720 427.610 819.730 ;
        RECT 428.450 815.720 431.750 819.730 ;
        RECT 432.590 815.720 435.890 819.730 ;
        RECT 436.730 815.720 440.030 819.730 ;
        RECT 440.870 815.720 444.170 819.730 ;
        RECT 445.010 815.720 448.310 819.730 ;
        RECT 449.150 815.720 452.450 819.730 ;
        RECT 453.290 815.720 456.590 819.730 ;
        RECT 457.430 815.720 460.730 819.730 ;
        RECT 461.570 815.720 464.870 819.730 ;
        RECT 465.710 815.720 469.010 819.730 ;
        RECT 469.850 815.720 473.150 819.730 ;
        RECT 473.990 815.720 477.290 819.730 ;
        RECT 478.130 815.720 481.430 819.730 ;
        RECT 482.270 815.720 485.570 819.730 ;
        RECT 486.410 815.720 489.710 819.730 ;
        RECT 490.550 815.720 493.850 819.730 ;
        RECT 494.690 815.720 497.990 819.730 ;
        RECT 498.830 815.720 502.130 819.730 ;
        RECT 502.970 815.720 506.270 819.730 ;
        RECT 507.110 815.720 510.410 819.730 ;
        RECT 511.250 815.720 514.550 819.730 ;
        RECT 515.390 815.720 518.690 819.730 ;
        RECT 519.530 815.720 522.830 819.730 ;
        RECT 523.670 815.720 526.970 819.730 ;
        RECT 527.810 815.720 531.110 819.730 ;
        RECT 531.950 815.720 535.250 819.730 ;
        RECT 536.090 815.720 539.390 819.730 ;
        RECT 540.230 815.720 543.530 819.730 ;
        RECT 544.370 815.720 547.670 819.730 ;
        RECT 548.510 815.720 551.810 819.730 ;
        RECT 552.650 815.720 555.950 819.730 ;
        RECT 556.790 815.720 560.090 819.730 ;
        RECT 560.930 815.720 564.230 819.730 ;
        RECT 565.070 815.720 568.370 819.730 ;
        RECT 569.210 815.720 572.510 819.730 ;
        RECT 573.350 815.720 576.650 819.730 ;
        RECT 577.490 815.720 580.790 819.730 ;
        RECT 581.630 815.720 584.930 819.730 ;
        RECT 585.770 815.720 589.070 819.730 ;
        RECT 589.910 815.720 593.210 819.730 ;
        RECT 594.050 815.720 597.350 819.730 ;
        RECT 598.190 815.720 601.490 819.730 ;
        RECT 602.330 815.720 605.630 819.730 ;
        RECT 606.470 815.720 609.770 819.730 ;
        RECT 610.610 815.720 613.910 819.730 ;
        RECT 614.750 815.720 618.050 819.730 ;
        RECT 618.890 815.720 622.190 819.730 ;
        RECT 623.030 815.720 626.330 819.730 ;
        RECT 627.170 815.720 630.470 819.730 ;
        RECT 631.310 815.720 634.610 819.730 ;
        RECT 635.450 815.720 638.750 819.730 ;
        RECT 639.590 815.720 642.890 819.730 ;
        RECT 643.730 815.720 647.030 819.730 ;
        RECT 647.870 815.720 651.170 819.730 ;
        RECT 652.010 815.720 655.310 819.730 ;
        RECT 656.150 815.720 659.450 819.730 ;
        RECT 660.290 815.720 663.590 819.730 ;
        RECT 664.430 815.720 667.730 819.730 ;
        RECT 668.570 815.720 671.870 819.730 ;
        RECT 672.710 815.720 676.010 819.730 ;
        RECT 676.850 815.720 680.150 819.730 ;
        RECT 680.990 815.720 684.290 819.730 ;
        RECT 685.130 815.720 688.430 819.730 ;
        RECT 689.270 815.720 692.570 819.730 ;
        RECT 693.410 815.720 696.710 819.730 ;
        RECT 697.550 815.720 700.850 819.730 ;
        RECT 701.690 815.720 704.990 819.730 ;
        RECT 705.830 815.720 709.130 819.730 ;
        RECT 709.970 815.720 713.270 819.730 ;
        RECT 714.110 815.720 717.410 819.730 ;
        RECT 718.250 815.720 721.550 819.730 ;
        RECT 722.390 815.720 725.690 819.730 ;
        RECT 726.530 815.720 729.830 819.730 ;
        RECT 730.670 815.720 733.970 819.730 ;
        RECT 734.810 815.720 738.110 819.730 ;
        RECT 738.950 815.720 742.250 819.730 ;
        RECT 743.090 815.720 746.390 819.730 ;
        RECT 747.230 815.720 750.530 819.730 ;
        RECT 751.370 815.720 754.670 819.730 ;
        RECT 755.510 815.720 758.810 819.730 ;
        RECT 759.650 815.720 762.950 819.730 ;
        RECT 763.790 815.720 767.090 819.730 ;
        RECT 767.930 815.720 771.230 819.730 ;
        RECT 772.070 815.720 775.370 819.730 ;
        RECT 776.210 815.720 779.510 819.730 ;
        RECT 780.350 815.720 783.650 819.730 ;
        RECT 784.490 815.720 787.790 819.730 ;
        RECT 788.630 815.720 791.930 819.730 ;
        RECT 792.770 815.720 796.070 819.730 ;
        RECT 796.910 815.720 800.210 819.730 ;
        RECT 801.050 815.720 804.350 819.730 ;
        RECT 805.190 815.720 808.490 819.730 ;
        RECT 809.330 815.720 812.630 819.730 ;
        RECT 813.470 815.720 816.770 819.730 ;
        RECT 817.610 815.720 820.910 819.730 ;
        RECT 821.750 815.720 825.050 819.730 ;
        RECT 825.890 815.720 829.190 819.730 ;
        RECT 830.030 815.720 833.330 819.730 ;
        RECT 834.170 815.720 837.470 819.730 ;
        RECT 838.310 815.720 841.610 819.730 ;
        RECT 842.450 815.720 845.750 819.730 ;
        RECT 846.590 815.720 849.890 819.730 ;
        RECT 850.730 815.720 854.030 819.730 ;
        RECT 854.870 815.720 858.170 819.730 ;
        RECT 859.010 815.720 862.310 819.730 ;
        RECT 863.150 815.720 866.450 819.730 ;
        RECT 867.290 815.720 870.590 819.730 ;
        RECT 871.430 815.720 874.730 819.730 ;
        RECT 875.570 815.720 878.870 819.730 ;
        RECT 879.710 815.720 883.010 819.730 ;
        RECT 883.850 815.720 887.150 819.730 ;
        RECT 887.990 815.720 891.290 819.730 ;
        RECT 892.130 815.720 895.430 819.730 ;
        RECT 896.270 815.720 899.570 819.730 ;
        RECT 900.410 815.720 903.710 819.730 ;
        RECT 904.550 815.720 907.850 819.730 ;
        RECT 908.690 815.720 911.990 819.730 ;
        RECT 912.830 815.720 916.130 819.730 ;
        RECT 916.970 815.720 920.270 819.730 ;
        RECT 921.110 815.720 924.410 819.730 ;
        RECT 925.250 815.720 928.550 819.730 ;
        RECT 929.390 815.720 932.690 819.730 ;
        RECT 933.530 815.720 936.830 819.730 ;
        RECT 937.670 815.720 940.970 819.730 ;
        RECT 941.810 815.720 945.110 819.730 ;
        RECT 945.950 815.720 949.250 819.730 ;
        RECT 950.090 815.720 953.390 819.730 ;
        RECT 954.230 815.720 957.530 819.730 ;
        RECT 958.370 815.720 961.670 819.730 ;
        RECT 962.510 815.720 965.810 819.730 ;
        RECT 966.650 815.720 969.950 819.730 ;
        RECT 970.790 815.720 974.090 819.730 ;
        RECT 974.930 815.720 978.230 819.730 ;
        RECT 979.070 815.720 982.370 819.730 ;
        RECT 983.210 815.720 986.510 819.730 ;
        RECT 987.350 815.720 990.650 819.730 ;
        RECT 991.490 815.720 994.790 819.730 ;
        RECT 995.630 815.720 998.930 819.730 ;
        RECT 999.770 815.720 1003.070 819.730 ;
        RECT 1003.910 815.720 1007.210 819.730 ;
        RECT 1008.050 815.720 1011.350 819.730 ;
        RECT 1012.190 815.720 1015.490 819.730 ;
        RECT 1016.330 815.720 1019.630 819.730 ;
        RECT 1020.470 815.720 1023.770 819.730 ;
        RECT 1024.610 815.720 1027.910 819.730 ;
        RECT 1028.750 815.720 1032.050 819.730 ;
        RECT 1032.890 815.720 1036.190 819.730 ;
        RECT 1037.030 815.720 1040.330 819.730 ;
        RECT 1041.170 815.720 1044.470 819.730 ;
        RECT 1045.310 815.720 1048.610 819.730 ;
        RECT 1049.450 815.720 1052.750 819.730 ;
        RECT 1053.590 815.720 1056.890 819.730 ;
        RECT 1057.730 815.720 1061.030 819.730 ;
        RECT 1061.870 815.720 1065.170 819.730 ;
        RECT 1066.010 815.720 1069.310 819.730 ;
        RECT 1070.150 815.720 1073.450 819.730 ;
        RECT 1074.290 815.720 1077.590 819.730 ;
        RECT 1078.430 815.720 1081.730 819.730 ;
        RECT 1082.570 815.720 1085.870 819.730 ;
        RECT 1086.710 815.720 1090.010 819.730 ;
        RECT 1090.850 815.720 1094.150 819.730 ;
        RECT 1094.990 815.720 1098.290 819.730 ;
        RECT 1099.130 815.720 1102.430 819.730 ;
        RECT 1103.270 815.720 1106.570 819.730 ;
        RECT 1107.410 815.720 1110.710 819.730 ;
        RECT 1111.550 815.720 1114.850 819.730 ;
        RECT 1115.690 815.720 1118.990 819.730 ;
        RECT 1119.830 815.720 1123.130 819.730 ;
        RECT 1123.970 815.720 1127.270 819.730 ;
        RECT 1128.110 815.720 1131.410 819.730 ;
        RECT 1132.250 815.720 1135.550 819.730 ;
        RECT 1136.390 815.720 1139.690 819.730 ;
        RECT 1140.530 815.720 1143.830 819.730 ;
        RECT 1144.670 815.720 1147.970 819.730 ;
        RECT 1148.810 815.720 1152.110 819.730 ;
        RECT 1152.950 815.720 1156.250 819.730 ;
        RECT 1157.090 815.720 1160.390 819.730 ;
        RECT 1161.230 815.720 1164.530 819.730 ;
        RECT 1165.370 815.720 1168.670 819.730 ;
        RECT 1169.510 815.720 1172.810 819.730 ;
        RECT 1173.650 815.720 1176.950 819.730 ;
        RECT 1177.790 815.720 1181.090 819.730 ;
        RECT 1181.930 815.720 1185.230 819.730 ;
        RECT 1186.070 815.720 1189.370 819.730 ;
        RECT 1190.210 815.720 1193.510 819.730 ;
        RECT 1194.350 815.720 1197.650 819.730 ;
        RECT 1198.490 815.720 1201.790 819.730 ;
        RECT 1202.630 815.720 1205.930 819.730 ;
        RECT 1206.770 815.720 1210.070 819.730 ;
        RECT 1210.910 815.720 1214.210 819.730 ;
        RECT 1215.050 815.720 1218.350 819.730 ;
        RECT 1219.190 815.720 1222.490 819.730 ;
        RECT 1223.330 815.720 1226.630 819.730 ;
        RECT 1227.470 815.720 1230.770 819.730 ;
        RECT 1231.610 815.720 1234.910 819.730 ;
        RECT 1235.750 815.720 1239.050 819.730 ;
        RECT 1239.890 815.720 1243.190 819.730 ;
        RECT 1244.030 815.720 1247.330 819.730 ;
        RECT 1248.170 815.720 1251.470 819.730 ;
        RECT 1252.310 815.720 1255.610 819.730 ;
        RECT 1256.450 815.720 1259.750 819.730 ;
        RECT 1260.590 815.720 1263.890 819.730 ;
        RECT 1264.730 815.720 1268.030 819.730 ;
        RECT 1268.870 815.720 1272.170 819.730 ;
        RECT 1273.010 815.720 1276.310 819.730 ;
        RECT 1277.150 815.720 1280.450 819.730 ;
        RECT 1281.290 815.720 1284.590 819.730 ;
        RECT 1285.430 815.720 1288.730 819.730 ;
        RECT 1289.570 815.720 1292.870 819.730 ;
        RECT 1293.710 815.720 1297.010 819.730 ;
        RECT 1297.850 815.720 1301.150 819.730 ;
        RECT 1301.990 815.720 1305.290 819.730 ;
        RECT 1306.130 815.720 1309.430 819.730 ;
        RECT 1310.270 815.720 1313.570 819.730 ;
        RECT 1314.410 815.720 1317.710 819.730 ;
        RECT 1318.550 815.720 1321.850 819.730 ;
        RECT 1322.690 815.720 1325.990 819.730 ;
        RECT 1326.830 815.720 1330.130 819.730 ;
        RECT 1330.970 815.720 1334.270 819.730 ;
        RECT 1335.110 815.720 1338.410 819.730 ;
        RECT 1339.250 815.720 1342.550 819.730 ;
        RECT 1343.390 815.720 1346.690 819.730 ;
        RECT 1347.530 815.720 1350.830 819.730 ;
        RECT 1351.670 815.720 1354.970 819.730 ;
        RECT 1355.810 815.720 1359.110 819.730 ;
        RECT 1359.950 815.720 1363.250 819.730 ;
        RECT 1364.090 815.720 1367.390 819.730 ;
        RECT 1368.230 815.720 1371.530 819.730 ;
        RECT 1372.370 815.720 1375.670 819.730 ;
        RECT 1376.510 815.720 1379.810 819.730 ;
        RECT 1380.650 815.720 1383.950 819.730 ;
        RECT 1384.790 815.720 1388.090 819.730 ;
        RECT 1388.930 815.720 1392.230 819.730 ;
        RECT 1393.070 815.720 1396.370 819.730 ;
        RECT 1397.210 815.720 1400.510 819.730 ;
        RECT 1401.350 815.720 1404.650 819.730 ;
        RECT 1405.490 815.720 1408.790 819.730 ;
        RECT 1409.630 815.720 1412.930 819.730 ;
        RECT 1413.770 815.720 1417.070 819.730 ;
        RECT 1417.910 815.720 1421.210 819.730 ;
        RECT 1422.050 815.720 1425.350 819.730 ;
        RECT 1426.190 815.720 1429.490 819.730 ;
        RECT 1430.330 815.720 1433.630 819.730 ;
        RECT 1434.470 815.720 1437.770 819.730 ;
        RECT 1438.610 815.720 1441.910 819.730 ;
        RECT 1442.750 815.720 1446.050 819.730 ;
        RECT 1446.890 815.720 1450.190 819.730 ;
        RECT 1451.030 815.720 1454.330 819.730 ;
        RECT 1455.170 815.720 1458.470 819.730 ;
        RECT 1459.310 815.720 1462.610 819.730 ;
        RECT 1463.450 815.720 1466.750 819.730 ;
        RECT 1467.590 815.720 1470.890 819.730 ;
        RECT 1471.730 815.720 1475.030 819.730 ;
        RECT 1475.870 815.720 1479.170 819.730 ;
        RECT 1480.010 815.720 1483.310 819.730 ;
        RECT 1484.150 815.720 1487.450 819.730 ;
        RECT 1488.290 815.720 1491.590 819.730 ;
        RECT 1492.430 815.720 1495.730 819.730 ;
        RECT 1496.570 815.720 1499.870 819.730 ;
        RECT 1500.710 815.720 1504.010 819.730 ;
        RECT 1504.850 815.720 1508.150 819.730 ;
        RECT 1508.990 815.720 1512.290 819.730 ;
        RECT 1513.130 815.720 1516.430 819.730 ;
        RECT 1517.270 815.720 1520.570 819.730 ;
        RECT 1521.410 815.720 1524.710 819.730 ;
        RECT 1525.550 815.720 1528.850 819.730 ;
        RECT 1529.690 815.720 1532.990 819.730 ;
        RECT 1533.830 815.720 1537.130 819.730 ;
        RECT 1537.970 815.720 1541.270 819.730 ;
        RECT 1542.110 815.720 1545.410 819.730 ;
        RECT 1546.250 815.720 1549.550 819.730 ;
        RECT 1550.390 815.720 1553.690 819.730 ;
        RECT 1554.530 815.720 1557.830 819.730 ;
        RECT 1558.670 815.720 1561.970 819.730 ;
        RECT 1562.810 815.720 1566.110 819.730 ;
        RECT 1566.950 815.720 1570.250 819.730 ;
        RECT 1571.090 815.720 1574.390 819.730 ;
        RECT 1575.230 815.720 1578.530 819.730 ;
        RECT 1579.370 815.720 1582.670 819.730 ;
        RECT 1583.510 815.720 1586.810 819.730 ;
        RECT 1587.650 815.720 1590.950 819.730 ;
        RECT 1591.790 815.720 1595.090 819.730 ;
        RECT 1595.930 815.720 1599.230 819.730 ;
        RECT 1600.070 815.720 1603.370 819.730 ;
        RECT 1604.210 815.720 1607.510 819.730 ;
        RECT 1608.350 815.720 1611.650 819.730 ;
        RECT 1612.490 815.720 1615.790 819.730 ;
        RECT 1616.630 815.720 1619.930 819.730 ;
        RECT 1620.770 815.720 1624.070 819.730 ;
        RECT 1624.910 815.720 1628.210 819.730 ;
        RECT 1629.050 815.720 1632.350 819.730 ;
        RECT 1633.190 815.720 1636.490 819.730 ;
        RECT 1637.330 815.720 1640.630 819.730 ;
        RECT 1641.470 815.720 1644.770 819.730 ;
        RECT 1645.610 815.720 1648.910 819.730 ;
        RECT 1649.750 815.720 1653.050 819.730 ;
        RECT 1653.890 815.720 1657.190 819.730 ;
        RECT 1658.030 815.720 1661.330 819.730 ;
        RECT 1662.170 815.720 1665.470 819.730 ;
        RECT 1666.310 815.720 1669.610 819.730 ;
        RECT 1670.450 815.720 1673.750 819.730 ;
        RECT 1674.590 815.720 1677.890 819.730 ;
        RECT 1678.730 815.720 1682.030 819.730 ;
        RECT 1682.870 815.720 1686.170 819.730 ;
        RECT 1687.010 815.720 1690.310 819.730 ;
        RECT 1691.150 815.720 1694.450 819.730 ;
        RECT 1695.290 815.720 1698.590 819.730 ;
        RECT 1699.430 815.720 1702.730 819.730 ;
        RECT 1703.570 815.720 1706.870 819.730 ;
        RECT 1707.710 815.720 1711.010 819.730 ;
        RECT 1711.850 815.720 1715.150 819.730 ;
        RECT 1715.990 815.720 1719.290 819.730 ;
        RECT 1720.130 815.720 1723.430 819.730 ;
        RECT 1724.270 815.720 1727.570 819.730 ;
        RECT 1728.410 815.720 1731.710 819.730 ;
        RECT 1732.550 815.720 1735.850 819.730 ;
        RECT 1736.690 815.720 1739.990 819.730 ;
        RECT 1740.830 815.720 1744.130 819.730 ;
        RECT 1744.970 815.720 1748.270 819.730 ;
        RECT 1749.110 815.720 1752.410 819.730 ;
        RECT 1753.250 815.720 1756.550 819.730 ;
        RECT 1757.390 815.720 1760.690 819.730 ;
        RECT 1761.530 815.720 1764.830 819.730 ;
        RECT 1765.670 815.720 1768.970 819.730 ;
        RECT 1769.810 815.720 1773.110 819.730 ;
        RECT 1773.950 815.720 1777.250 819.730 ;
        RECT 1778.090 815.720 1781.390 819.730 ;
        RECT 1782.230 815.720 1785.530 819.730 ;
        RECT 1786.370 815.720 1789.670 819.730 ;
        RECT 1790.510 815.720 1793.810 819.730 ;
        RECT 1794.650 815.720 1797.950 819.730 ;
        RECT 1798.790 815.720 1802.090 819.730 ;
        RECT 1802.930 815.720 1806.230 819.730 ;
        RECT 1807.070 815.720 1810.370 819.730 ;
        RECT 1811.210 815.720 1814.510 819.730 ;
        RECT 1815.350 815.720 1818.650 819.730 ;
        RECT 1819.490 815.720 1822.790 819.730 ;
        RECT 1823.630 815.720 1826.930 819.730 ;
        RECT 1827.770 815.720 1831.070 819.730 ;
        RECT 1831.910 815.720 1835.210 819.730 ;
        RECT 1836.050 815.720 1839.350 819.730 ;
        RECT 1840.190 815.720 1843.490 819.730 ;
        RECT 1844.330 815.720 1847.630 819.730 ;
        RECT 1848.470 815.720 1851.770 819.730 ;
        RECT 1852.610 815.720 1855.910 819.730 ;
        RECT 1856.750 815.720 1860.050 819.730 ;
        RECT 1860.890 815.720 1864.190 819.730 ;
        RECT 1865.030 815.720 1868.330 819.730 ;
        RECT 1869.170 815.720 1872.470 819.730 ;
        RECT 1873.310 815.720 1876.610 819.730 ;
        RECT 1877.450 815.720 1880.750 819.730 ;
        RECT 1881.590 815.720 1884.890 819.730 ;
        RECT 1885.730 815.720 1889.030 819.730 ;
        RECT 1889.870 815.720 1893.170 819.730 ;
        RECT 1894.010 815.720 1897.310 819.730 ;
        RECT 1898.150 815.720 1901.450 819.730 ;
        RECT 1902.290 815.720 1905.590 819.730 ;
        RECT 1906.430 815.720 1909.730 819.730 ;
        RECT 1910.570 815.720 1913.870 819.730 ;
        RECT 1914.710 815.720 1918.010 819.730 ;
        RECT 1918.850 815.720 1922.150 819.730 ;
        RECT 1922.990 815.720 1926.290 819.730 ;
        RECT 1927.130 815.720 1930.430 819.730 ;
        RECT 1931.270 815.720 1934.570 819.730 ;
        RECT 1935.410 815.720 1938.710 819.730 ;
        RECT 1939.550 815.720 1942.850 819.730 ;
        RECT 1943.690 815.720 1946.990 819.730 ;
        RECT 1947.830 815.720 1951.130 819.730 ;
        RECT 1951.970 815.720 1955.270 819.730 ;
        RECT 1956.110 815.720 1959.410 819.730 ;
        RECT 1960.250 815.720 1963.550 819.730 ;
        RECT 1964.390 815.720 1967.690 819.730 ;
        RECT 1968.530 815.720 1971.830 819.730 ;
        RECT 1972.670 815.720 1975.970 819.730 ;
        RECT 1976.810 815.720 1980.110 819.730 ;
        RECT 1980.950 815.720 1984.250 819.730 ;
        RECT 1985.090 815.720 1988.390 819.730 ;
        RECT 1989.230 815.720 1992.530 819.730 ;
        RECT 1993.370 815.720 1996.670 819.730 ;
        RECT 1997.510 815.720 2000.810 819.730 ;
        RECT 2001.650 815.720 2004.950 819.730 ;
        RECT 2005.790 815.720 2009.090 819.730 ;
        RECT 2009.930 815.720 2013.230 819.730 ;
        RECT 2014.070 815.720 2017.370 819.730 ;
        RECT 2018.210 815.720 2021.510 819.730 ;
        RECT 2022.350 815.720 2025.650 819.730 ;
        RECT 2026.490 815.720 2029.790 819.730 ;
        RECT 2030.630 815.720 2033.930 819.730 ;
        RECT 2034.770 815.720 2038.070 819.730 ;
        RECT 2038.910 815.720 2042.210 819.730 ;
        RECT 2043.050 815.720 2046.350 819.730 ;
        RECT 2047.190 815.720 2050.490 819.730 ;
        RECT 2051.330 815.720 2054.630 819.730 ;
        RECT 2055.470 815.720 2058.770 819.730 ;
        RECT 2059.610 815.720 2062.910 819.730 ;
        RECT 2063.750 815.720 2067.050 819.730 ;
        RECT 2067.890 815.720 2071.190 819.730 ;
        RECT 2072.030 815.720 2075.330 819.730 ;
        RECT 2076.170 815.720 2079.470 819.730 ;
        RECT 2080.310 815.720 2083.610 819.730 ;
        RECT 2084.450 815.720 2087.750 819.730 ;
        RECT 2088.590 815.720 2091.890 819.730 ;
        RECT 2092.730 815.720 2096.030 819.730 ;
        RECT 2096.870 815.720 2100.170 819.730 ;
        RECT 2101.010 815.720 2104.310 819.730 ;
        RECT 2105.150 815.720 2108.450 819.730 ;
        RECT 2109.290 815.720 2112.590 819.730 ;
        RECT 2113.430 815.720 2116.730 819.730 ;
        RECT 2117.570 815.720 2120.870 819.730 ;
        RECT 2121.710 815.720 2125.010 819.730 ;
        RECT 2125.850 815.720 2129.150 819.730 ;
        RECT 2129.990 815.720 2133.290 819.730 ;
        RECT 2134.130 815.720 2137.430 819.730 ;
        RECT 2138.270 815.720 2141.570 819.730 ;
        RECT 2142.410 815.720 2145.710 819.730 ;
        RECT 2146.550 815.720 2149.850 819.730 ;
        RECT 2150.690 815.720 2153.990 819.730 ;
        RECT 2154.830 815.720 2158.130 819.730 ;
        RECT 2158.970 815.720 2162.270 819.730 ;
        RECT 2163.110 815.720 2166.410 819.730 ;
        RECT 2167.250 815.720 2170.550 819.730 ;
        RECT 2171.390 815.720 2174.690 819.730 ;
        RECT 2175.530 815.720 2178.830 819.730 ;
        RECT 2179.670 815.720 2182.970 819.730 ;
        RECT 2183.810 815.720 2187.110 819.730 ;
        RECT 2187.950 815.720 2191.250 819.730 ;
        RECT 2192.090 815.720 2195.390 819.730 ;
        RECT 2196.230 815.720 2199.530 819.730 ;
        RECT 2200.370 815.720 2203.670 819.730 ;
        RECT 2204.510 815.720 2207.810 819.730 ;
        RECT 2208.650 815.720 2211.950 819.730 ;
        RECT 2212.790 815.720 2216.090 819.730 ;
        RECT 2216.930 815.720 2220.230 819.730 ;
        RECT 2221.070 815.720 2224.370 819.730 ;
        RECT 2225.210 815.720 2228.510 819.730 ;
        RECT 2229.350 815.720 2232.650 819.730 ;
        RECT 2233.490 815.720 2236.790 819.730 ;
        RECT 2237.630 815.720 2240.930 819.730 ;
        RECT 2241.770 815.720 2245.070 819.730 ;
        RECT 2245.910 815.720 2249.210 819.730 ;
        RECT 2250.050 815.720 2253.350 819.730 ;
        RECT 2254.190 815.720 2257.490 819.730 ;
        RECT 2258.330 815.720 2261.630 819.730 ;
        RECT 2262.470 815.720 2265.770 819.730 ;
        RECT 2266.610 815.720 2269.910 819.730 ;
        RECT 2270.750 815.720 2274.050 819.730 ;
        RECT 2274.890 815.720 2278.190 819.730 ;
        RECT 2279.030 815.720 2282.330 819.730 ;
        RECT 2283.170 815.720 2286.470 819.730 ;
        RECT 2287.310 815.720 2290.610 819.730 ;
        RECT 2291.450 815.720 2294.750 819.730 ;
        RECT 2295.590 815.720 2298.890 819.730 ;
        RECT 2299.730 815.720 2303.030 819.730 ;
        RECT 2303.870 815.720 2307.170 819.730 ;
        RECT 2308.010 815.720 2311.310 819.730 ;
        RECT 2312.150 815.720 2315.450 819.730 ;
        RECT 2316.290 815.720 2319.590 819.730 ;
        RECT 2320.430 815.720 2323.730 819.730 ;
        RECT 2324.570 815.720 2327.870 819.730 ;
        RECT 2328.710 815.720 2332.010 819.730 ;
        RECT 2332.850 815.720 2336.150 819.730 ;
        RECT 2336.990 815.720 2340.290 819.730 ;
        RECT 2341.130 815.720 2344.430 819.730 ;
        RECT 2345.270 815.720 2348.570 819.730 ;
        RECT 2349.410 815.720 2352.710 819.730 ;
        RECT 2353.550 815.720 2356.850 819.730 ;
        RECT 2357.690 815.720 2360.990 819.730 ;
        RECT 2361.830 815.720 2365.130 819.730 ;
        RECT 2365.970 815.720 2369.270 819.730 ;
        RECT 2370.110 815.720 2373.410 819.730 ;
        RECT 2374.250 815.720 2377.550 819.730 ;
        RECT 2378.390 815.720 2381.690 819.730 ;
        RECT 2382.530 815.720 2385.830 819.730 ;
        RECT 2386.670 815.720 2389.970 819.730 ;
        RECT 2390.810 815.720 2394.110 819.730 ;
        RECT 2394.950 815.720 2398.250 819.730 ;
        RECT 2399.090 815.720 2402.390 819.730 ;
        RECT 2403.230 815.720 2406.530 819.730 ;
        RECT 2407.370 815.720 2410.670 819.730 ;
        RECT 2411.510 815.720 2414.810 819.730 ;
        RECT 2415.650 815.720 2418.950 819.730 ;
        RECT 2419.790 815.720 2423.090 819.730 ;
        RECT 2423.930 815.720 2427.230 819.730 ;
        RECT 2428.070 815.720 2431.370 819.730 ;
        RECT 2432.210 815.720 2435.510 819.730 ;
        RECT 2436.350 815.720 2439.650 819.730 ;
        RECT 2440.490 815.720 2443.790 819.730 ;
        RECT 2444.630 815.720 2447.930 819.730 ;
        RECT 2448.770 815.720 2452.070 819.730 ;
        RECT 2452.910 815.720 2456.210 819.730 ;
        RECT 2457.050 815.720 2460.350 819.730 ;
        RECT 2461.190 815.720 2464.490 819.730 ;
        RECT 2465.330 815.720 2468.630 819.730 ;
        RECT 2469.470 815.720 2472.770 819.730 ;
        RECT 2473.610 815.720 2476.910 819.730 ;
        RECT 2477.750 815.720 2481.050 819.730 ;
        RECT 2481.890 815.720 2485.190 819.730 ;
        RECT 2486.030 815.720 2489.330 819.730 ;
        RECT 2490.170 815.720 2493.470 819.730 ;
        RECT 2494.310 815.720 2497.610 819.730 ;
        RECT 2498.450 815.720 2501.750 819.730 ;
        RECT 2502.590 815.720 2505.890 819.730 ;
        RECT 2506.730 815.720 2510.030 819.730 ;
        RECT 2510.870 815.720 2514.170 819.730 ;
        RECT 2515.010 815.720 2518.310 819.730 ;
        RECT 2519.150 815.720 2522.450 819.730 ;
        RECT 2523.290 815.720 2526.590 819.730 ;
        RECT 2527.430 815.720 2530.730 819.730 ;
        RECT 2531.570 815.720 2534.870 819.730 ;
        RECT 2535.710 815.720 2539.010 819.730 ;
        RECT 2539.850 815.720 2543.150 819.730 ;
        RECT 2543.990 815.720 2547.290 819.730 ;
        RECT 2548.130 815.720 2551.430 819.730 ;
        RECT 2552.270 815.720 2555.570 819.730 ;
        RECT 2556.410 815.720 2559.710 819.730 ;
        RECT 2560.550 815.720 2563.850 819.730 ;
        RECT 2564.690 815.720 2567.990 819.730 ;
        RECT 2568.830 815.720 2572.130 819.730 ;
        RECT 2572.970 815.720 2576.270 819.730 ;
        RECT 2577.110 815.720 2580.410 819.730 ;
        RECT 2581.250 815.720 2584.550 819.730 ;
        RECT 2585.390 815.720 2588.690 819.730 ;
        RECT 2589.530 815.720 2592.830 819.730 ;
        RECT 2593.670 815.720 2596.970 819.730 ;
        RECT 2597.810 815.720 2601.110 819.730 ;
        RECT 2601.950 815.720 2609.480 819.730 ;
        RECT 14.350 4.280 2609.480 815.720 ;
        RECT 14.350 3.740 1269.580 4.280 ;
        RECT 1270.420 3.740 1279.580 4.280 ;
        RECT 1280.420 3.740 1289.580 4.280 ;
        RECT 1290.420 3.740 1299.580 4.280 ;
        RECT 1300.420 3.740 1309.580 4.280 ;
        RECT 1310.420 3.740 1319.580 4.280 ;
        RECT 1320.420 3.740 1329.580 4.280 ;
        RECT 1330.420 3.740 2459.580 4.280 ;
        RECT 2460.420 3.740 2469.580 4.280 ;
        RECT 2470.420 3.740 2479.580 4.280 ;
        RECT 2480.420 3.740 2489.580 4.280 ;
        RECT 2490.420 3.740 2499.580 4.280 ;
        RECT 2500.420 3.740 2509.580 4.280 ;
        RECT 2510.420 3.740 2609.480 4.280 ;
      LAYER met3 ;
        RECT 3.220 807.520 2616.000 809.705 ;
        RECT 3.220 806.120 2615.600 807.520 ;
        RECT 3.220 796.640 2616.000 806.120 ;
        RECT 3.220 795.240 2615.600 796.640 ;
        RECT 3.220 785.760 2616.000 795.240 ;
        RECT 3.220 784.360 2615.600 785.760 ;
        RECT 3.220 774.880 2616.000 784.360 ;
        RECT 3.220 773.480 2615.600 774.880 ;
        RECT 3.220 764.000 2616.000 773.480 ;
        RECT 3.220 762.600 2615.600 764.000 ;
        RECT 3.220 753.120 2616.000 762.600 ;
        RECT 3.220 751.720 2615.600 753.120 ;
        RECT 3.220 742.240 2616.000 751.720 ;
        RECT 3.220 740.840 2615.600 742.240 ;
        RECT 3.220 731.360 2616.000 740.840 ;
        RECT 3.220 729.960 2615.600 731.360 ;
        RECT 3.220 720.480 2616.000 729.960 ;
        RECT 3.220 719.080 2615.600 720.480 ;
        RECT 3.220 717.760 2616.000 719.080 ;
        RECT 4.400 716.360 2616.000 717.760 ;
        RECT 3.220 709.600 2616.000 716.360 ;
        RECT 3.220 708.200 2615.600 709.600 ;
        RECT 3.220 707.760 2616.000 708.200 ;
        RECT 4.400 706.360 2616.000 707.760 ;
        RECT 3.220 698.720 2616.000 706.360 ;
        RECT 3.220 697.760 2615.600 698.720 ;
        RECT 4.400 697.320 2615.600 697.760 ;
        RECT 4.400 696.360 2616.000 697.320 ;
        RECT 3.220 687.840 2616.000 696.360 ;
        RECT 3.220 687.760 2615.600 687.840 ;
        RECT 4.400 686.440 2615.600 687.760 ;
        RECT 4.400 686.360 2616.000 686.440 ;
        RECT 3.220 676.960 2616.000 686.360 ;
        RECT 3.220 675.560 2615.600 676.960 ;
        RECT 3.220 666.080 2616.000 675.560 ;
        RECT 3.220 664.680 2615.600 666.080 ;
        RECT 3.220 655.200 2616.000 664.680 ;
        RECT 3.220 653.800 2615.600 655.200 ;
        RECT 3.220 644.320 2616.000 653.800 ;
        RECT 3.220 642.920 2615.600 644.320 ;
        RECT 3.220 633.440 2616.000 642.920 ;
        RECT 3.220 632.040 2615.600 633.440 ;
        RECT 3.220 622.560 2616.000 632.040 ;
        RECT 3.220 621.160 2615.600 622.560 ;
        RECT 3.220 611.680 2616.000 621.160 ;
        RECT 3.220 610.280 2615.600 611.680 ;
        RECT 3.220 600.800 2616.000 610.280 ;
        RECT 3.220 599.400 2615.600 600.800 ;
        RECT 3.220 589.920 2616.000 599.400 ;
        RECT 3.220 588.520 2615.600 589.920 ;
        RECT 3.220 579.040 2616.000 588.520 ;
        RECT 3.220 577.640 2615.600 579.040 ;
        RECT 3.220 568.160 2616.000 577.640 ;
        RECT 3.220 566.760 2615.600 568.160 ;
        RECT 3.220 557.280 2616.000 566.760 ;
        RECT 3.220 555.880 2615.600 557.280 ;
        RECT 3.220 546.400 2616.000 555.880 ;
        RECT 3.220 545.000 2615.600 546.400 ;
        RECT 3.220 535.520 2616.000 545.000 ;
        RECT 3.220 534.120 2615.600 535.520 ;
        RECT 3.220 524.640 2616.000 534.120 ;
        RECT 3.220 523.240 2615.600 524.640 ;
        RECT 3.220 513.760 2616.000 523.240 ;
        RECT 3.220 512.360 2615.600 513.760 ;
        RECT 3.220 502.880 2616.000 512.360 ;
        RECT 3.220 501.480 2615.600 502.880 ;
        RECT 3.220 492.000 2616.000 501.480 ;
        RECT 3.220 490.600 2615.600 492.000 ;
        RECT 3.220 481.120 2616.000 490.600 ;
        RECT 3.220 479.720 2615.600 481.120 ;
        RECT 3.220 470.240 2616.000 479.720 ;
        RECT 3.220 468.840 2615.600 470.240 ;
        RECT 3.220 459.360 2616.000 468.840 ;
        RECT 3.220 457.960 2615.600 459.360 ;
        RECT 3.220 448.480 2616.000 457.960 ;
        RECT 3.220 447.080 2615.600 448.480 ;
        RECT 3.220 437.600 2616.000 447.080 ;
        RECT 3.220 436.200 2615.600 437.600 ;
        RECT 3.220 426.720 2616.000 436.200 ;
        RECT 3.220 425.320 2615.600 426.720 ;
        RECT 3.220 415.840 2616.000 425.320 ;
        RECT 3.220 414.440 2615.600 415.840 ;
        RECT 3.220 404.960 2616.000 414.440 ;
        RECT 3.220 403.560 2615.600 404.960 ;
        RECT 3.220 394.080 2616.000 403.560 ;
        RECT 3.220 392.680 2615.600 394.080 ;
        RECT 3.220 383.200 2616.000 392.680 ;
        RECT 3.220 381.800 2615.600 383.200 ;
        RECT 3.220 372.320 2616.000 381.800 ;
        RECT 3.220 370.920 2615.600 372.320 ;
        RECT 3.220 361.440 2616.000 370.920 ;
        RECT 3.220 360.040 2615.600 361.440 ;
        RECT 3.220 350.560 2616.000 360.040 ;
        RECT 3.220 349.160 2615.600 350.560 ;
        RECT 3.220 339.680 2616.000 349.160 ;
        RECT 3.220 338.280 2615.600 339.680 ;
        RECT 3.220 328.800 2616.000 338.280 ;
        RECT 3.220 327.400 2615.600 328.800 ;
        RECT 3.220 317.920 2616.000 327.400 ;
        RECT 3.220 316.520 2615.600 317.920 ;
        RECT 3.220 307.040 2616.000 316.520 ;
        RECT 3.220 305.640 2615.600 307.040 ;
        RECT 3.220 296.160 2616.000 305.640 ;
        RECT 3.220 294.760 2615.600 296.160 ;
        RECT 3.220 285.280 2616.000 294.760 ;
        RECT 3.220 283.880 2615.600 285.280 ;
        RECT 3.220 274.400 2616.000 283.880 ;
        RECT 3.220 273.000 2615.600 274.400 ;
        RECT 3.220 263.520 2616.000 273.000 ;
        RECT 3.220 262.120 2615.600 263.520 ;
        RECT 3.220 252.640 2616.000 262.120 ;
        RECT 3.220 251.240 2615.600 252.640 ;
        RECT 3.220 241.760 2616.000 251.240 ;
        RECT 3.220 240.360 2615.600 241.760 ;
        RECT 3.220 230.880 2616.000 240.360 ;
        RECT 3.220 229.480 2615.600 230.880 ;
        RECT 3.220 220.000 2616.000 229.480 ;
        RECT 3.220 218.600 2615.600 220.000 ;
        RECT 3.220 209.120 2616.000 218.600 ;
        RECT 3.220 207.720 2615.600 209.120 ;
        RECT 3.220 198.240 2616.000 207.720 ;
        RECT 3.220 196.840 2615.600 198.240 ;
        RECT 3.220 187.360 2616.000 196.840 ;
        RECT 3.220 185.960 2615.600 187.360 ;
        RECT 3.220 176.480 2616.000 185.960 ;
        RECT 3.220 175.080 2615.600 176.480 ;
        RECT 3.220 165.600 2616.000 175.080 ;
        RECT 3.220 164.200 2615.600 165.600 ;
        RECT 3.220 154.720 2616.000 164.200 ;
        RECT 3.220 153.320 2615.600 154.720 ;
        RECT 3.220 143.840 2616.000 153.320 ;
        RECT 3.220 142.440 2615.600 143.840 ;
        RECT 3.220 132.960 2616.000 142.440 ;
        RECT 3.220 131.560 2615.600 132.960 ;
        RECT 3.220 122.080 2616.000 131.560 ;
        RECT 3.220 120.680 2615.600 122.080 ;
        RECT 3.220 111.200 2616.000 120.680 ;
        RECT 3.220 109.800 2615.600 111.200 ;
        RECT 3.220 100.320 2616.000 109.800 ;
        RECT 3.220 98.920 2615.600 100.320 ;
        RECT 3.220 89.440 2616.000 98.920 ;
        RECT 3.220 88.040 2615.600 89.440 ;
        RECT 3.220 78.560 2616.000 88.040 ;
        RECT 3.220 77.160 2615.600 78.560 ;
        RECT 3.220 67.680 2616.000 77.160 ;
        RECT 3.220 66.280 2615.600 67.680 ;
        RECT 3.220 56.800 2616.000 66.280 ;
        RECT 3.220 55.400 2615.600 56.800 ;
        RECT 3.220 45.920 2616.000 55.400 ;
        RECT 3.220 44.520 2615.600 45.920 ;
        RECT 3.220 35.040 2616.000 44.520 ;
        RECT 3.220 33.640 2615.600 35.040 ;
        RECT 3.220 24.160 2616.000 33.640 ;
        RECT 3.220 22.760 2615.600 24.160 ;
        RECT 3.220 13.280 2616.000 22.760 ;
        RECT 3.220 12.415 2615.600 13.280 ;
      LAYER met4 ;
        RECT 56.025 658.205 75.240 809.705 ;
        RECT 77.640 658.205 86.840 809.705 ;
        RECT 89.240 658.205 125.240 809.705 ;
        RECT 127.640 658.205 136.840 809.705 ;
        RECT 139.240 658.205 175.240 809.705 ;
        RECT 177.640 658.205 186.840 809.705 ;
        RECT 189.240 658.205 225.240 809.705 ;
        RECT 227.640 658.205 236.840 809.705 ;
        RECT 239.240 658.205 275.240 809.705 ;
        RECT 277.640 658.205 286.840 809.705 ;
        RECT 289.240 658.205 325.240 809.705 ;
        RECT 327.640 658.205 336.840 809.705 ;
        RECT 339.240 659.980 375.240 809.705 ;
        RECT 377.640 659.980 386.840 809.705 ;
        RECT 339.240 658.205 386.840 659.980 ;
        RECT 389.240 658.205 425.240 809.705 ;
        RECT 427.640 658.205 436.840 809.705 ;
        RECT 439.240 658.205 475.240 809.705 ;
        RECT 477.640 658.205 486.840 809.705 ;
        RECT 489.240 658.205 525.240 809.705 ;
        RECT 527.640 658.205 536.840 809.705 ;
        RECT 539.240 658.205 575.240 809.705 ;
        RECT 577.640 658.205 586.840 809.705 ;
        RECT 589.240 658.205 625.240 809.705 ;
        RECT 627.640 658.205 636.840 809.705 ;
        RECT 639.240 658.205 675.240 809.705 ;
        RECT 677.640 658.205 686.840 809.705 ;
        RECT 689.240 658.205 725.240 809.705 ;
        RECT 727.640 658.205 736.840 809.705 ;
        RECT 739.240 658.205 775.240 809.705 ;
        RECT 777.640 658.205 786.840 809.705 ;
        RECT 789.240 658.205 825.240 809.705 ;
        RECT 827.640 659.980 836.840 809.705 ;
        RECT 839.240 659.980 875.240 809.705 ;
        RECT 827.640 658.205 875.240 659.980 ;
        RECT 56.025 240.275 875.240 658.205 ;
        RECT 56.025 148.415 75.240 240.275 ;
        RECT 77.640 148.415 86.840 240.275 ;
        RECT 89.240 148.415 125.240 240.275 ;
        RECT 127.640 148.415 136.840 240.275 ;
        RECT 139.240 148.415 175.240 240.275 ;
        RECT 177.640 148.415 186.840 240.275 ;
        RECT 189.240 148.415 225.240 240.275 ;
        RECT 227.640 148.415 236.840 240.275 ;
        RECT 239.240 148.415 275.240 240.275 ;
        RECT 277.640 148.415 286.840 240.275 ;
        RECT 289.240 148.415 325.240 240.275 ;
        RECT 327.640 148.415 336.840 240.275 ;
        RECT 339.240 148.415 375.240 240.275 ;
        RECT 377.640 148.415 386.840 240.275 ;
        RECT 389.240 148.415 425.240 240.275 ;
        RECT 427.640 148.415 436.840 240.275 ;
        RECT 439.240 148.415 475.240 240.275 ;
        RECT 477.640 148.415 486.840 240.275 ;
        RECT 489.240 148.415 525.240 240.275 ;
        RECT 527.640 148.415 536.840 240.275 ;
        RECT 539.240 148.415 575.240 240.275 ;
        RECT 577.640 148.415 586.840 240.275 ;
        RECT 589.240 148.415 625.240 240.275 ;
        RECT 627.640 148.415 636.840 240.275 ;
        RECT 639.240 148.415 675.240 240.275 ;
        RECT 677.640 148.415 686.840 240.275 ;
        RECT 689.240 148.415 725.240 240.275 ;
        RECT 727.640 148.415 736.840 240.275 ;
        RECT 739.240 148.415 775.240 240.275 ;
        RECT 777.640 148.415 786.840 240.275 ;
        RECT 789.240 148.415 825.240 240.275 ;
        RECT 827.640 148.415 836.840 240.275 ;
        RECT 839.240 148.415 875.240 240.275 ;
        RECT 877.640 148.415 886.840 809.705 ;
        RECT 889.240 148.415 925.240 809.705 ;
        RECT 927.640 148.415 936.840 809.705 ;
        RECT 939.240 148.415 975.240 809.705 ;
        RECT 977.640 148.415 986.840 809.705 ;
        RECT 989.240 148.415 1025.240 809.705 ;
        RECT 1027.640 148.415 1036.840 809.705 ;
        RECT 1039.240 148.415 1075.240 809.705 ;
        RECT 1077.640 148.415 1086.840 809.705 ;
        RECT 1089.240 148.415 1125.240 809.705 ;
        RECT 1127.640 148.415 1136.840 809.705 ;
        RECT 1139.240 148.415 1175.240 809.705 ;
        RECT 1177.640 148.415 1186.840 809.705 ;
        RECT 1189.240 148.415 1225.240 809.705 ;
        RECT 1227.640 148.415 1236.840 809.705 ;
        RECT 1239.240 148.415 1275.240 809.705 ;
        RECT 1277.640 148.415 1286.840 809.705 ;
        RECT 1289.240 148.415 1325.240 809.705 ;
        RECT 1327.640 148.415 1336.840 809.705 ;
        RECT 1339.240 148.415 1375.240 809.705 ;
        RECT 1377.640 148.415 1386.840 809.705 ;
        RECT 1389.240 148.415 1425.240 809.705 ;
        RECT 1427.640 148.415 1436.840 809.705 ;
        RECT 1439.240 148.415 1475.240 809.705 ;
        RECT 1477.640 148.415 1486.840 809.705 ;
        RECT 1489.240 148.415 1525.240 809.705 ;
        RECT 1527.640 148.415 1536.840 809.705 ;
        RECT 1539.240 148.415 1575.240 809.705 ;
        RECT 1577.640 148.415 1586.840 809.705 ;
        RECT 1589.240 148.415 1625.240 809.705 ;
        RECT 1627.640 148.415 1636.840 809.705 ;
        RECT 1639.240 148.415 1675.240 809.705 ;
        RECT 1677.640 148.415 1686.840 809.705 ;
        RECT 1689.240 148.415 1725.240 809.705 ;
        RECT 1727.640 148.415 1736.840 809.705 ;
        RECT 1739.240 148.415 1775.240 809.705 ;
        RECT 1777.640 148.415 1786.840 809.705 ;
        RECT 1789.240 148.415 1825.240 809.705 ;
        RECT 1827.640 148.415 1836.840 809.705 ;
        RECT 1839.240 148.415 1875.240 809.705 ;
        RECT 1877.640 148.415 1886.840 809.705 ;
        RECT 1889.240 148.415 1925.240 809.705 ;
        RECT 1927.640 148.415 1936.840 809.705 ;
        RECT 1939.240 148.415 1975.240 809.705 ;
        RECT 1977.640 148.415 1986.840 809.705 ;
        RECT 1989.240 148.415 2025.240 809.705 ;
        RECT 2027.640 148.415 2036.840 809.705 ;
        RECT 2039.240 148.415 2075.240 809.705 ;
        RECT 2077.640 148.415 2086.840 809.705 ;
        RECT 2089.240 148.415 2125.240 809.705 ;
        RECT 2127.640 148.415 2136.840 809.705 ;
        RECT 2139.240 148.415 2175.240 809.705 ;
        RECT 2177.640 651.820 2186.840 809.705 ;
        RECT 2189.240 654.125 2225.240 809.705 ;
        RECT 2227.640 654.125 2236.840 809.705 ;
        RECT 2239.240 654.125 2275.240 809.705 ;
        RECT 2277.640 654.125 2286.840 809.705 ;
        RECT 2289.240 654.125 2325.240 809.705 ;
        RECT 2327.640 654.125 2336.840 809.705 ;
        RECT 2339.240 654.125 2375.240 809.705 ;
        RECT 2377.640 654.125 2386.840 809.705 ;
        RECT 2389.240 654.125 2425.240 809.705 ;
        RECT 2427.640 654.125 2436.840 809.705 ;
        RECT 2439.240 654.125 2475.240 809.705 ;
        RECT 2477.640 654.125 2486.840 809.705 ;
        RECT 2489.240 654.125 2525.240 809.705 ;
        RECT 2527.640 654.125 2536.840 809.705 ;
        RECT 2539.240 654.125 2575.240 809.705 ;
        RECT 2189.240 651.820 2575.240 654.125 ;
        RECT 2177.640 258.635 2575.240 651.820 ;
        RECT 2177.640 242.580 2225.240 258.635 ;
        RECT 2177.640 148.415 2186.840 242.580 ;
        RECT 2189.240 148.415 2225.240 242.580 ;
        RECT 2227.640 148.415 2236.840 258.635 ;
        RECT 2239.240 148.415 2275.240 258.635 ;
        RECT 2277.640 148.415 2286.840 258.635 ;
        RECT 2289.240 148.415 2325.240 258.635 ;
        RECT 2327.640 148.415 2336.840 258.635 ;
        RECT 2339.240 148.415 2375.240 258.635 ;
        RECT 2377.640 148.415 2386.840 258.635 ;
        RECT 2389.240 148.415 2425.240 258.635 ;
        RECT 2427.640 148.415 2436.840 258.635 ;
        RECT 2439.240 148.415 2475.240 258.635 ;
        RECT 2477.640 148.415 2486.840 258.635 ;
        RECT 2489.240 148.415 2525.240 258.635 ;
        RECT 2527.640 148.415 2536.840 258.635 ;
        RECT 2539.240 148.415 2575.240 258.635 ;
        RECT 2577.640 148.415 2586.840 809.705 ;
        RECT 2589.240 658.880 2605.145 809.705 ;
        RECT 2589.240 238.720 2594.580 658.880 ;
        RECT 2596.980 238.720 2605.145 658.880 ;
        RECT 2589.240 148.415 2605.145 238.720 ;
      LAYER met5 ;
        RECT 457.820 794.250 2591.060 798.100 ;
        RECT 457.820 782.650 2591.060 789.450 ;
        RECT 457.820 744.250 2591.060 777.850 ;
        RECT 457.820 732.650 2591.060 739.450 ;
        RECT 457.820 694.250 2591.060 727.850 ;
        RECT 457.820 682.650 2591.060 689.450 ;
        RECT 457.820 644.250 2591.060 677.850 ;
        RECT 457.820 632.650 2591.060 639.450 ;
        RECT 457.820 594.250 2591.060 627.850 ;
        RECT 457.820 582.650 2591.060 589.450 ;
        RECT 457.820 544.250 2591.060 577.850 ;
        RECT 457.820 532.650 2591.060 539.450 ;
        RECT 457.820 494.250 2591.060 527.850 ;
        RECT 457.820 482.650 2591.060 489.450 ;
        RECT 457.820 444.250 2591.060 477.850 ;
        RECT 457.820 432.650 2591.060 439.450 ;
        RECT 457.820 394.250 2591.060 427.850 ;
        RECT 457.820 382.650 2591.060 389.450 ;
        RECT 457.820 344.250 2591.060 377.850 ;
        RECT 457.820 332.650 2591.060 339.450 ;
        RECT 457.820 317.100 2591.060 327.850 ;
  END
END mgmt_core_wrapper
END LIBRARY

