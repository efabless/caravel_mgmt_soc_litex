VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_core_wrapper
  CLASS BLOCK ;
  FOREIGN mgmt_core_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2500.000 BY 720.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -5.380 -0.020 -3.780 718.100 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 -0.020 2505.020 1.580 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 716.500 2505.020 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2503.420 -0.020 2505.020 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 32.640 -0.020 34.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.640 -0.020 84.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 132.640 -0.020 134.240 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 132.640 585.510 134.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 182.640 -0.020 184.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 232.640 -0.020 234.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 232.640 554.875 234.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 282.640 -0.020 284.240 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 282.640 585.510 284.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 332.640 -0.020 334.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 332.640 554.875 334.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 382.640 -0.020 384.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 382.640 554.875 384.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 432.640 -0.020 434.240 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 432.640 585.510 434.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 482.640 -0.020 484.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 482.640 554.875 484.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 532.640 -0.020 534.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 532.640 554.875 534.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 582.640 -0.020 584.240 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 582.640 585.510 584.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.640 -0.020 634.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 632.640 554.875 634.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 682.640 -0.020 684.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 682.640 554.875 684.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 732.640 -0.020 734.240 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 732.640 585.510 734.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 782.640 -0.020 784.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 782.640 554.875 784.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 832.640 -0.020 834.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 832.640 554.875 834.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 882.640 -0.020 884.240 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 882.640 585.510 884.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 932.640 -0.020 934.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 932.640 554.875 934.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 982.640 -0.020 984.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 982.640 554.875 984.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1032.640 -0.020 1034.240 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 1032.640 585.510 1034.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1082.640 -0.020 1084.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 1082.640 554.875 1084.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1132.640 -0.020 1134.240 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 1132.640 554.875 1134.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1182.640 -0.020 1184.240 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 1182.640 585.510 1184.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1232.640 -0.020 1234.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1282.640 -0.020 1284.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1332.640 -0.020 1334.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1382.640 -0.020 1384.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1432.640 -0.020 1434.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1482.640 -0.020 1484.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1532.640 -0.020 1534.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1582.640 -0.020 1584.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1632.640 -0.020 1634.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1682.640 -0.020 1684.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1732.640 -0.020 1734.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1782.640 -0.020 1784.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1832.640 -0.020 1834.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1882.640 -0.020 1884.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1932.640 -0.020 1934.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1982.640 -0.020 1984.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2032.640 -0.020 2034.240 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2032.640 581.160 2034.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2082.640 -0.020 2084.240 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2082.640 581.160 2084.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2132.640 -0.020 2134.240 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2132.640 581.160 2134.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2182.640 -0.020 2184.240 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2182.640 581.160 2184.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.640 -0.020 2234.240 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2232.640 581.160 2234.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2282.640 -0.020 2284.240 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2282.640 581.160 2284.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2332.640 -0.020 2334.240 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2332.640 581.160 2334.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2382.640 -0.020 2384.240 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2382.640 581.160 2384.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2432.640 -0.020 2434.240 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2432.640 581.160 2434.240 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2482.640 -0.020 2484.240 718.100 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 38.330 2505.020 39.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 88.330 2505.020 89.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 138.330 2505.020 139.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 188.330 2505.020 189.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 238.330 2505.020 239.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 288.330 2505.020 289.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 338.330 2505.020 339.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 388.330 2505.020 389.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 438.330 2505.020 439.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 488.330 2505.020 489.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 538.330 2505.020 539.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 588.330 2505.020 589.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 638.330 2505.020 639.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 688.330 2505.020 689.930 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -2.080 3.280 -0.480 714.800 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 3.280 2501.720 4.880 ;
    END
    PORT
      LAYER met5 ;
        RECT -2.080 713.200 2501.720 714.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 2500.120 3.280 2501.720 714.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 -0.020 22.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.040 -0.020 72.640 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 71.040 585.510 72.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.040 -0.020 122.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.040 -0.020 172.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.040 -0.020 222.640 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 221.040 585.510 222.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 271.040 -0.020 272.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 271.040 554.875 272.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 -0.020 322.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 321.040 554.875 322.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.040 -0.020 372.640 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 371.040 585.510 372.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 421.040 -0.020 422.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 421.040 554.875 422.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 -0.020 472.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 471.040 554.875 472.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 521.040 -0.020 522.640 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 521.040 585.510 522.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.040 -0.020 572.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.040 554.875 572.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 -0.020 622.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 621.040 554.875 622.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.040 -0.020 672.640 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 671.040 585.510 672.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 721.040 -0.020 722.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 721.040 554.875 722.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 -0.020 772.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 771.040 554.875 772.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 821.040 -0.020 822.640 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 821.040 585.510 822.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 871.040 -0.020 872.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 871.040 554.875 872.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 -0.020 922.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 921.040 554.875 922.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 971.040 -0.020 972.640 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 971.040 585.510 972.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.040 -0.020 1022.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.040 554.875 1022.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1071.040 -0.020 1072.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 1071.040 554.875 1072.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1121.040 -0.020 1122.640 52.470 ;
    END
    PORT
      LAYER met4 ;
        RECT 1121.040 585.510 1122.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1171.040 -0.020 1172.640 104.185 ;
    END
    PORT
      LAYER met4 ;
        RECT 1171.040 554.875 1172.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1221.040 -0.020 1222.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1271.040 -0.020 1272.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1321.040 -0.020 1322.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1371.040 -0.020 1372.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1421.040 -0.020 1422.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1471.040 -0.020 1472.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1521.040 -0.020 1522.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.040 -0.020 1572.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1621.040 -0.020 1622.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1671.040 -0.020 1672.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1721.040 -0.020 1722.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1771.040 -0.020 1772.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1821.040 -0.020 1822.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1871.040 -0.020 1872.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1921.040 -0.020 1922.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 1971.040 -0.020 1972.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2021.040 -0.020 2022.640 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2021.040 581.160 2022.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2071.040 -0.020 2072.640 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2071.040 581.160 2072.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2121.040 -0.020 2122.640 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2121.040 581.160 2122.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.040 -0.020 2172.640 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.040 581.160 2172.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2221.040 -0.020 2222.640 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2221.040 581.160 2222.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2271.040 -0.020 2272.640 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2271.040 581.160 2272.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2321.040 -0.020 2322.640 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2321.040 581.160 2322.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2371.040 -0.020 2372.640 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2371.040 581.160 2372.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2421.040 -0.020 2422.640 69.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2421.040 581.160 2422.640 718.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2471.040 -0.020 2472.640 718.100 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 26.730 2505.020 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 76.730 2505.020 78.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 126.730 2505.020 128.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 176.730 2505.020 178.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 226.730 2505.020 228.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 276.730 2505.020 278.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 326.730 2505.020 328.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 376.730 2505.020 378.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 426.730 2505.020 428.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 476.730 2505.020 478.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 526.730 2505.020 528.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 576.730 2505.020 578.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 626.730 2505.020 628.330 ;
    END
    PORT
      LAYER met5 ;
        RECT -5.380 676.730 2505.020 678.330 ;
    END
  END VPWR
  PIN core_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1717.730 0.000 1718.010 4.000 ;
    END
  END core_clk
  PIN core_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1821.690 0.000 1821.970 4.000 ;
    END
  END core_rstn
  PIN debug_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 44.920 2500.000 45.520 ;
    END
  END debug_in
  PIN debug_mode
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 54.440 2500.000 55.040 ;
    END
  END debug_mode
  PIN debug_oeb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 63.960 2500.000 64.560 ;
    END
  END debug_oeb
  PIN debug_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 73.480 2500.000 74.080 ;
    END
  END debug_out
  PIN flash_clk
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 559.000 2500.000 559.600 ;
    END
  END flash_clk
  PIN flash_csb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 549.480 2500.000 550.080 ;
    END
  END flash_csb
  PIN flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 568.520 2500.000 569.120 ;
    END
  END flash_io0_di
  PIN flash_io0_do
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 578.040 2500.000 578.640 ;
    END
  END flash_io0_do
  PIN flash_io0_oeb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 587.560 2500.000 588.160 ;
    END
  END flash_io0_oeb
  PIN flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 597.080 2500.000 597.680 ;
    END
  END flash_io1_di
  PIN flash_io1_do
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 606.600 2500.000 607.200 ;
    END
  END flash_io1_do
  PIN flash_io1_oeb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 616.120 2500.000 616.720 ;
    END
  END flash_io1_oeb
  PIN flash_io2_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 625.640 2500.000 626.240 ;
    END
  END flash_io2_di
  PIN flash_io2_do
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 635.160 2500.000 635.760 ;
    END
  END flash_io2_do
  PIN flash_io2_oeb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 644.680 2500.000 645.280 ;
    END
  END flash_io2_oeb
  PIN flash_io3_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 654.200 2500.000 654.800 ;
    END
  END flash_io3_di
  PIN flash_io3_do
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 663.720 2500.000 664.320 ;
    END
  END flash_io3_do
  PIN flash_io3_oeb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 673.240 2500.000 673.840 ;
    END
  END flash_io3_oeb
  PIN gpio_in_pad
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1925.650 0.000 1925.930 4.000 ;
    END
  END gpio_in_pad
  PIN gpio_inenb_pad
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.610 0.000 2029.890 4.000 ;
    END
  END gpio_inenb_pad
  PIN gpio_mode0_pad
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2133.570 0.000 2133.850 4.000 ;
    END
  END gpio_mode0_pad
  PIN gpio_mode1_pad
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2237.530 0.000 2237.810 4.000 ;
    END
  END gpio_mode1_pad
  PIN gpio_out_pad
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2341.490 0.000 2341.770 4.000 ;
    END
  END gpio_out_pad
  PIN gpio_outenb_pad
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2445.450 0.000 2445.730 4.000 ;
    END
  END gpio_outenb_pad
  PIN hk_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 216.280 2500.000 216.880 ;
    END
  END hk_ack_i
  PIN hk_cyc_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 235.320 2500.000 235.920 ;
    END
  END hk_cyc_o
  PIN hk_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 244.840 2500.000 245.440 ;
    END
  END hk_dat_i[0]
  PIN hk_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 340.040 2500.000 340.640 ;
    END
  END hk_dat_i[10]
  PIN hk_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 349.560 2500.000 350.160 ;
    END
  END hk_dat_i[11]
  PIN hk_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 359.080 2500.000 359.680 ;
    END
  END hk_dat_i[12]
  PIN hk_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 368.600 2500.000 369.200 ;
    END
  END hk_dat_i[13]
  PIN hk_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 378.120 2500.000 378.720 ;
    END
  END hk_dat_i[14]
  PIN hk_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 387.640 2500.000 388.240 ;
    END
  END hk_dat_i[15]
  PIN hk_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 397.160 2500.000 397.760 ;
    END
  END hk_dat_i[16]
  PIN hk_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 406.680 2500.000 407.280 ;
    END
  END hk_dat_i[17]
  PIN hk_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 416.200 2500.000 416.800 ;
    END
  END hk_dat_i[18]
  PIN hk_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 425.720 2500.000 426.320 ;
    END
  END hk_dat_i[19]
  PIN hk_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 254.360 2500.000 254.960 ;
    END
  END hk_dat_i[1]
  PIN hk_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 435.240 2500.000 435.840 ;
    END
  END hk_dat_i[20]
  PIN hk_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 444.760 2500.000 445.360 ;
    END
  END hk_dat_i[21]
  PIN hk_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 454.280 2500.000 454.880 ;
    END
  END hk_dat_i[22]
  PIN hk_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 463.800 2500.000 464.400 ;
    END
  END hk_dat_i[23]
  PIN hk_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 473.320 2500.000 473.920 ;
    END
  END hk_dat_i[24]
  PIN hk_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 482.840 2500.000 483.440 ;
    END
  END hk_dat_i[25]
  PIN hk_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 492.360 2500.000 492.960 ;
    END
  END hk_dat_i[26]
  PIN hk_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 501.880 2500.000 502.480 ;
    END
  END hk_dat_i[27]
  PIN hk_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 511.400 2500.000 512.000 ;
    END
  END hk_dat_i[28]
  PIN hk_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 520.920 2500.000 521.520 ;
    END
  END hk_dat_i[29]
  PIN hk_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 263.880 2500.000 264.480 ;
    END
  END hk_dat_i[2]
  PIN hk_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 530.440 2500.000 531.040 ;
    END
  END hk_dat_i[30]
  PIN hk_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 539.960 2500.000 540.560 ;
    END
  END hk_dat_i[31]
  PIN hk_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 273.400 2500.000 274.000 ;
    END
  END hk_dat_i[3]
  PIN hk_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 282.920 2500.000 283.520 ;
    END
  END hk_dat_i[4]
  PIN hk_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 292.440 2500.000 293.040 ;
    END
  END hk_dat_i[5]
  PIN hk_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 301.960 2500.000 302.560 ;
    END
  END hk_dat_i[6]
  PIN hk_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 311.480 2500.000 312.080 ;
    END
  END hk_dat_i[7]
  PIN hk_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 321.000 2500.000 321.600 ;
    END
  END hk_dat_i[8]
  PIN hk_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 330.520 2500.000 331.120 ;
    END
  END hk_dat_i[9]
  PIN hk_stb_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 225.800 2500.000 226.400 ;
    END
  END hk_stb_o
  PIN irq[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2387.030 716.000 2387.310 720.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.710 716.000 2390.990 720.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2394.390 716.000 2394.670 720.000 ;
    END
  END irq[2]
  PIN irq[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 111.560 2500.000 112.160 ;
    END
  END irq[3]
  PIN irq[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 102.040 2500.000 102.640 ;
    END
  END irq[4]
  PIN irq[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 92.520 2500.000 93.120 ;
    END
  END irq[5]
  PIN la_iena[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 716.000 105.710 720.000 ;
    END
  END la_iena[0]
  PIN la_iena[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1577.430 716.000 1577.710 720.000 ;
    END
  END la_iena[100]
  PIN la_iena[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.150 716.000 1592.430 720.000 ;
    END
  END la_iena[101]
  PIN la_iena[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1606.870 716.000 1607.150 720.000 ;
    END
  END la_iena[102]
  PIN la_iena[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.590 716.000 1621.870 720.000 ;
    END
  END la_iena[103]
  PIN la_iena[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1636.310 716.000 1636.590 720.000 ;
    END
  END la_iena[104]
  PIN la_iena[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.030 716.000 1651.310 720.000 ;
    END
  END la_iena[105]
  PIN la_iena[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1665.750 716.000 1666.030 720.000 ;
    END
  END la_iena[106]
  PIN la_iena[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1680.470 716.000 1680.750 720.000 ;
    END
  END la_iena[107]
  PIN la_iena[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1695.190 716.000 1695.470 720.000 ;
    END
  END la_iena[108]
  PIN la_iena[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1709.910 716.000 1710.190 720.000 ;
    END
  END la_iena[109]
  PIN la_iena[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 716.000 252.910 720.000 ;
    END
  END la_iena[10]
  PIN la_iena[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1724.630 716.000 1724.910 720.000 ;
    END
  END la_iena[110]
  PIN la_iena[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1739.350 716.000 1739.630 720.000 ;
    END
  END la_iena[111]
  PIN la_iena[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.070 716.000 1754.350 720.000 ;
    END
  END la_iena[112]
  PIN la_iena[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1768.790 716.000 1769.070 720.000 ;
    END
  END la_iena[113]
  PIN la_iena[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.510 716.000 1783.790 720.000 ;
    END
  END la_iena[114]
  PIN la_iena[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1798.230 716.000 1798.510 720.000 ;
    END
  END la_iena[115]
  PIN la_iena[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1812.950 716.000 1813.230 720.000 ;
    END
  END la_iena[116]
  PIN la_iena[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1827.670 716.000 1827.950 720.000 ;
    END
  END la_iena[117]
  PIN la_iena[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1842.390 716.000 1842.670 720.000 ;
    END
  END la_iena[118]
  PIN la_iena[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1857.110 716.000 1857.390 720.000 ;
    END
  END la_iena[119]
  PIN la_iena[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 716.000 267.630 720.000 ;
    END
  END la_iena[11]
  PIN la_iena[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1871.830 716.000 1872.110 720.000 ;
    END
  END la_iena[120]
  PIN la_iena[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1886.550 716.000 1886.830 720.000 ;
    END
  END la_iena[121]
  PIN la_iena[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1901.270 716.000 1901.550 720.000 ;
    END
  END la_iena[122]
  PIN la_iena[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1915.990 716.000 1916.270 720.000 ;
    END
  END la_iena[123]
  PIN la_iena[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1930.710 716.000 1930.990 720.000 ;
    END
  END la_iena[124]
  PIN la_iena[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1945.430 716.000 1945.710 720.000 ;
    END
  END la_iena[125]
  PIN la_iena[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1960.150 716.000 1960.430 720.000 ;
    END
  END la_iena[126]
  PIN la_iena[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1974.870 716.000 1975.150 720.000 ;
    END
  END la_iena[127]
  PIN la_iena[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.070 716.000 282.350 720.000 ;
    END
  END la_iena[12]
  PIN la_iena[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 716.000 297.070 720.000 ;
    END
  END la_iena[13]
  PIN la_iena[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.510 716.000 311.790 720.000 ;
    END
  END la_iena[14]
  PIN la_iena[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 716.000 326.510 720.000 ;
    END
  END la_iena[15]
  PIN la_iena[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.950 716.000 341.230 720.000 ;
    END
  END la_iena[16]
  PIN la_iena[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 716.000 355.950 720.000 ;
    END
  END la_iena[17]
  PIN la_iena[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 716.000 370.670 720.000 ;
    END
  END la_iena[18]
  PIN la_iena[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 716.000 385.390 720.000 ;
    END
  END la_iena[19]
  PIN la_iena[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 716.000 120.430 720.000 ;
    END
  END la_iena[1]
  PIN la_iena[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.830 716.000 400.110 720.000 ;
    END
  END la_iena[20]
  PIN la_iena[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.550 716.000 414.830 720.000 ;
    END
  END la_iena[21]
  PIN la_iena[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.270 716.000 429.550 720.000 ;
    END
  END la_iena[22]
  PIN la_iena[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 716.000 444.270 720.000 ;
    END
  END la_iena[23]
  PIN la_iena[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.710 716.000 458.990 720.000 ;
    END
  END la_iena[24]
  PIN la_iena[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 716.000 473.710 720.000 ;
    END
  END la_iena[25]
  PIN la_iena[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 716.000 488.430 720.000 ;
    END
  END la_iena[26]
  PIN la_iena[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.870 716.000 503.150 720.000 ;
    END
  END la_iena[27]
  PIN la_iena[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 716.000 517.870 720.000 ;
    END
  END la_iena[28]
  PIN la_iena[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 716.000 532.590 720.000 ;
    END
  END la_iena[29]
  PIN la_iena[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.870 716.000 135.150 720.000 ;
    END
  END la_iena[2]
  PIN la_iena[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.030 716.000 547.310 720.000 ;
    END
  END la_iena[30]
  PIN la_iena[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 716.000 562.030 720.000 ;
    END
  END la_iena[31]
  PIN la_iena[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 716.000 576.750 720.000 ;
    END
  END la_iena[32]
  PIN la_iena[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.190 716.000 591.470 720.000 ;
    END
  END la_iena[33]
  PIN la_iena[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.910 716.000 606.190 720.000 ;
    END
  END la_iena[34]
  PIN la_iena[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.630 716.000 620.910 720.000 ;
    END
  END la_iena[35]
  PIN la_iena[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 716.000 635.630 720.000 ;
    END
  END la_iena[36]
  PIN la_iena[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 716.000 650.350 720.000 ;
    END
  END la_iena[37]
  PIN la_iena[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.790 716.000 665.070 720.000 ;
    END
  END la_iena[38]
  PIN la_iena[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 679.510 716.000 679.790 720.000 ;
    END
  END la_iena[39]
  PIN la_iena[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 716.000 149.870 720.000 ;
    END
  END la_iena[3]
  PIN la_iena[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.230 716.000 694.510 720.000 ;
    END
  END la_iena[40]
  PIN la_iena[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.950 716.000 709.230 720.000 ;
    END
  END la_iena[41]
  PIN la_iena[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.670 716.000 723.950 720.000 ;
    END
  END la_iena[42]
  PIN la_iena[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.390 716.000 738.670 720.000 ;
    END
  END la_iena[43]
  PIN la_iena[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.110 716.000 753.390 720.000 ;
    END
  END la_iena[44]
  PIN la_iena[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 716.000 768.110 720.000 ;
    END
  END la_iena[45]
  PIN la_iena[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 716.000 782.830 720.000 ;
    END
  END la_iena[46]
  PIN la_iena[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 797.270 716.000 797.550 720.000 ;
    END
  END la_iena[47]
  PIN la_iena[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.990 716.000 812.270 720.000 ;
    END
  END la_iena[48]
  PIN la_iena[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 826.710 716.000 826.990 720.000 ;
    END
  END la_iena[49]
  PIN la_iena[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 716.000 164.590 720.000 ;
    END
  END la_iena[4]
  PIN la_iena[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.430 716.000 841.710 720.000 ;
    END
  END la_iena[50]
  PIN la_iena[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.150 716.000 856.430 720.000 ;
    END
  END la_iena[51]
  PIN la_iena[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.870 716.000 871.150 720.000 ;
    END
  END la_iena[52]
  PIN la_iena[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.590 716.000 885.870 720.000 ;
    END
  END la_iena[53]
  PIN la_iena[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.310 716.000 900.590 720.000 ;
    END
  END la_iena[54]
  PIN la_iena[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.030 716.000 915.310 720.000 ;
    END
  END la_iena[55]
  PIN la_iena[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.750 716.000 930.030 720.000 ;
    END
  END la_iena[56]
  PIN la_iena[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.470 716.000 944.750 720.000 ;
    END
  END la_iena[57]
  PIN la_iena[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.190 716.000 959.470 720.000 ;
    END
  END la_iena[58]
  PIN la_iena[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 973.910 716.000 974.190 720.000 ;
    END
  END la_iena[59]
  PIN la_iena[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 716.000 179.310 720.000 ;
    END
  END la_iena[5]
  PIN la_iena[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 988.630 716.000 988.910 720.000 ;
    END
  END la_iena[60]
  PIN la_iena[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1003.350 716.000 1003.630 720.000 ;
    END
  END la_iena[61]
  PIN la_iena[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.070 716.000 1018.350 720.000 ;
    END
  END la_iena[62]
  PIN la_iena[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1032.790 716.000 1033.070 720.000 ;
    END
  END la_iena[63]
  PIN la_iena[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.510 716.000 1047.790 720.000 ;
    END
  END la_iena[64]
  PIN la_iena[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1062.230 716.000 1062.510 720.000 ;
    END
  END la_iena[65]
  PIN la_iena[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1076.950 716.000 1077.230 720.000 ;
    END
  END la_iena[66]
  PIN la_iena[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.670 716.000 1091.950 720.000 ;
    END
  END la_iena[67]
  PIN la_iena[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.390 716.000 1106.670 720.000 ;
    END
  END la_iena[68]
  PIN la_iena[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1121.110 716.000 1121.390 720.000 ;
    END
  END la_iena[69]
  PIN la_iena[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 716.000 194.030 720.000 ;
    END
  END la_iena[6]
  PIN la_iena[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1135.830 716.000 1136.110 720.000 ;
    END
  END la_iena[70]
  PIN la_iena[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1150.550 716.000 1150.830 720.000 ;
    END
  END la_iena[71]
  PIN la_iena[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.270 716.000 1165.550 720.000 ;
    END
  END la_iena[72]
  PIN la_iena[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1179.990 716.000 1180.270 720.000 ;
    END
  END la_iena[73]
  PIN la_iena[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.710 716.000 1194.990 720.000 ;
    END
  END la_iena[74]
  PIN la_iena[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1209.430 716.000 1209.710 720.000 ;
    END
  END la_iena[75]
  PIN la_iena[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.150 716.000 1224.430 720.000 ;
    END
  END la_iena[76]
  PIN la_iena[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.870 716.000 1239.150 720.000 ;
    END
  END la_iena[77]
  PIN la_iena[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.590 716.000 1253.870 720.000 ;
    END
  END la_iena[78]
  PIN la_iena[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.310 716.000 1268.590 720.000 ;
    END
  END la_iena[79]
  PIN la_iena[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.470 716.000 208.750 720.000 ;
    END
  END la_iena[7]
  PIN la_iena[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1283.030 716.000 1283.310 720.000 ;
    END
  END la_iena[80]
  PIN la_iena[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.750 716.000 1298.030 720.000 ;
    END
  END la_iena[81]
  PIN la_iena[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.470 716.000 1312.750 720.000 ;
    END
  END la_iena[82]
  PIN la_iena[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1327.190 716.000 1327.470 720.000 ;
    END
  END la_iena[83]
  PIN la_iena[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1341.910 716.000 1342.190 720.000 ;
    END
  END la_iena[84]
  PIN la_iena[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.630 716.000 1356.910 720.000 ;
    END
  END la_iena[85]
  PIN la_iena[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1371.350 716.000 1371.630 720.000 ;
    END
  END la_iena[86]
  PIN la_iena[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.070 716.000 1386.350 720.000 ;
    END
  END la_iena[87]
  PIN la_iena[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1400.790 716.000 1401.070 720.000 ;
    END
  END la_iena[88]
  PIN la_iena[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.510 716.000 1415.790 720.000 ;
    END
  END la_iena[89]
  PIN la_iena[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 716.000 223.470 720.000 ;
    END
  END la_iena[8]
  PIN la_iena[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1430.230 716.000 1430.510 720.000 ;
    END
  END la_iena[90]
  PIN la_iena[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.950 716.000 1445.230 720.000 ;
    END
  END la_iena[91]
  PIN la_iena[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.670 716.000 1459.950 720.000 ;
    END
  END la_iena[92]
  PIN la_iena[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.390 716.000 1474.670 720.000 ;
    END
  END la_iena[93]
  PIN la_iena[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.110 716.000 1489.390 720.000 ;
    END
  END la_iena[94]
  PIN la_iena[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.830 716.000 1504.110 720.000 ;
    END
  END la_iena[95]
  PIN la_iena[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1518.550 716.000 1518.830 720.000 ;
    END
  END la_iena[96]
  PIN la_iena[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.270 716.000 1533.550 720.000 ;
    END
  END la_iena[97]
  PIN la_iena[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1547.990 716.000 1548.270 720.000 ;
    END
  END la_iena[98]
  PIN la_iena[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1562.710 716.000 1562.990 720.000 ;
    END
  END la_iena[99]
  PIN la_iena[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.910 716.000 238.190 720.000 ;
    END
  END la_iena[9]
  PIN la_input[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 716.000 109.390 720.000 ;
    END
  END la_input[0]
  PIN la_input[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.110 716.000 1581.390 720.000 ;
    END
  END la_input[100]
  PIN la_input[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1595.830 716.000 1596.110 720.000 ;
    END
  END la_input[101]
  PIN la_input[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.550 716.000 1610.830 720.000 ;
    END
  END la_input[102]
  PIN la_input[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1625.270 716.000 1625.550 720.000 ;
    END
  END la_input[103]
  PIN la_input[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.990 716.000 1640.270 720.000 ;
    END
  END la_input[104]
  PIN la_input[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1654.710 716.000 1654.990 720.000 ;
    END
  END la_input[105]
  PIN la_input[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.430 716.000 1669.710 720.000 ;
    END
  END la_input[106]
  PIN la_input[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1684.150 716.000 1684.430 720.000 ;
    END
  END la_input[107]
  PIN la_input[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1698.870 716.000 1699.150 720.000 ;
    END
  END la_input[108]
  PIN la_input[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1713.590 716.000 1713.870 720.000 ;
    END
  END la_input[109]
  PIN la_input[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.310 716.000 256.590 720.000 ;
    END
  END la_input[10]
  PIN la_input[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.310 716.000 1728.590 720.000 ;
    END
  END la_input[110]
  PIN la_input[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.030 716.000 1743.310 720.000 ;
    END
  END la_input[111]
  PIN la_input[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1757.750 716.000 1758.030 720.000 ;
    END
  END la_input[112]
  PIN la_input[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1772.470 716.000 1772.750 720.000 ;
    END
  END la_input[113]
  PIN la_input[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.190 716.000 1787.470 720.000 ;
    END
  END la_input[114]
  PIN la_input[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1801.910 716.000 1802.190 720.000 ;
    END
  END la_input[115]
  PIN la_input[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.630 716.000 1816.910 720.000 ;
    END
  END la_input[116]
  PIN la_input[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1831.350 716.000 1831.630 720.000 ;
    END
  END la_input[117]
  PIN la_input[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.070 716.000 1846.350 720.000 ;
    END
  END la_input[118]
  PIN la_input[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1860.790 716.000 1861.070 720.000 ;
    END
  END la_input[119]
  PIN la_input[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 716.000 271.310 720.000 ;
    END
  END la_input[11]
  PIN la_input[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1875.510 716.000 1875.790 720.000 ;
    END
  END la_input[120]
  PIN la_input[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.230 716.000 1890.510 720.000 ;
    END
  END la_input[121]
  PIN la_input[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.950 716.000 1905.230 720.000 ;
    END
  END la_input[122]
  PIN la_input[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1919.670 716.000 1919.950 720.000 ;
    END
  END la_input[123]
  PIN la_input[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1934.390 716.000 1934.670 720.000 ;
    END
  END la_input[124]
  PIN la_input[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1949.110 716.000 1949.390 720.000 ;
    END
  END la_input[125]
  PIN la_input[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1963.830 716.000 1964.110 720.000 ;
    END
  END la_input[126]
  PIN la_input[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1978.550 716.000 1978.830 720.000 ;
    END
  END la_input[127]
  PIN la_input[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 716.000 286.030 720.000 ;
    END
  END la_input[12]
  PIN la_input[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 716.000 300.750 720.000 ;
    END
  END la_input[13]
  PIN la_input[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.190 716.000 315.470 720.000 ;
    END
  END la_input[14]
  PIN la_input[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 716.000 330.190 720.000 ;
    END
  END la_input[15]
  PIN la_input[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 716.000 344.910 720.000 ;
    END
  END la_input[16]
  PIN la_input[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.350 716.000 359.630 720.000 ;
    END
  END la_input[17]
  PIN la_input[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.070 716.000 374.350 720.000 ;
    END
  END la_input[18]
  PIN la_input[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.790 716.000 389.070 720.000 ;
    END
  END la_input[19]
  PIN la_input[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.830 716.000 124.110 720.000 ;
    END
  END la_input[1]
  PIN la_input[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.510 716.000 403.790 720.000 ;
    END
  END la_input[20]
  PIN la_input[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 716.000 418.510 720.000 ;
    END
  END la_input[21]
  PIN la_input[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 716.000 433.230 720.000 ;
    END
  END la_input[22]
  PIN la_input[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 716.000 447.950 720.000 ;
    END
  END la_input[23]
  PIN la_input[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 716.000 462.670 720.000 ;
    END
  END la_input[24]
  PIN la_input[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 716.000 477.390 720.000 ;
    END
  END la_input[25]
  PIN la_input[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 716.000 492.110 720.000 ;
    END
  END la_input[26]
  PIN la_input[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.550 716.000 506.830 720.000 ;
    END
  END la_input[27]
  PIN la_input[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.270 716.000 521.550 720.000 ;
    END
  END la_input[28]
  PIN la_input[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 535.990 716.000 536.270 720.000 ;
    END
  END la_input[29]
  PIN la_input[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 716.000 138.830 720.000 ;
    END
  END la_input[2]
  PIN la_input[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 716.000 550.990 720.000 ;
    END
  END la_input[30]
  PIN la_input[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.430 716.000 565.710 720.000 ;
    END
  END la_input[31]
  PIN la_input[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 716.000 580.430 720.000 ;
    END
  END la_input[32]
  PIN la_input[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 594.870 716.000 595.150 720.000 ;
    END
  END la_input[33]
  PIN la_input[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 716.000 609.870 720.000 ;
    END
  END la_input[34]
  PIN la_input[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.310 716.000 624.590 720.000 ;
    END
  END la_input[35]
  PIN la_input[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 716.000 639.310 720.000 ;
    END
  END la_input[36]
  PIN la_input[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.750 716.000 654.030 720.000 ;
    END
  END la_input[37]
  PIN la_input[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.470 716.000 668.750 720.000 ;
    END
  END la_input[38]
  PIN la_input[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 716.000 683.470 720.000 ;
    END
  END la_input[39]
  PIN la_input[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.270 716.000 153.550 720.000 ;
    END
  END la_input[3]
  PIN la_input[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.910 716.000 698.190 720.000 ;
    END
  END la_input[40]
  PIN la_input[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.630 716.000 712.910 720.000 ;
    END
  END la_input[41]
  PIN la_input[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.350 716.000 727.630 720.000 ;
    END
  END la_input[42]
  PIN la_input[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.070 716.000 742.350 720.000 ;
    END
  END la_input[43]
  PIN la_input[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 756.790 716.000 757.070 720.000 ;
    END
  END la_input[44]
  PIN la_input[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 716.000 771.790 720.000 ;
    END
  END la_input[45]
  PIN la_input[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.230 716.000 786.510 720.000 ;
    END
  END la_input[46]
  PIN la_input[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.950 716.000 801.230 720.000 ;
    END
  END la_input[47]
  PIN la_input[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.670 716.000 815.950 720.000 ;
    END
  END la_input[48]
  PIN la_input[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.390 716.000 830.670 720.000 ;
    END
  END la_input[49]
  PIN la_input[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 716.000 168.270 720.000 ;
    END
  END la_input[4]
  PIN la_input[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 845.110 716.000 845.390 720.000 ;
    END
  END la_input[50]
  PIN la_input[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 716.000 860.110 720.000 ;
    END
  END la_input[51]
  PIN la_input[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 874.550 716.000 874.830 720.000 ;
    END
  END la_input[52]
  PIN la_input[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.270 716.000 889.550 720.000 ;
    END
  END la_input[53]
  PIN la_input[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 903.990 716.000 904.270 720.000 ;
    END
  END la_input[54]
  PIN la_input[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.710 716.000 918.990 720.000 ;
    END
  END la_input[55]
  PIN la_input[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.430 716.000 933.710 720.000 ;
    END
  END la_input[56]
  PIN la_input[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.150 716.000 948.430 720.000 ;
    END
  END la_input[57]
  PIN la_input[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.870 716.000 963.150 720.000 ;
    END
  END la_input[58]
  PIN la_input[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.590 716.000 977.870 720.000 ;
    END
  END la_input[59]
  PIN la_input[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.710 716.000 182.990 720.000 ;
    END
  END la_input[5]
  PIN la_input[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.310 716.000 992.590 720.000 ;
    END
  END la_input[60]
  PIN la_input[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.030 716.000 1007.310 720.000 ;
    END
  END la_input[61]
  PIN la_input[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1021.750 716.000 1022.030 720.000 ;
    END
  END la_input[62]
  PIN la_input[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.470 716.000 1036.750 720.000 ;
    END
  END la_input[63]
  PIN la_input[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.190 716.000 1051.470 720.000 ;
    END
  END la_input[64]
  PIN la_input[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.910 716.000 1066.190 720.000 ;
    END
  END la_input[65]
  PIN la_input[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.630 716.000 1080.910 720.000 ;
    END
  END la_input[66]
  PIN la_input[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.350 716.000 1095.630 720.000 ;
    END
  END la_input[67]
  PIN la_input[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.070 716.000 1110.350 720.000 ;
    END
  END la_input[68]
  PIN la_input[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.790 716.000 1125.070 720.000 ;
    END
  END la_input[69]
  PIN la_input[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.430 716.000 197.710 720.000 ;
    END
  END la_input[6]
  PIN la_input[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.510 716.000 1139.790 720.000 ;
    END
  END la_input[70]
  PIN la_input[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1154.230 716.000 1154.510 720.000 ;
    END
  END la_input[71]
  PIN la_input[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.950 716.000 1169.230 720.000 ;
    END
  END la_input[72]
  PIN la_input[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.670 716.000 1183.950 720.000 ;
    END
  END la_input[73]
  PIN la_input[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1198.390 716.000 1198.670 720.000 ;
    END
  END la_input[74]
  PIN la_input[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1213.110 716.000 1213.390 720.000 ;
    END
  END la_input[75]
  PIN la_input[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.830 716.000 1228.110 720.000 ;
    END
  END la_input[76]
  PIN la_input[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1242.550 716.000 1242.830 720.000 ;
    END
  END la_input[77]
  PIN la_input[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.270 716.000 1257.550 720.000 ;
    END
  END la_input[78]
  PIN la_input[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.990 716.000 1272.270 720.000 ;
    END
  END la_input[79]
  PIN la_input[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 716.000 212.430 720.000 ;
    END
  END la_input[7]
  PIN la_input[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1286.710 716.000 1286.990 720.000 ;
    END
  END la_input[80]
  PIN la_input[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.430 716.000 1301.710 720.000 ;
    END
  END la_input[81]
  PIN la_input[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1316.150 716.000 1316.430 720.000 ;
    END
  END la_input[82]
  PIN la_input[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1330.870 716.000 1331.150 720.000 ;
    END
  END la_input[83]
  PIN la_input[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1345.590 716.000 1345.870 720.000 ;
    END
  END la_input[84]
  PIN la_input[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1360.310 716.000 1360.590 720.000 ;
    END
  END la_input[85]
  PIN la_input[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1375.030 716.000 1375.310 720.000 ;
    END
  END la_input[86]
  PIN la_input[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1389.750 716.000 1390.030 720.000 ;
    END
  END la_input[87]
  PIN la_input[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1404.470 716.000 1404.750 720.000 ;
    END
  END la_input[88]
  PIN la_input[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.190 716.000 1419.470 720.000 ;
    END
  END la_input[89]
  PIN la_input[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 716.000 227.150 720.000 ;
    END
  END la_input[8]
  PIN la_input[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1433.910 716.000 1434.190 720.000 ;
    END
  END la_input[90]
  PIN la_input[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1448.630 716.000 1448.910 720.000 ;
    END
  END la_input[91]
  PIN la_input[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1463.350 716.000 1463.630 720.000 ;
    END
  END la_input[92]
  PIN la_input[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.070 716.000 1478.350 720.000 ;
    END
  END la_input[93]
  PIN la_input[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.790 716.000 1493.070 720.000 ;
    END
  END la_input[94]
  PIN la_input[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.510 716.000 1507.790 720.000 ;
    END
  END la_input[95]
  PIN la_input[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1522.230 716.000 1522.510 720.000 ;
    END
  END la_input[96]
  PIN la_input[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.950 716.000 1537.230 720.000 ;
    END
  END la_input[97]
  PIN la_input[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.670 716.000 1551.950 720.000 ;
    END
  END la_input[98]
  PIN la_input[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1566.390 716.000 1566.670 720.000 ;
    END
  END la_input[99]
  PIN la_input[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 716.000 241.870 720.000 ;
    END
  END la_input[9]
  PIN la_oenb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 716.000 113.070 720.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1584.790 716.000 1585.070 720.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1599.510 716.000 1599.790 720.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1614.230 716.000 1614.510 720.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1628.950 716.000 1629.230 720.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.670 716.000 1643.950 720.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1658.390 716.000 1658.670 720.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1673.110 716.000 1673.390 720.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.830 716.000 1688.110 720.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1702.550 716.000 1702.830 720.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1717.270 716.000 1717.550 720.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 716.000 260.270 720.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1731.990 716.000 1732.270 720.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.710 716.000 1746.990 720.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.430 716.000 1761.710 720.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.150 716.000 1776.430 720.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1790.870 716.000 1791.150 720.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.590 716.000 1805.870 720.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1820.310 716.000 1820.590 720.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1835.030 716.000 1835.310 720.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1849.750 716.000 1850.030 720.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.470 716.000 1864.750 720.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 716.000 274.990 720.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1879.190 716.000 1879.470 720.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1893.910 716.000 1894.190 720.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1908.630 716.000 1908.910 720.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.350 716.000 1923.630 720.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1938.070 716.000 1938.350 720.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1952.790 716.000 1953.070 720.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1967.510 716.000 1967.790 720.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1982.230 716.000 1982.510 720.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 716.000 289.710 720.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 716.000 304.430 720.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 716.000 319.150 720.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 716.000 333.870 720.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 348.310 716.000 348.590 720.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.030 716.000 363.310 720.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 716.000 378.030 720.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.470 716.000 392.750 720.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 716.000 127.790 720.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.190 716.000 407.470 720.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 716.000 422.190 720.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 436.630 716.000 436.910 720.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 716.000 451.630 720.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 716.000 466.350 720.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.790 716.000 481.070 720.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 716.000 495.790 720.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.230 716.000 510.510 720.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 716.000 525.230 720.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.670 716.000 539.950 720.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.230 716.000 142.510 720.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.390 716.000 554.670 720.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.110 716.000 569.390 720.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 716.000 584.110 720.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.550 716.000 598.830 720.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 716.000 613.550 720.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.990 716.000 628.270 720.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.710 716.000 642.990 720.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 716.000 657.710 720.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.150 716.000 672.430 720.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.870 716.000 687.150 720.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 716.000 157.230 720.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 701.590 716.000 701.870 720.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.310 716.000 716.590 720.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 716.000 731.310 720.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 745.750 716.000 746.030 720.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.470 716.000 760.750 720.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.190 716.000 775.470 720.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 789.910 716.000 790.190 720.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.630 716.000 804.910 720.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.350 716.000 819.630 720.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 834.070 716.000 834.350 720.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 171.670 716.000 171.950 720.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.790 716.000 849.070 720.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.510 716.000 863.790 720.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.230 716.000 878.510 720.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.950 716.000 893.230 720.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.670 716.000 907.950 720.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.390 716.000 922.670 720.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.110 716.000 937.390 720.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.830 716.000 952.110 720.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.550 716.000 966.830 720.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.270 716.000 981.550 720.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 716.000 186.670 720.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.990 716.000 996.270 720.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1010.710 716.000 1010.990 720.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.430 716.000 1025.710 720.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1040.150 716.000 1040.430 720.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.870 716.000 1055.150 720.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.590 716.000 1069.870 720.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.310 716.000 1084.590 720.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.030 716.000 1099.310 720.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.750 716.000 1114.030 720.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1128.470 716.000 1128.750 720.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 716.000 201.390 720.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.190 716.000 1143.470 720.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1157.910 716.000 1158.190 720.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.630 716.000 1172.910 720.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1187.350 716.000 1187.630 720.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.070 716.000 1202.350 720.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1216.790 716.000 1217.070 720.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.510 716.000 1231.790 720.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.230 716.000 1246.510 720.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.950 716.000 1261.230 720.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1275.670 716.000 1275.950 720.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 716.000 216.110 720.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1290.390 716.000 1290.670 720.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1305.110 716.000 1305.390 720.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1319.830 716.000 1320.110 720.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1334.550 716.000 1334.830 720.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1349.270 716.000 1349.550 720.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.990 716.000 1364.270 720.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1378.710 716.000 1378.990 720.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1393.430 716.000 1393.710 720.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1408.150 716.000 1408.430 720.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1422.870 716.000 1423.150 720.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 716.000 230.830 720.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1437.590 716.000 1437.870 720.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1452.310 716.000 1452.590 720.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.030 716.000 1467.310 720.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.750 716.000 1482.030 720.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1496.470 716.000 1496.750 720.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1511.190 716.000 1511.470 720.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1525.910 716.000 1526.190 720.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1540.630 716.000 1540.910 720.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.350 716.000 1555.630 720.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1570.070 716.000 1570.350 720.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 716.000 245.550 720.000 ;
    END
  END la_oenb[9]
  PIN la_output[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.470 716.000 116.750 720.000 ;
    END
  END la_output[0]
  PIN la_output[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.470 716.000 1588.750 720.000 ;
    END
  END la_output[100]
  PIN la_output[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1603.190 716.000 1603.470 720.000 ;
    END
  END la_output[101]
  PIN la_output[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1617.910 716.000 1618.190 720.000 ;
    END
  END la_output[102]
  PIN la_output[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.630 716.000 1632.910 720.000 ;
    END
  END la_output[103]
  PIN la_output[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1647.350 716.000 1647.630 720.000 ;
    END
  END la_output[104]
  PIN la_output[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.070 716.000 1662.350 720.000 ;
    END
  END la_output[105]
  PIN la_output[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1676.790 716.000 1677.070 720.000 ;
    END
  END la_output[106]
  PIN la_output[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1691.510 716.000 1691.790 720.000 ;
    END
  END la_output[107]
  PIN la_output[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1706.230 716.000 1706.510 720.000 ;
    END
  END la_output[108]
  PIN la_output[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1720.950 716.000 1721.230 720.000 ;
    END
  END la_output[109]
  PIN la_output[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.670 716.000 263.950 720.000 ;
    END
  END la_output[10]
  PIN la_output[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1735.670 716.000 1735.950 720.000 ;
    END
  END la_output[110]
  PIN la_output[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1750.390 716.000 1750.670 720.000 ;
    END
  END la_output[111]
  PIN la_output[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1765.110 716.000 1765.390 720.000 ;
    END
  END la_output[112]
  PIN la_output[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1779.830 716.000 1780.110 720.000 ;
    END
  END la_output[113]
  PIN la_output[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1794.550 716.000 1794.830 720.000 ;
    END
  END la_output[114]
  PIN la_output[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1809.270 716.000 1809.550 720.000 ;
    END
  END la_output[115]
  PIN la_output[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1823.990 716.000 1824.270 720.000 ;
    END
  END la_output[116]
  PIN la_output[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1838.710 716.000 1838.990 720.000 ;
    END
  END la_output[117]
  PIN la_output[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1853.430 716.000 1853.710 720.000 ;
    END
  END la_output[118]
  PIN la_output[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1868.150 716.000 1868.430 720.000 ;
    END
  END la_output[119]
  PIN la_output[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.390 716.000 278.670 720.000 ;
    END
  END la_output[11]
  PIN la_output[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.870 716.000 1883.150 720.000 ;
    END
  END la_output[120]
  PIN la_output[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1897.590 716.000 1897.870 720.000 ;
    END
  END la_output[121]
  PIN la_output[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1912.310 716.000 1912.590 720.000 ;
    END
  END la_output[122]
  PIN la_output[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1927.030 716.000 1927.310 720.000 ;
    END
  END la_output[123]
  PIN la_output[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.750 716.000 1942.030 720.000 ;
    END
  END la_output[124]
  PIN la_output[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1956.470 716.000 1956.750 720.000 ;
    END
  END la_output[125]
  PIN la_output[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.190 716.000 1971.470 720.000 ;
    END
  END la_output[126]
  PIN la_output[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1985.910 716.000 1986.190 720.000 ;
    END
  END la_output[127]
  PIN la_output[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 716.000 293.390 720.000 ;
    END
  END la_output[12]
  PIN la_output[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.830 716.000 308.110 720.000 ;
    END
  END la_output[13]
  PIN la_output[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 716.000 322.830 720.000 ;
    END
  END la_output[14]
  PIN la_output[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 716.000 337.550 720.000 ;
    END
  END la_output[15]
  PIN la_output[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 716.000 352.270 720.000 ;
    END
  END la_output[16]
  PIN la_output[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 716.000 366.990 720.000 ;
    END
  END la_output[17]
  PIN la_output[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.430 716.000 381.710 720.000 ;
    END
  END la_output[18]
  PIN la_output[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.150 716.000 396.430 720.000 ;
    END
  END la_output[19]
  PIN la_output[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 716.000 131.470 720.000 ;
    END
  END la_output[1]
  PIN la_output[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 716.000 411.150 720.000 ;
    END
  END la_output[20]
  PIN la_output[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 716.000 425.870 720.000 ;
    END
  END la_output[21]
  PIN la_output[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 716.000 440.590 720.000 ;
    END
  END la_output[22]
  PIN la_output[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 716.000 455.310 720.000 ;
    END
  END la_output[23]
  PIN la_output[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 716.000 470.030 720.000 ;
    END
  END la_output[24]
  PIN la_output[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 716.000 484.750 720.000 ;
    END
  END la_output[25]
  PIN la_output[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 716.000 499.470 720.000 ;
    END
  END la_output[26]
  PIN la_output[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 716.000 514.190 720.000 ;
    END
  END la_output[27]
  PIN la_output[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 716.000 528.910 720.000 ;
    END
  END la_output[28]
  PIN la_output[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 543.350 716.000 543.630 720.000 ;
    END
  END la_output[29]
  PIN la_output[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 716.000 146.190 720.000 ;
    END
  END la_output[2]
  PIN la_output[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.070 716.000 558.350 720.000 ;
    END
  END la_output[30]
  PIN la_output[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 716.000 573.070 720.000 ;
    END
  END la_output[31]
  PIN la_output[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.510 716.000 587.790 720.000 ;
    END
  END la_output[32]
  PIN la_output[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 716.000 602.510 720.000 ;
    END
  END la_output[33]
  PIN la_output[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.950 716.000 617.230 720.000 ;
    END
  END la_output[34]
  PIN la_output[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.670 716.000 631.950 720.000 ;
    END
  END la_output[35]
  PIN la_output[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.390 716.000 646.670 720.000 ;
    END
  END la_output[36]
  PIN la_output[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.110 716.000 661.390 720.000 ;
    END
  END la_output[37]
  PIN la_output[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.830 716.000 676.110 720.000 ;
    END
  END la_output[38]
  PIN la_output[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.550 716.000 690.830 720.000 ;
    END
  END la_output[39]
  PIN la_output[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 716.000 160.910 720.000 ;
    END
  END la_output[3]
  PIN la_output[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 716.000 705.550 720.000 ;
    END
  END la_output[40]
  PIN la_output[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.990 716.000 720.270 720.000 ;
    END
  END la_output[41]
  PIN la_output[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.710 716.000 734.990 720.000 ;
    END
  END la_output[42]
  PIN la_output[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 716.000 749.710 720.000 ;
    END
  END la_output[43]
  PIN la_output[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.150 716.000 764.430 720.000 ;
    END
  END la_output[44]
  PIN la_output[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.870 716.000 779.150 720.000 ;
    END
  END la_output[45]
  PIN la_output[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 716.000 793.870 720.000 ;
    END
  END la_output[46]
  PIN la_output[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 808.310 716.000 808.590 720.000 ;
    END
  END la_output[47]
  PIN la_output[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.030 716.000 823.310 720.000 ;
    END
  END la_output[48]
  PIN la_output[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.750 716.000 838.030 720.000 ;
    END
  END la_output[49]
  PIN la_output[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 716.000 175.630 720.000 ;
    END
  END la_output[4]
  PIN la_output[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.470 716.000 852.750 720.000 ;
    END
  END la_output[50]
  PIN la_output[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 867.190 716.000 867.470 720.000 ;
    END
  END la_output[51]
  PIN la_output[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.910 716.000 882.190 720.000 ;
    END
  END la_output[52]
  PIN la_output[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.630 716.000 896.910 720.000 ;
    END
  END la_output[53]
  PIN la_output[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.350 716.000 911.630 720.000 ;
    END
  END la_output[54]
  PIN la_output[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.070 716.000 926.350 720.000 ;
    END
  END la_output[55]
  PIN la_output[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.790 716.000 941.070 720.000 ;
    END
  END la_output[56]
  PIN la_output[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 955.510 716.000 955.790 720.000 ;
    END
  END la_output[57]
  PIN la_output[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.230 716.000 970.510 720.000 ;
    END
  END la_output[58]
  PIN la_output[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.950 716.000 985.230 720.000 ;
    END
  END la_output[59]
  PIN la_output[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 716.000 190.350 720.000 ;
    END
  END la_output[5]
  PIN la_output[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.670 716.000 999.950 720.000 ;
    END
  END la_output[60]
  PIN la_output[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.390 716.000 1014.670 720.000 ;
    END
  END la_output[61]
  PIN la_output[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.110 716.000 1029.390 720.000 ;
    END
  END la_output[62]
  PIN la_output[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1043.830 716.000 1044.110 720.000 ;
    END
  END la_output[63]
  PIN la_output[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.550 716.000 1058.830 720.000 ;
    END
  END la_output[64]
  PIN la_output[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1073.270 716.000 1073.550 720.000 ;
    END
  END la_output[65]
  PIN la_output[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.990 716.000 1088.270 720.000 ;
    END
  END la_output[66]
  PIN la_output[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.710 716.000 1102.990 720.000 ;
    END
  END la_output[67]
  PIN la_output[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.430 716.000 1117.710 720.000 ;
    END
  END la_output[68]
  PIN la_output[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1132.150 716.000 1132.430 720.000 ;
    END
  END la_output[69]
  PIN la_output[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.790 716.000 205.070 720.000 ;
    END
  END la_output[6]
  PIN la_output[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1146.870 716.000 1147.150 720.000 ;
    END
  END la_output[70]
  PIN la_output[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1161.590 716.000 1161.870 720.000 ;
    END
  END la_output[71]
  PIN la_output[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.310 716.000 1176.590 720.000 ;
    END
  END la_output[72]
  PIN la_output[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.030 716.000 1191.310 720.000 ;
    END
  END la_output[73]
  PIN la_output[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.750 716.000 1206.030 720.000 ;
    END
  END la_output[74]
  PIN la_output[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.470 716.000 1220.750 720.000 ;
    END
  END la_output[75]
  PIN la_output[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1235.190 716.000 1235.470 720.000 ;
    END
  END la_output[76]
  PIN la_output[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.910 716.000 1250.190 720.000 ;
    END
  END la_output[77]
  PIN la_output[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1264.630 716.000 1264.910 720.000 ;
    END
  END la_output[78]
  PIN la_output[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.350 716.000 1279.630 720.000 ;
    END
  END la_output[79]
  PIN la_output[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 716.000 219.790 720.000 ;
    END
  END la_output[7]
  PIN la_output[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1294.070 716.000 1294.350 720.000 ;
    END
  END la_output[80]
  PIN la_output[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.790 716.000 1309.070 720.000 ;
    END
  END la_output[81]
  PIN la_output[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.510 716.000 1323.790 720.000 ;
    END
  END la_output[82]
  PIN la_output[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.230 716.000 1338.510 720.000 ;
    END
  END la_output[83]
  PIN la_output[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.950 716.000 1353.230 720.000 ;
    END
  END la_output[84]
  PIN la_output[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.670 716.000 1367.950 720.000 ;
    END
  END la_output[85]
  PIN la_output[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1382.390 716.000 1382.670 720.000 ;
    END
  END la_output[86]
  PIN la_output[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.110 716.000 1397.390 720.000 ;
    END
  END la_output[87]
  PIN la_output[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1411.830 716.000 1412.110 720.000 ;
    END
  END la_output[88]
  PIN la_output[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.550 716.000 1426.830 720.000 ;
    END
  END la_output[89]
  PIN la_output[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 716.000 234.510 720.000 ;
    END
  END la_output[8]
  PIN la_output[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1441.270 716.000 1441.550 720.000 ;
    END
  END la_output[90]
  PIN la_output[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.990 716.000 1456.270 720.000 ;
    END
  END la_output[91]
  PIN la_output[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1470.710 716.000 1470.990 720.000 ;
    END
  END la_output[92]
  PIN la_output[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1485.430 716.000 1485.710 720.000 ;
    END
  END la_output[93]
  PIN la_output[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.150 716.000 1500.430 720.000 ;
    END
  END la_output[94]
  PIN la_output[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1514.870 716.000 1515.150 720.000 ;
    END
  END la_output[95]
  PIN la_output[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1529.590 716.000 1529.870 720.000 ;
    END
  END la_output[96]
  PIN la_output[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1544.310 716.000 1544.590 720.000 ;
    END
  END la_output[97]
  PIN la_output[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1559.030 716.000 1559.310 720.000 ;
    END
  END la_output[98]
  PIN la_output[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1573.750 716.000 1574.030 720.000 ;
    END
  END la_output[99]
  PIN la_output[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 716.000 249.230 720.000 ;
    END
  END la_output[9]
  PIN mprj_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1989.590 716.000 1989.870 720.000 ;
    END
  END mprj_ack_i
  PIN mprj_adr_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2007.990 716.000 2008.270 720.000 ;
    END
  END mprj_adr_o[0]
  PIN mprj_adr_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2133.110 716.000 2133.390 720.000 ;
    END
  END mprj_adr_o[10]
  PIN mprj_adr_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2144.150 716.000 2144.430 720.000 ;
    END
  END mprj_adr_o[11]
  PIN mprj_adr_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2155.190 716.000 2155.470 720.000 ;
    END
  END mprj_adr_o[12]
  PIN mprj_adr_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2166.230 716.000 2166.510 720.000 ;
    END
  END mprj_adr_o[13]
  PIN mprj_adr_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.270 716.000 2177.550 720.000 ;
    END
  END mprj_adr_o[14]
  PIN mprj_adr_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2188.310 716.000 2188.590 720.000 ;
    END
  END mprj_adr_o[15]
  PIN mprj_adr_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2199.350 716.000 2199.630 720.000 ;
    END
  END mprj_adr_o[16]
  PIN mprj_adr_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2210.390 716.000 2210.670 720.000 ;
    END
  END mprj_adr_o[17]
  PIN mprj_adr_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2221.430 716.000 2221.710 720.000 ;
    END
  END mprj_adr_o[18]
  PIN mprj_adr_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2232.470 716.000 2232.750 720.000 ;
    END
  END mprj_adr_o[19]
  PIN mprj_adr_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2022.710 716.000 2022.990 720.000 ;
    END
  END mprj_adr_o[1]
  PIN mprj_adr_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2243.510 716.000 2243.790 720.000 ;
    END
  END mprj_adr_o[20]
  PIN mprj_adr_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2254.550 716.000 2254.830 720.000 ;
    END
  END mprj_adr_o[21]
  PIN mprj_adr_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2265.590 716.000 2265.870 720.000 ;
    END
  END mprj_adr_o[22]
  PIN mprj_adr_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2276.630 716.000 2276.910 720.000 ;
    END
  END mprj_adr_o[23]
  PIN mprj_adr_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2287.670 716.000 2287.950 720.000 ;
    END
  END mprj_adr_o[24]
  PIN mprj_adr_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2298.710 716.000 2298.990 720.000 ;
    END
  END mprj_adr_o[25]
  PIN mprj_adr_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2309.750 716.000 2310.030 720.000 ;
    END
  END mprj_adr_o[26]
  PIN mprj_adr_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2320.790 716.000 2321.070 720.000 ;
    END
  END mprj_adr_o[27]
  PIN mprj_adr_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.830 716.000 2332.110 720.000 ;
    END
  END mprj_adr_o[28]
  PIN mprj_adr_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2342.870 716.000 2343.150 720.000 ;
    END
  END mprj_adr_o[29]
  PIN mprj_adr_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2037.430 716.000 2037.710 720.000 ;
    END
  END mprj_adr_o[2]
  PIN mprj_adr_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2353.910 716.000 2354.190 720.000 ;
    END
  END mprj_adr_o[30]
  PIN mprj_adr_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2364.950 716.000 2365.230 720.000 ;
    END
  END mprj_adr_o[31]
  PIN mprj_adr_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2052.150 716.000 2052.430 720.000 ;
    END
  END mprj_adr_o[3]
  PIN mprj_adr_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2066.870 716.000 2067.150 720.000 ;
    END
  END mprj_adr_o[4]
  PIN mprj_adr_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.910 716.000 2078.190 720.000 ;
    END
  END mprj_adr_o[5]
  PIN mprj_adr_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2088.950 716.000 2089.230 720.000 ;
    END
  END mprj_adr_o[6]
  PIN mprj_adr_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2099.990 716.000 2100.270 720.000 ;
    END
  END mprj_adr_o[7]
  PIN mprj_adr_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2111.030 716.000 2111.310 720.000 ;
    END
  END mprj_adr_o[8]
  PIN mprj_adr_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2122.070 716.000 2122.350 720.000 ;
    END
  END mprj_adr_o[9]
  PIN mprj_cyc_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1993.270 716.000 1993.550 720.000 ;
    END
  END mprj_cyc_o
  PIN mprj_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2011.670 716.000 2011.950 720.000 ;
    END
  END mprj_dat_i[0]
  PIN mprj_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.790 716.000 2137.070 720.000 ;
    END
  END mprj_dat_i[10]
  PIN mprj_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2147.830 716.000 2148.110 720.000 ;
    END
  END mprj_dat_i[11]
  PIN mprj_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2158.870 716.000 2159.150 720.000 ;
    END
  END mprj_dat_i[12]
  PIN mprj_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2169.910 716.000 2170.190 720.000 ;
    END
  END mprj_dat_i[13]
  PIN mprj_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2180.950 716.000 2181.230 720.000 ;
    END
  END mprj_dat_i[14]
  PIN mprj_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2191.990 716.000 2192.270 720.000 ;
    END
  END mprj_dat_i[15]
  PIN mprj_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2203.030 716.000 2203.310 720.000 ;
    END
  END mprj_dat_i[16]
  PIN mprj_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2214.070 716.000 2214.350 720.000 ;
    END
  END mprj_dat_i[17]
  PIN mprj_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2225.110 716.000 2225.390 720.000 ;
    END
  END mprj_dat_i[18]
  PIN mprj_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2236.150 716.000 2236.430 720.000 ;
    END
  END mprj_dat_i[19]
  PIN mprj_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2026.390 716.000 2026.670 720.000 ;
    END
  END mprj_dat_i[1]
  PIN mprj_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2247.190 716.000 2247.470 720.000 ;
    END
  END mprj_dat_i[20]
  PIN mprj_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2258.230 716.000 2258.510 720.000 ;
    END
  END mprj_dat_i[21]
  PIN mprj_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2269.270 716.000 2269.550 720.000 ;
    END
  END mprj_dat_i[22]
  PIN mprj_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2280.310 716.000 2280.590 720.000 ;
    END
  END mprj_dat_i[23]
  PIN mprj_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2291.350 716.000 2291.630 720.000 ;
    END
  END mprj_dat_i[24]
  PIN mprj_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2302.390 716.000 2302.670 720.000 ;
    END
  END mprj_dat_i[25]
  PIN mprj_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2313.430 716.000 2313.710 720.000 ;
    END
  END mprj_dat_i[26]
  PIN mprj_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2324.470 716.000 2324.750 720.000 ;
    END
  END mprj_dat_i[27]
  PIN mprj_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2335.510 716.000 2335.790 720.000 ;
    END
  END mprj_dat_i[28]
  PIN mprj_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2346.550 716.000 2346.830 720.000 ;
    END
  END mprj_dat_i[29]
  PIN mprj_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.110 716.000 2041.390 720.000 ;
    END
  END mprj_dat_i[2]
  PIN mprj_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2357.590 716.000 2357.870 720.000 ;
    END
  END mprj_dat_i[30]
  PIN mprj_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2368.630 716.000 2368.910 720.000 ;
    END
  END mprj_dat_i[31]
  PIN mprj_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2055.830 716.000 2056.110 720.000 ;
    END
  END mprj_dat_i[3]
  PIN mprj_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2070.550 716.000 2070.830 720.000 ;
    END
  END mprj_dat_i[4]
  PIN mprj_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2081.590 716.000 2081.870 720.000 ;
    END
  END mprj_dat_i[5]
  PIN mprj_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2092.630 716.000 2092.910 720.000 ;
    END
  END mprj_dat_i[6]
  PIN mprj_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2103.670 716.000 2103.950 720.000 ;
    END
  END mprj_dat_i[7]
  PIN mprj_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2114.710 716.000 2114.990 720.000 ;
    END
  END mprj_dat_i[8]
  PIN mprj_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2125.750 716.000 2126.030 720.000 ;
    END
  END mprj_dat_i[9]
  PIN mprj_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2015.350 716.000 2015.630 720.000 ;
    END
  END mprj_dat_o[0]
  PIN mprj_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2140.470 716.000 2140.750 720.000 ;
    END
  END mprj_dat_o[10]
  PIN mprj_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2151.510 716.000 2151.790 720.000 ;
    END
  END mprj_dat_o[11]
  PIN mprj_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2162.550 716.000 2162.830 720.000 ;
    END
  END mprj_dat_o[12]
  PIN mprj_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2173.590 716.000 2173.870 720.000 ;
    END
  END mprj_dat_o[13]
  PIN mprj_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2184.630 716.000 2184.910 720.000 ;
    END
  END mprj_dat_o[14]
  PIN mprj_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.670 716.000 2195.950 720.000 ;
    END
  END mprj_dat_o[15]
  PIN mprj_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2206.710 716.000 2206.990 720.000 ;
    END
  END mprj_dat_o[16]
  PIN mprj_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2217.750 716.000 2218.030 720.000 ;
    END
  END mprj_dat_o[17]
  PIN mprj_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2228.790 716.000 2229.070 720.000 ;
    END
  END mprj_dat_o[18]
  PIN mprj_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2239.830 716.000 2240.110 720.000 ;
    END
  END mprj_dat_o[19]
  PIN mprj_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.070 716.000 2030.350 720.000 ;
    END
  END mprj_dat_o[1]
  PIN mprj_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2250.870 716.000 2251.150 720.000 ;
    END
  END mprj_dat_o[20]
  PIN mprj_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2261.910 716.000 2262.190 720.000 ;
    END
  END mprj_dat_o[21]
  PIN mprj_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2272.950 716.000 2273.230 720.000 ;
    END
  END mprj_dat_o[22]
  PIN mprj_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2283.990 716.000 2284.270 720.000 ;
    END
  END mprj_dat_o[23]
  PIN mprj_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.030 716.000 2295.310 720.000 ;
    END
  END mprj_dat_o[24]
  PIN mprj_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2306.070 716.000 2306.350 720.000 ;
    END
  END mprj_dat_o[25]
  PIN mprj_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2317.110 716.000 2317.390 720.000 ;
    END
  END mprj_dat_o[26]
  PIN mprj_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.150 716.000 2328.430 720.000 ;
    END
  END mprj_dat_o[27]
  PIN mprj_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2339.190 716.000 2339.470 720.000 ;
    END
  END mprj_dat_o[28]
  PIN mprj_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2350.230 716.000 2350.510 720.000 ;
    END
  END mprj_dat_o[29]
  PIN mprj_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2044.790 716.000 2045.070 720.000 ;
    END
  END mprj_dat_o[2]
  PIN mprj_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.270 716.000 2361.550 720.000 ;
    END
  END mprj_dat_o[30]
  PIN mprj_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2372.310 716.000 2372.590 720.000 ;
    END
  END mprj_dat_o[31]
  PIN mprj_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.510 716.000 2059.790 720.000 ;
    END
  END mprj_dat_o[3]
  PIN mprj_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2074.230 716.000 2074.510 720.000 ;
    END
  END mprj_dat_o[4]
  PIN mprj_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2085.270 716.000 2085.550 720.000 ;
    END
  END mprj_dat_o[5]
  PIN mprj_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2096.310 716.000 2096.590 720.000 ;
    END
  END mprj_dat_o[6]
  PIN mprj_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2107.350 716.000 2107.630 720.000 ;
    END
  END mprj_dat_o[7]
  PIN mprj_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.390 716.000 2118.670 720.000 ;
    END
  END mprj_dat_o[8]
  PIN mprj_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2129.430 716.000 2129.710 720.000 ;
    END
  END mprj_dat_o[9]
  PIN mprj_sel_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.030 716.000 2019.310 720.000 ;
    END
  END mprj_sel_o[0]
  PIN mprj_sel_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2033.750 716.000 2034.030 720.000 ;
    END
  END mprj_sel_o[1]
  PIN mprj_sel_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.470 716.000 2048.750 720.000 ;
    END
  END mprj_sel_o[2]
  PIN mprj_sel_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2063.190 716.000 2063.470 720.000 ;
    END
  END mprj_sel_o[3]
  PIN mprj_stb_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1996.950 716.000 1997.230 720.000 ;
    END
  END mprj_stb_o
  PIN mprj_wb_iena
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.630 716.000 2000.910 720.000 ;
    END
  END mprj_wb_iena
  PIN mprj_we_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2004.310 716.000 2004.590 720.000 ;
    END
  END mprj_we_o
  PIN qspi_enabled
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 206.760 2500.000 207.360 ;
    END
  END qspi_enabled
  PIN ser_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 168.680 2500.000 169.280 ;
    END
  END ser_rx
  PIN ser_tx
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 178.200 2500.000 178.800 ;
    END
  END ser_tx
  PIN spi_csb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 149.640 2500.000 150.240 ;
    END
  END spi_csb
  PIN spi_enabled
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 187.720 2500.000 188.320 ;
    END
  END spi_enabled
  PIN spi_sck
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 140.120 2500.000 140.720 ;
    END
  END spi_sck
  PIN spi_sdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 159.160 2500.000 159.760 ;
    END
  END spi_sdi
  PIN spi_sdo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 130.600 2500.000 131.200 ;
    END
  END spi_sdo
  PIN spi_sdoenb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 121.080 2500.000 121.680 ;
    END
  END spi_sdoenb
  PIN tck
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END tck
  PIN tdi
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 0.000 262.570 4.000 ;
    END
  END tdi
  PIN tdo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END tdo
  PIN tdo_paden_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.170 0.000 574.450 4.000 ;
    END
  END tdo_paden_o
  PIN tms
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 0.000 54.650 4.000 ;
    END
  END tms
  PIN trap
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 83.000 2500.000 83.600 ;
    END
  END trap
  PIN trst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 0.000 470.490 4.000 ;
    END
  END trst
  PIN uart_enabled
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2496.000 197.240 2500.000 197.840 ;
    END
  END uart_enabled
  PIN user_irq_ena[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2375.990 716.000 2376.270 720.000 ;
    END
  END user_irq_ena[0]
  PIN user_irq_ena[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2379.670 716.000 2379.950 720.000 ;
    END
  END user_irq_ena[1]
  PIN user_irq_ena[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2383.350 716.000 2383.630 720.000 ;
    END
  END user_irq_ena[2]
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2494.120 707.285 ;
      LAYER met1 ;
        RECT 5.520 2.420 2499.570 718.040 ;
      LAYER met2 ;
        RECT 13.900 715.720 105.150 718.070 ;
        RECT 105.990 715.720 108.830 718.070 ;
        RECT 109.670 715.720 112.510 718.070 ;
        RECT 113.350 715.720 116.190 718.070 ;
        RECT 117.030 715.720 119.870 718.070 ;
        RECT 120.710 715.720 123.550 718.070 ;
        RECT 124.390 715.720 127.230 718.070 ;
        RECT 128.070 715.720 130.910 718.070 ;
        RECT 131.750 715.720 134.590 718.070 ;
        RECT 135.430 715.720 138.270 718.070 ;
        RECT 139.110 715.720 141.950 718.070 ;
        RECT 142.790 715.720 145.630 718.070 ;
        RECT 146.470 715.720 149.310 718.070 ;
        RECT 150.150 715.720 152.990 718.070 ;
        RECT 153.830 715.720 156.670 718.070 ;
        RECT 157.510 715.720 160.350 718.070 ;
        RECT 161.190 715.720 164.030 718.070 ;
        RECT 164.870 715.720 167.710 718.070 ;
        RECT 168.550 715.720 171.390 718.070 ;
        RECT 172.230 715.720 175.070 718.070 ;
        RECT 175.910 715.720 178.750 718.070 ;
        RECT 179.590 715.720 182.430 718.070 ;
        RECT 183.270 715.720 186.110 718.070 ;
        RECT 186.950 715.720 189.790 718.070 ;
        RECT 190.630 715.720 193.470 718.070 ;
        RECT 194.310 715.720 197.150 718.070 ;
        RECT 197.990 715.720 200.830 718.070 ;
        RECT 201.670 715.720 204.510 718.070 ;
        RECT 205.350 715.720 208.190 718.070 ;
        RECT 209.030 715.720 211.870 718.070 ;
        RECT 212.710 715.720 215.550 718.070 ;
        RECT 216.390 715.720 219.230 718.070 ;
        RECT 220.070 715.720 222.910 718.070 ;
        RECT 223.750 715.720 226.590 718.070 ;
        RECT 227.430 715.720 230.270 718.070 ;
        RECT 231.110 715.720 233.950 718.070 ;
        RECT 234.790 715.720 237.630 718.070 ;
        RECT 238.470 715.720 241.310 718.070 ;
        RECT 242.150 715.720 244.990 718.070 ;
        RECT 245.830 715.720 248.670 718.070 ;
        RECT 249.510 715.720 252.350 718.070 ;
        RECT 253.190 715.720 256.030 718.070 ;
        RECT 256.870 715.720 259.710 718.070 ;
        RECT 260.550 715.720 263.390 718.070 ;
        RECT 264.230 715.720 267.070 718.070 ;
        RECT 267.910 715.720 270.750 718.070 ;
        RECT 271.590 715.720 274.430 718.070 ;
        RECT 275.270 715.720 278.110 718.070 ;
        RECT 278.950 715.720 281.790 718.070 ;
        RECT 282.630 715.720 285.470 718.070 ;
        RECT 286.310 715.720 289.150 718.070 ;
        RECT 289.990 715.720 292.830 718.070 ;
        RECT 293.670 715.720 296.510 718.070 ;
        RECT 297.350 715.720 300.190 718.070 ;
        RECT 301.030 715.720 303.870 718.070 ;
        RECT 304.710 715.720 307.550 718.070 ;
        RECT 308.390 715.720 311.230 718.070 ;
        RECT 312.070 715.720 314.910 718.070 ;
        RECT 315.750 715.720 318.590 718.070 ;
        RECT 319.430 715.720 322.270 718.070 ;
        RECT 323.110 715.720 325.950 718.070 ;
        RECT 326.790 715.720 329.630 718.070 ;
        RECT 330.470 715.720 333.310 718.070 ;
        RECT 334.150 715.720 336.990 718.070 ;
        RECT 337.830 715.720 340.670 718.070 ;
        RECT 341.510 715.720 344.350 718.070 ;
        RECT 345.190 715.720 348.030 718.070 ;
        RECT 348.870 715.720 351.710 718.070 ;
        RECT 352.550 715.720 355.390 718.070 ;
        RECT 356.230 715.720 359.070 718.070 ;
        RECT 359.910 715.720 362.750 718.070 ;
        RECT 363.590 715.720 366.430 718.070 ;
        RECT 367.270 715.720 370.110 718.070 ;
        RECT 370.950 715.720 373.790 718.070 ;
        RECT 374.630 715.720 377.470 718.070 ;
        RECT 378.310 715.720 381.150 718.070 ;
        RECT 381.990 715.720 384.830 718.070 ;
        RECT 385.670 715.720 388.510 718.070 ;
        RECT 389.350 715.720 392.190 718.070 ;
        RECT 393.030 715.720 395.870 718.070 ;
        RECT 396.710 715.720 399.550 718.070 ;
        RECT 400.390 715.720 403.230 718.070 ;
        RECT 404.070 715.720 406.910 718.070 ;
        RECT 407.750 715.720 410.590 718.070 ;
        RECT 411.430 715.720 414.270 718.070 ;
        RECT 415.110 715.720 417.950 718.070 ;
        RECT 418.790 715.720 421.630 718.070 ;
        RECT 422.470 715.720 425.310 718.070 ;
        RECT 426.150 715.720 428.990 718.070 ;
        RECT 429.830 715.720 432.670 718.070 ;
        RECT 433.510 715.720 436.350 718.070 ;
        RECT 437.190 715.720 440.030 718.070 ;
        RECT 440.870 715.720 443.710 718.070 ;
        RECT 444.550 715.720 447.390 718.070 ;
        RECT 448.230 715.720 451.070 718.070 ;
        RECT 451.910 715.720 454.750 718.070 ;
        RECT 455.590 715.720 458.430 718.070 ;
        RECT 459.270 715.720 462.110 718.070 ;
        RECT 462.950 715.720 465.790 718.070 ;
        RECT 466.630 715.720 469.470 718.070 ;
        RECT 470.310 715.720 473.150 718.070 ;
        RECT 473.990 715.720 476.830 718.070 ;
        RECT 477.670 715.720 480.510 718.070 ;
        RECT 481.350 715.720 484.190 718.070 ;
        RECT 485.030 715.720 487.870 718.070 ;
        RECT 488.710 715.720 491.550 718.070 ;
        RECT 492.390 715.720 495.230 718.070 ;
        RECT 496.070 715.720 498.910 718.070 ;
        RECT 499.750 715.720 502.590 718.070 ;
        RECT 503.430 715.720 506.270 718.070 ;
        RECT 507.110 715.720 509.950 718.070 ;
        RECT 510.790 715.720 513.630 718.070 ;
        RECT 514.470 715.720 517.310 718.070 ;
        RECT 518.150 715.720 520.990 718.070 ;
        RECT 521.830 715.720 524.670 718.070 ;
        RECT 525.510 715.720 528.350 718.070 ;
        RECT 529.190 715.720 532.030 718.070 ;
        RECT 532.870 715.720 535.710 718.070 ;
        RECT 536.550 715.720 539.390 718.070 ;
        RECT 540.230 715.720 543.070 718.070 ;
        RECT 543.910 715.720 546.750 718.070 ;
        RECT 547.590 715.720 550.430 718.070 ;
        RECT 551.270 715.720 554.110 718.070 ;
        RECT 554.950 715.720 557.790 718.070 ;
        RECT 558.630 715.720 561.470 718.070 ;
        RECT 562.310 715.720 565.150 718.070 ;
        RECT 565.990 715.720 568.830 718.070 ;
        RECT 569.670 715.720 572.510 718.070 ;
        RECT 573.350 715.720 576.190 718.070 ;
        RECT 577.030 715.720 579.870 718.070 ;
        RECT 580.710 715.720 583.550 718.070 ;
        RECT 584.390 715.720 587.230 718.070 ;
        RECT 588.070 715.720 590.910 718.070 ;
        RECT 591.750 715.720 594.590 718.070 ;
        RECT 595.430 715.720 598.270 718.070 ;
        RECT 599.110 715.720 601.950 718.070 ;
        RECT 602.790 715.720 605.630 718.070 ;
        RECT 606.470 715.720 609.310 718.070 ;
        RECT 610.150 715.720 612.990 718.070 ;
        RECT 613.830 715.720 616.670 718.070 ;
        RECT 617.510 715.720 620.350 718.070 ;
        RECT 621.190 715.720 624.030 718.070 ;
        RECT 624.870 715.720 627.710 718.070 ;
        RECT 628.550 715.720 631.390 718.070 ;
        RECT 632.230 715.720 635.070 718.070 ;
        RECT 635.910 715.720 638.750 718.070 ;
        RECT 639.590 715.720 642.430 718.070 ;
        RECT 643.270 715.720 646.110 718.070 ;
        RECT 646.950 715.720 649.790 718.070 ;
        RECT 650.630 715.720 653.470 718.070 ;
        RECT 654.310 715.720 657.150 718.070 ;
        RECT 657.990 715.720 660.830 718.070 ;
        RECT 661.670 715.720 664.510 718.070 ;
        RECT 665.350 715.720 668.190 718.070 ;
        RECT 669.030 715.720 671.870 718.070 ;
        RECT 672.710 715.720 675.550 718.070 ;
        RECT 676.390 715.720 679.230 718.070 ;
        RECT 680.070 715.720 682.910 718.070 ;
        RECT 683.750 715.720 686.590 718.070 ;
        RECT 687.430 715.720 690.270 718.070 ;
        RECT 691.110 715.720 693.950 718.070 ;
        RECT 694.790 715.720 697.630 718.070 ;
        RECT 698.470 715.720 701.310 718.070 ;
        RECT 702.150 715.720 704.990 718.070 ;
        RECT 705.830 715.720 708.670 718.070 ;
        RECT 709.510 715.720 712.350 718.070 ;
        RECT 713.190 715.720 716.030 718.070 ;
        RECT 716.870 715.720 719.710 718.070 ;
        RECT 720.550 715.720 723.390 718.070 ;
        RECT 724.230 715.720 727.070 718.070 ;
        RECT 727.910 715.720 730.750 718.070 ;
        RECT 731.590 715.720 734.430 718.070 ;
        RECT 735.270 715.720 738.110 718.070 ;
        RECT 738.950 715.720 741.790 718.070 ;
        RECT 742.630 715.720 745.470 718.070 ;
        RECT 746.310 715.720 749.150 718.070 ;
        RECT 749.990 715.720 752.830 718.070 ;
        RECT 753.670 715.720 756.510 718.070 ;
        RECT 757.350 715.720 760.190 718.070 ;
        RECT 761.030 715.720 763.870 718.070 ;
        RECT 764.710 715.720 767.550 718.070 ;
        RECT 768.390 715.720 771.230 718.070 ;
        RECT 772.070 715.720 774.910 718.070 ;
        RECT 775.750 715.720 778.590 718.070 ;
        RECT 779.430 715.720 782.270 718.070 ;
        RECT 783.110 715.720 785.950 718.070 ;
        RECT 786.790 715.720 789.630 718.070 ;
        RECT 790.470 715.720 793.310 718.070 ;
        RECT 794.150 715.720 796.990 718.070 ;
        RECT 797.830 715.720 800.670 718.070 ;
        RECT 801.510 715.720 804.350 718.070 ;
        RECT 805.190 715.720 808.030 718.070 ;
        RECT 808.870 715.720 811.710 718.070 ;
        RECT 812.550 715.720 815.390 718.070 ;
        RECT 816.230 715.720 819.070 718.070 ;
        RECT 819.910 715.720 822.750 718.070 ;
        RECT 823.590 715.720 826.430 718.070 ;
        RECT 827.270 715.720 830.110 718.070 ;
        RECT 830.950 715.720 833.790 718.070 ;
        RECT 834.630 715.720 837.470 718.070 ;
        RECT 838.310 715.720 841.150 718.070 ;
        RECT 841.990 715.720 844.830 718.070 ;
        RECT 845.670 715.720 848.510 718.070 ;
        RECT 849.350 715.720 852.190 718.070 ;
        RECT 853.030 715.720 855.870 718.070 ;
        RECT 856.710 715.720 859.550 718.070 ;
        RECT 860.390 715.720 863.230 718.070 ;
        RECT 864.070 715.720 866.910 718.070 ;
        RECT 867.750 715.720 870.590 718.070 ;
        RECT 871.430 715.720 874.270 718.070 ;
        RECT 875.110 715.720 877.950 718.070 ;
        RECT 878.790 715.720 881.630 718.070 ;
        RECT 882.470 715.720 885.310 718.070 ;
        RECT 886.150 715.720 888.990 718.070 ;
        RECT 889.830 715.720 892.670 718.070 ;
        RECT 893.510 715.720 896.350 718.070 ;
        RECT 897.190 715.720 900.030 718.070 ;
        RECT 900.870 715.720 903.710 718.070 ;
        RECT 904.550 715.720 907.390 718.070 ;
        RECT 908.230 715.720 911.070 718.070 ;
        RECT 911.910 715.720 914.750 718.070 ;
        RECT 915.590 715.720 918.430 718.070 ;
        RECT 919.270 715.720 922.110 718.070 ;
        RECT 922.950 715.720 925.790 718.070 ;
        RECT 926.630 715.720 929.470 718.070 ;
        RECT 930.310 715.720 933.150 718.070 ;
        RECT 933.990 715.720 936.830 718.070 ;
        RECT 937.670 715.720 940.510 718.070 ;
        RECT 941.350 715.720 944.190 718.070 ;
        RECT 945.030 715.720 947.870 718.070 ;
        RECT 948.710 715.720 951.550 718.070 ;
        RECT 952.390 715.720 955.230 718.070 ;
        RECT 956.070 715.720 958.910 718.070 ;
        RECT 959.750 715.720 962.590 718.070 ;
        RECT 963.430 715.720 966.270 718.070 ;
        RECT 967.110 715.720 969.950 718.070 ;
        RECT 970.790 715.720 973.630 718.070 ;
        RECT 974.470 715.720 977.310 718.070 ;
        RECT 978.150 715.720 980.990 718.070 ;
        RECT 981.830 715.720 984.670 718.070 ;
        RECT 985.510 715.720 988.350 718.070 ;
        RECT 989.190 715.720 992.030 718.070 ;
        RECT 992.870 715.720 995.710 718.070 ;
        RECT 996.550 715.720 999.390 718.070 ;
        RECT 1000.230 715.720 1003.070 718.070 ;
        RECT 1003.910 715.720 1006.750 718.070 ;
        RECT 1007.590 715.720 1010.430 718.070 ;
        RECT 1011.270 715.720 1014.110 718.070 ;
        RECT 1014.950 715.720 1017.790 718.070 ;
        RECT 1018.630 715.720 1021.470 718.070 ;
        RECT 1022.310 715.720 1025.150 718.070 ;
        RECT 1025.990 715.720 1028.830 718.070 ;
        RECT 1029.670 715.720 1032.510 718.070 ;
        RECT 1033.350 715.720 1036.190 718.070 ;
        RECT 1037.030 715.720 1039.870 718.070 ;
        RECT 1040.710 715.720 1043.550 718.070 ;
        RECT 1044.390 715.720 1047.230 718.070 ;
        RECT 1048.070 715.720 1050.910 718.070 ;
        RECT 1051.750 715.720 1054.590 718.070 ;
        RECT 1055.430 715.720 1058.270 718.070 ;
        RECT 1059.110 715.720 1061.950 718.070 ;
        RECT 1062.790 715.720 1065.630 718.070 ;
        RECT 1066.470 715.720 1069.310 718.070 ;
        RECT 1070.150 715.720 1072.990 718.070 ;
        RECT 1073.830 715.720 1076.670 718.070 ;
        RECT 1077.510 715.720 1080.350 718.070 ;
        RECT 1081.190 715.720 1084.030 718.070 ;
        RECT 1084.870 715.720 1087.710 718.070 ;
        RECT 1088.550 715.720 1091.390 718.070 ;
        RECT 1092.230 715.720 1095.070 718.070 ;
        RECT 1095.910 715.720 1098.750 718.070 ;
        RECT 1099.590 715.720 1102.430 718.070 ;
        RECT 1103.270 715.720 1106.110 718.070 ;
        RECT 1106.950 715.720 1109.790 718.070 ;
        RECT 1110.630 715.720 1113.470 718.070 ;
        RECT 1114.310 715.720 1117.150 718.070 ;
        RECT 1117.990 715.720 1120.830 718.070 ;
        RECT 1121.670 715.720 1124.510 718.070 ;
        RECT 1125.350 715.720 1128.190 718.070 ;
        RECT 1129.030 715.720 1131.870 718.070 ;
        RECT 1132.710 715.720 1135.550 718.070 ;
        RECT 1136.390 715.720 1139.230 718.070 ;
        RECT 1140.070 715.720 1142.910 718.070 ;
        RECT 1143.750 715.720 1146.590 718.070 ;
        RECT 1147.430 715.720 1150.270 718.070 ;
        RECT 1151.110 715.720 1153.950 718.070 ;
        RECT 1154.790 715.720 1157.630 718.070 ;
        RECT 1158.470 715.720 1161.310 718.070 ;
        RECT 1162.150 715.720 1164.990 718.070 ;
        RECT 1165.830 715.720 1168.670 718.070 ;
        RECT 1169.510 715.720 1172.350 718.070 ;
        RECT 1173.190 715.720 1176.030 718.070 ;
        RECT 1176.870 715.720 1179.710 718.070 ;
        RECT 1180.550 715.720 1183.390 718.070 ;
        RECT 1184.230 715.720 1187.070 718.070 ;
        RECT 1187.910 715.720 1190.750 718.070 ;
        RECT 1191.590 715.720 1194.430 718.070 ;
        RECT 1195.270 715.720 1198.110 718.070 ;
        RECT 1198.950 715.720 1201.790 718.070 ;
        RECT 1202.630 715.720 1205.470 718.070 ;
        RECT 1206.310 715.720 1209.150 718.070 ;
        RECT 1209.990 715.720 1212.830 718.070 ;
        RECT 1213.670 715.720 1216.510 718.070 ;
        RECT 1217.350 715.720 1220.190 718.070 ;
        RECT 1221.030 715.720 1223.870 718.070 ;
        RECT 1224.710 715.720 1227.550 718.070 ;
        RECT 1228.390 715.720 1231.230 718.070 ;
        RECT 1232.070 715.720 1234.910 718.070 ;
        RECT 1235.750 715.720 1238.590 718.070 ;
        RECT 1239.430 715.720 1242.270 718.070 ;
        RECT 1243.110 715.720 1245.950 718.070 ;
        RECT 1246.790 715.720 1249.630 718.070 ;
        RECT 1250.470 715.720 1253.310 718.070 ;
        RECT 1254.150 715.720 1256.990 718.070 ;
        RECT 1257.830 715.720 1260.670 718.070 ;
        RECT 1261.510 715.720 1264.350 718.070 ;
        RECT 1265.190 715.720 1268.030 718.070 ;
        RECT 1268.870 715.720 1271.710 718.070 ;
        RECT 1272.550 715.720 1275.390 718.070 ;
        RECT 1276.230 715.720 1279.070 718.070 ;
        RECT 1279.910 715.720 1282.750 718.070 ;
        RECT 1283.590 715.720 1286.430 718.070 ;
        RECT 1287.270 715.720 1290.110 718.070 ;
        RECT 1290.950 715.720 1293.790 718.070 ;
        RECT 1294.630 715.720 1297.470 718.070 ;
        RECT 1298.310 715.720 1301.150 718.070 ;
        RECT 1301.990 715.720 1304.830 718.070 ;
        RECT 1305.670 715.720 1308.510 718.070 ;
        RECT 1309.350 715.720 1312.190 718.070 ;
        RECT 1313.030 715.720 1315.870 718.070 ;
        RECT 1316.710 715.720 1319.550 718.070 ;
        RECT 1320.390 715.720 1323.230 718.070 ;
        RECT 1324.070 715.720 1326.910 718.070 ;
        RECT 1327.750 715.720 1330.590 718.070 ;
        RECT 1331.430 715.720 1334.270 718.070 ;
        RECT 1335.110 715.720 1337.950 718.070 ;
        RECT 1338.790 715.720 1341.630 718.070 ;
        RECT 1342.470 715.720 1345.310 718.070 ;
        RECT 1346.150 715.720 1348.990 718.070 ;
        RECT 1349.830 715.720 1352.670 718.070 ;
        RECT 1353.510 715.720 1356.350 718.070 ;
        RECT 1357.190 715.720 1360.030 718.070 ;
        RECT 1360.870 715.720 1363.710 718.070 ;
        RECT 1364.550 715.720 1367.390 718.070 ;
        RECT 1368.230 715.720 1371.070 718.070 ;
        RECT 1371.910 715.720 1374.750 718.070 ;
        RECT 1375.590 715.720 1378.430 718.070 ;
        RECT 1379.270 715.720 1382.110 718.070 ;
        RECT 1382.950 715.720 1385.790 718.070 ;
        RECT 1386.630 715.720 1389.470 718.070 ;
        RECT 1390.310 715.720 1393.150 718.070 ;
        RECT 1393.990 715.720 1396.830 718.070 ;
        RECT 1397.670 715.720 1400.510 718.070 ;
        RECT 1401.350 715.720 1404.190 718.070 ;
        RECT 1405.030 715.720 1407.870 718.070 ;
        RECT 1408.710 715.720 1411.550 718.070 ;
        RECT 1412.390 715.720 1415.230 718.070 ;
        RECT 1416.070 715.720 1418.910 718.070 ;
        RECT 1419.750 715.720 1422.590 718.070 ;
        RECT 1423.430 715.720 1426.270 718.070 ;
        RECT 1427.110 715.720 1429.950 718.070 ;
        RECT 1430.790 715.720 1433.630 718.070 ;
        RECT 1434.470 715.720 1437.310 718.070 ;
        RECT 1438.150 715.720 1440.990 718.070 ;
        RECT 1441.830 715.720 1444.670 718.070 ;
        RECT 1445.510 715.720 1448.350 718.070 ;
        RECT 1449.190 715.720 1452.030 718.070 ;
        RECT 1452.870 715.720 1455.710 718.070 ;
        RECT 1456.550 715.720 1459.390 718.070 ;
        RECT 1460.230 715.720 1463.070 718.070 ;
        RECT 1463.910 715.720 1466.750 718.070 ;
        RECT 1467.590 715.720 1470.430 718.070 ;
        RECT 1471.270 715.720 1474.110 718.070 ;
        RECT 1474.950 715.720 1477.790 718.070 ;
        RECT 1478.630 715.720 1481.470 718.070 ;
        RECT 1482.310 715.720 1485.150 718.070 ;
        RECT 1485.990 715.720 1488.830 718.070 ;
        RECT 1489.670 715.720 1492.510 718.070 ;
        RECT 1493.350 715.720 1496.190 718.070 ;
        RECT 1497.030 715.720 1499.870 718.070 ;
        RECT 1500.710 715.720 1503.550 718.070 ;
        RECT 1504.390 715.720 1507.230 718.070 ;
        RECT 1508.070 715.720 1510.910 718.070 ;
        RECT 1511.750 715.720 1514.590 718.070 ;
        RECT 1515.430 715.720 1518.270 718.070 ;
        RECT 1519.110 715.720 1521.950 718.070 ;
        RECT 1522.790 715.720 1525.630 718.070 ;
        RECT 1526.470 715.720 1529.310 718.070 ;
        RECT 1530.150 715.720 1532.990 718.070 ;
        RECT 1533.830 715.720 1536.670 718.070 ;
        RECT 1537.510 715.720 1540.350 718.070 ;
        RECT 1541.190 715.720 1544.030 718.070 ;
        RECT 1544.870 715.720 1547.710 718.070 ;
        RECT 1548.550 715.720 1551.390 718.070 ;
        RECT 1552.230 715.720 1555.070 718.070 ;
        RECT 1555.910 715.720 1558.750 718.070 ;
        RECT 1559.590 715.720 1562.430 718.070 ;
        RECT 1563.270 715.720 1566.110 718.070 ;
        RECT 1566.950 715.720 1569.790 718.070 ;
        RECT 1570.630 715.720 1573.470 718.070 ;
        RECT 1574.310 715.720 1577.150 718.070 ;
        RECT 1577.990 715.720 1580.830 718.070 ;
        RECT 1581.670 715.720 1584.510 718.070 ;
        RECT 1585.350 715.720 1588.190 718.070 ;
        RECT 1589.030 715.720 1591.870 718.070 ;
        RECT 1592.710 715.720 1595.550 718.070 ;
        RECT 1596.390 715.720 1599.230 718.070 ;
        RECT 1600.070 715.720 1602.910 718.070 ;
        RECT 1603.750 715.720 1606.590 718.070 ;
        RECT 1607.430 715.720 1610.270 718.070 ;
        RECT 1611.110 715.720 1613.950 718.070 ;
        RECT 1614.790 715.720 1617.630 718.070 ;
        RECT 1618.470 715.720 1621.310 718.070 ;
        RECT 1622.150 715.720 1624.990 718.070 ;
        RECT 1625.830 715.720 1628.670 718.070 ;
        RECT 1629.510 715.720 1632.350 718.070 ;
        RECT 1633.190 715.720 1636.030 718.070 ;
        RECT 1636.870 715.720 1639.710 718.070 ;
        RECT 1640.550 715.720 1643.390 718.070 ;
        RECT 1644.230 715.720 1647.070 718.070 ;
        RECT 1647.910 715.720 1650.750 718.070 ;
        RECT 1651.590 715.720 1654.430 718.070 ;
        RECT 1655.270 715.720 1658.110 718.070 ;
        RECT 1658.950 715.720 1661.790 718.070 ;
        RECT 1662.630 715.720 1665.470 718.070 ;
        RECT 1666.310 715.720 1669.150 718.070 ;
        RECT 1669.990 715.720 1672.830 718.070 ;
        RECT 1673.670 715.720 1676.510 718.070 ;
        RECT 1677.350 715.720 1680.190 718.070 ;
        RECT 1681.030 715.720 1683.870 718.070 ;
        RECT 1684.710 715.720 1687.550 718.070 ;
        RECT 1688.390 715.720 1691.230 718.070 ;
        RECT 1692.070 715.720 1694.910 718.070 ;
        RECT 1695.750 715.720 1698.590 718.070 ;
        RECT 1699.430 715.720 1702.270 718.070 ;
        RECT 1703.110 715.720 1705.950 718.070 ;
        RECT 1706.790 715.720 1709.630 718.070 ;
        RECT 1710.470 715.720 1713.310 718.070 ;
        RECT 1714.150 715.720 1716.990 718.070 ;
        RECT 1717.830 715.720 1720.670 718.070 ;
        RECT 1721.510 715.720 1724.350 718.070 ;
        RECT 1725.190 715.720 1728.030 718.070 ;
        RECT 1728.870 715.720 1731.710 718.070 ;
        RECT 1732.550 715.720 1735.390 718.070 ;
        RECT 1736.230 715.720 1739.070 718.070 ;
        RECT 1739.910 715.720 1742.750 718.070 ;
        RECT 1743.590 715.720 1746.430 718.070 ;
        RECT 1747.270 715.720 1750.110 718.070 ;
        RECT 1750.950 715.720 1753.790 718.070 ;
        RECT 1754.630 715.720 1757.470 718.070 ;
        RECT 1758.310 715.720 1761.150 718.070 ;
        RECT 1761.990 715.720 1764.830 718.070 ;
        RECT 1765.670 715.720 1768.510 718.070 ;
        RECT 1769.350 715.720 1772.190 718.070 ;
        RECT 1773.030 715.720 1775.870 718.070 ;
        RECT 1776.710 715.720 1779.550 718.070 ;
        RECT 1780.390 715.720 1783.230 718.070 ;
        RECT 1784.070 715.720 1786.910 718.070 ;
        RECT 1787.750 715.720 1790.590 718.070 ;
        RECT 1791.430 715.720 1794.270 718.070 ;
        RECT 1795.110 715.720 1797.950 718.070 ;
        RECT 1798.790 715.720 1801.630 718.070 ;
        RECT 1802.470 715.720 1805.310 718.070 ;
        RECT 1806.150 715.720 1808.990 718.070 ;
        RECT 1809.830 715.720 1812.670 718.070 ;
        RECT 1813.510 715.720 1816.350 718.070 ;
        RECT 1817.190 715.720 1820.030 718.070 ;
        RECT 1820.870 715.720 1823.710 718.070 ;
        RECT 1824.550 715.720 1827.390 718.070 ;
        RECT 1828.230 715.720 1831.070 718.070 ;
        RECT 1831.910 715.720 1834.750 718.070 ;
        RECT 1835.590 715.720 1838.430 718.070 ;
        RECT 1839.270 715.720 1842.110 718.070 ;
        RECT 1842.950 715.720 1845.790 718.070 ;
        RECT 1846.630 715.720 1849.470 718.070 ;
        RECT 1850.310 715.720 1853.150 718.070 ;
        RECT 1853.990 715.720 1856.830 718.070 ;
        RECT 1857.670 715.720 1860.510 718.070 ;
        RECT 1861.350 715.720 1864.190 718.070 ;
        RECT 1865.030 715.720 1867.870 718.070 ;
        RECT 1868.710 715.720 1871.550 718.070 ;
        RECT 1872.390 715.720 1875.230 718.070 ;
        RECT 1876.070 715.720 1878.910 718.070 ;
        RECT 1879.750 715.720 1882.590 718.070 ;
        RECT 1883.430 715.720 1886.270 718.070 ;
        RECT 1887.110 715.720 1889.950 718.070 ;
        RECT 1890.790 715.720 1893.630 718.070 ;
        RECT 1894.470 715.720 1897.310 718.070 ;
        RECT 1898.150 715.720 1900.990 718.070 ;
        RECT 1901.830 715.720 1904.670 718.070 ;
        RECT 1905.510 715.720 1908.350 718.070 ;
        RECT 1909.190 715.720 1912.030 718.070 ;
        RECT 1912.870 715.720 1915.710 718.070 ;
        RECT 1916.550 715.720 1919.390 718.070 ;
        RECT 1920.230 715.720 1923.070 718.070 ;
        RECT 1923.910 715.720 1926.750 718.070 ;
        RECT 1927.590 715.720 1930.430 718.070 ;
        RECT 1931.270 715.720 1934.110 718.070 ;
        RECT 1934.950 715.720 1937.790 718.070 ;
        RECT 1938.630 715.720 1941.470 718.070 ;
        RECT 1942.310 715.720 1945.150 718.070 ;
        RECT 1945.990 715.720 1948.830 718.070 ;
        RECT 1949.670 715.720 1952.510 718.070 ;
        RECT 1953.350 715.720 1956.190 718.070 ;
        RECT 1957.030 715.720 1959.870 718.070 ;
        RECT 1960.710 715.720 1963.550 718.070 ;
        RECT 1964.390 715.720 1967.230 718.070 ;
        RECT 1968.070 715.720 1970.910 718.070 ;
        RECT 1971.750 715.720 1974.590 718.070 ;
        RECT 1975.430 715.720 1978.270 718.070 ;
        RECT 1979.110 715.720 1981.950 718.070 ;
        RECT 1982.790 715.720 1985.630 718.070 ;
        RECT 1986.470 715.720 1989.310 718.070 ;
        RECT 1990.150 715.720 1992.990 718.070 ;
        RECT 1993.830 715.720 1996.670 718.070 ;
        RECT 1997.510 715.720 2000.350 718.070 ;
        RECT 2001.190 715.720 2004.030 718.070 ;
        RECT 2004.870 715.720 2007.710 718.070 ;
        RECT 2008.550 715.720 2011.390 718.070 ;
        RECT 2012.230 715.720 2015.070 718.070 ;
        RECT 2015.910 715.720 2018.750 718.070 ;
        RECT 2019.590 715.720 2022.430 718.070 ;
        RECT 2023.270 715.720 2026.110 718.070 ;
        RECT 2026.950 715.720 2029.790 718.070 ;
        RECT 2030.630 715.720 2033.470 718.070 ;
        RECT 2034.310 715.720 2037.150 718.070 ;
        RECT 2037.990 715.720 2040.830 718.070 ;
        RECT 2041.670 715.720 2044.510 718.070 ;
        RECT 2045.350 715.720 2048.190 718.070 ;
        RECT 2049.030 715.720 2051.870 718.070 ;
        RECT 2052.710 715.720 2055.550 718.070 ;
        RECT 2056.390 715.720 2059.230 718.070 ;
        RECT 2060.070 715.720 2062.910 718.070 ;
        RECT 2063.750 715.720 2066.590 718.070 ;
        RECT 2067.430 715.720 2070.270 718.070 ;
        RECT 2071.110 715.720 2073.950 718.070 ;
        RECT 2074.790 715.720 2077.630 718.070 ;
        RECT 2078.470 715.720 2081.310 718.070 ;
        RECT 2082.150 715.720 2084.990 718.070 ;
        RECT 2085.830 715.720 2088.670 718.070 ;
        RECT 2089.510 715.720 2092.350 718.070 ;
        RECT 2093.190 715.720 2096.030 718.070 ;
        RECT 2096.870 715.720 2099.710 718.070 ;
        RECT 2100.550 715.720 2103.390 718.070 ;
        RECT 2104.230 715.720 2107.070 718.070 ;
        RECT 2107.910 715.720 2110.750 718.070 ;
        RECT 2111.590 715.720 2114.430 718.070 ;
        RECT 2115.270 715.720 2118.110 718.070 ;
        RECT 2118.950 715.720 2121.790 718.070 ;
        RECT 2122.630 715.720 2125.470 718.070 ;
        RECT 2126.310 715.720 2129.150 718.070 ;
        RECT 2129.990 715.720 2132.830 718.070 ;
        RECT 2133.670 715.720 2136.510 718.070 ;
        RECT 2137.350 715.720 2140.190 718.070 ;
        RECT 2141.030 715.720 2143.870 718.070 ;
        RECT 2144.710 715.720 2147.550 718.070 ;
        RECT 2148.390 715.720 2151.230 718.070 ;
        RECT 2152.070 715.720 2154.910 718.070 ;
        RECT 2155.750 715.720 2158.590 718.070 ;
        RECT 2159.430 715.720 2162.270 718.070 ;
        RECT 2163.110 715.720 2165.950 718.070 ;
        RECT 2166.790 715.720 2169.630 718.070 ;
        RECT 2170.470 715.720 2173.310 718.070 ;
        RECT 2174.150 715.720 2176.990 718.070 ;
        RECT 2177.830 715.720 2180.670 718.070 ;
        RECT 2181.510 715.720 2184.350 718.070 ;
        RECT 2185.190 715.720 2188.030 718.070 ;
        RECT 2188.870 715.720 2191.710 718.070 ;
        RECT 2192.550 715.720 2195.390 718.070 ;
        RECT 2196.230 715.720 2199.070 718.070 ;
        RECT 2199.910 715.720 2202.750 718.070 ;
        RECT 2203.590 715.720 2206.430 718.070 ;
        RECT 2207.270 715.720 2210.110 718.070 ;
        RECT 2210.950 715.720 2213.790 718.070 ;
        RECT 2214.630 715.720 2217.470 718.070 ;
        RECT 2218.310 715.720 2221.150 718.070 ;
        RECT 2221.990 715.720 2224.830 718.070 ;
        RECT 2225.670 715.720 2228.510 718.070 ;
        RECT 2229.350 715.720 2232.190 718.070 ;
        RECT 2233.030 715.720 2235.870 718.070 ;
        RECT 2236.710 715.720 2239.550 718.070 ;
        RECT 2240.390 715.720 2243.230 718.070 ;
        RECT 2244.070 715.720 2246.910 718.070 ;
        RECT 2247.750 715.720 2250.590 718.070 ;
        RECT 2251.430 715.720 2254.270 718.070 ;
        RECT 2255.110 715.720 2257.950 718.070 ;
        RECT 2258.790 715.720 2261.630 718.070 ;
        RECT 2262.470 715.720 2265.310 718.070 ;
        RECT 2266.150 715.720 2268.990 718.070 ;
        RECT 2269.830 715.720 2272.670 718.070 ;
        RECT 2273.510 715.720 2276.350 718.070 ;
        RECT 2277.190 715.720 2280.030 718.070 ;
        RECT 2280.870 715.720 2283.710 718.070 ;
        RECT 2284.550 715.720 2287.390 718.070 ;
        RECT 2288.230 715.720 2291.070 718.070 ;
        RECT 2291.910 715.720 2294.750 718.070 ;
        RECT 2295.590 715.720 2298.430 718.070 ;
        RECT 2299.270 715.720 2302.110 718.070 ;
        RECT 2302.950 715.720 2305.790 718.070 ;
        RECT 2306.630 715.720 2309.470 718.070 ;
        RECT 2310.310 715.720 2313.150 718.070 ;
        RECT 2313.990 715.720 2316.830 718.070 ;
        RECT 2317.670 715.720 2320.510 718.070 ;
        RECT 2321.350 715.720 2324.190 718.070 ;
        RECT 2325.030 715.720 2327.870 718.070 ;
        RECT 2328.710 715.720 2331.550 718.070 ;
        RECT 2332.390 715.720 2335.230 718.070 ;
        RECT 2336.070 715.720 2338.910 718.070 ;
        RECT 2339.750 715.720 2342.590 718.070 ;
        RECT 2343.430 715.720 2346.270 718.070 ;
        RECT 2347.110 715.720 2349.950 718.070 ;
        RECT 2350.790 715.720 2353.630 718.070 ;
        RECT 2354.470 715.720 2357.310 718.070 ;
        RECT 2358.150 715.720 2360.990 718.070 ;
        RECT 2361.830 715.720 2364.670 718.070 ;
        RECT 2365.510 715.720 2368.350 718.070 ;
        RECT 2369.190 715.720 2372.030 718.070 ;
        RECT 2372.870 715.720 2375.710 718.070 ;
        RECT 2376.550 715.720 2379.390 718.070 ;
        RECT 2380.230 715.720 2383.070 718.070 ;
        RECT 2383.910 715.720 2386.750 718.070 ;
        RECT 2387.590 715.720 2390.430 718.070 ;
        RECT 2391.270 715.720 2394.110 718.070 ;
        RECT 2394.950 715.720 2499.550 718.070 ;
        RECT 13.900 4.280 2499.550 715.720 ;
        RECT 13.900 2.390 54.090 4.280 ;
        RECT 54.930 2.390 158.050 4.280 ;
        RECT 158.890 2.390 262.010 4.280 ;
        RECT 262.850 2.390 365.970 4.280 ;
        RECT 366.810 2.390 469.930 4.280 ;
        RECT 470.770 2.390 573.890 4.280 ;
        RECT 574.730 2.390 1717.450 4.280 ;
        RECT 1718.290 2.390 1821.410 4.280 ;
        RECT 1822.250 2.390 1925.370 4.280 ;
        RECT 1926.210 2.390 2029.330 4.280 ;
        RECT 2030.170 2.390 2133.290 4.280 ;
        RECT 2134.130 2.390 2237.250 4.280 ;
        RECT 2238.090 2.390 2341.210 4.280 ;
        RECT 2342.050 2.390 2445.170 4.280 ;
        RECT 2446.010 2.390 2499.550 4.280 ;
      LAYER met3 ;
        RECT 21.050 674.240 2499.575 711.105 ;
        RECT 21.050 672.840 2495.600 674.240 ;
        RECT 21.050 664.720 2499.575 672.840 ;
        RECT 21.050 663.320 2495.600 664.720 ;
        RECT 21.050 655.200 2499.575 663.320 ;
        RECT 21.050 653.800 2495.600 655.200 ;
        RECT 21.050 645.680 2499.575 653.800 ;
        RECT 21.050 644.280 2495.600 645.680 ;
        RECT 21.050 636.160 2499.575 644.280 ;
        RECT 21.050 634.760 2495.600 636.160 ;
        RECT 21.050 626.640 2499.575 634.760 ;
        RECT 21.050 625.240 2495.600 626.640 ;
        RECT 21.050 617.120 2499.575 625.240 ;
        RECT 21.050 615.720 2495.600 617.120 ;
        RECT 21.050 607.600 2499.575 615.720 ;
        RECT 21.050 606.200 2495.600 607.600 ;
        RECT 21.050 598.080 2499.575 606.200 ;
        RECT 21.050 596.680 2495.600 598.080 ;
        RECT 21.050 588.560 2499.575 596.680 ;
        RECT 21.050 587.160 2495.600 588.560 ;
        RECT 21.050 579.040 2499.575 587.160 ;
        RECT 21.050 577.640 2495.600 579.040 ;
        RECT 21.050 569.520 2499.575 577.640 ;
        RECT 21.050 568.120 2495.600 569.520 ;
        RECT 21.050 560.000 2499.575 568.120 ;
        RECT 21.050 558.600 2495.600 560.000 ;
        RECT 21.050 550.480 2499.575 558.600 ;
        RECT 21.050 549.080 2495.600 550.480 ;
        RECT 21.050 540.960 2499.575 549.080 ;
        RECT 21.050 539.560 2495.600 540.960 ;
        RECT 21.050 531.440 2499.575 539.560 ;
        RECT 21.050 530.040 2495.600 531.440 ;
        RECT 21.050 521.920 2499.575 530.040 ;
        RECT 21.050 520.520 2495.600 521.920 ;
        RECT 21.050 512.400 2499.575 520.520 ;
        RECT 21.050 511.000 2495.600 512.400 ;
        RECT 21.050 502.880 2499.575 511.000 ;
        RECT 21.050 501.480 2495.600 502.880 ;
        RECT 21.050 493.360 2499.575 501.480 ;
        RECT 21.050 491.960 2495.600 493.360 ;
        RECT 21.050 483.840 2499.575 491.960 ;
        RECT 21.050 482.440 2495.600 483.840 ;
        RECT 21.050 474.320 2499.575 482.440 ;
        RECT 21.050 472.920 2495.600 474.320 ;
        RECT 21.050 464.800 2499.575 472.920 ;
        RECT 21.050 463.400 2495.600 464.800 ;
        RECT 21.050 455.280 2499.575 463.400 ;
        RECT 21.050 453.880 2495.600 455.280 ;
        RECT 21.050 445.760 2499.575 453.880 ;
        RECT 21.050 444.360 2495.600 445.760 ;
        RECT 21.050 436.240 2499.575 444.360 ;
        RECT 21.050 434.840 2495.600 436.240 ;
        RECT 21.050 426.720 2499.575 434.840 ;
        RECT 21.050 425.320 2495.600 426.720 ;
        RECT 21.050 417.200 2499.575 425.320 ;
        RECT 21.050 415.800 2495.600 417.200 ;
        RECT 21.050 407.680 2499.575 415.800 ;
        RECT 21.050 406.280 2495.600 407.680 ;
        RECT 21.050 398.160 2499.575 406.280 ;
        RECT 21.050 396.760 2495.600 398.160 ;
        RECT 21.050 388.640 2499.575 396.760 ;
        RECT 21.050 387.240 2495.600 388.640 ;
        RECT 21.050 379.120 2499.575 387.240 ;
        RECT 21.050 377.720 2495.600 379.120 ;
        RECT 21.050 369.600 2499.575 377.720 ;
        RECT 21.050 368.200 2495.600 369.600 ;
        RECT 21.050 360.080 2499.575 368.200 ;
        RECT 21.050 358.680 2495.600 360.080 ;
        RECT 21.050 350.560 2499.575 358.680 ;
        RECT 21.050 349.160 2495.600 350.560 ;
        RECT 21.050 341.040 2499.575 349.160 ;
        RECT 21.050 339.640 2495.600 341.040 ;
        RECT 21.050 331.520 2499.575 339.640 ;
        RECT 21.050 330.120 2495.600 331.520 ;
        RECT 21.050 322.000 2499.575 330.120 ;
        RECT 21.050 320.600 2495.600 322.000 ;
        RECT 21.050 312.480 2499.575 320.600 ;
        RECT 21.050 311.080 2495.600 312.480 ;
        RECT 21.050 302.960 2499.575 311.080 ;
        RECT 21.050 301.560 2495.600 302.960 ;
        RECT 21.050 293.440 2499.575 301.560 ;
        RECT 21.050 292.040 2495.600 293.440 ;
        RECT 21.050 283.920 2499.575 292.040 ;
        RECT 21.050 282.520 2495.600 283.920 ;
        RECT 21.050 274.400 2499.575 282.520 ;
        RECT 21.050 273.000 2495.600 274.400 ;
        RECT 21.050 264.880 2499.575 273.000 ;
        RECT 21.050 263.480 2495.600 264.880 ;
        RECT 21.050 255.360 2499.575 263.480 ;
        RECT 21.050 253.960 2495.600 255.360 ;
        RECT 21.050 245.840 2499.575 253.960 ;
        RECT 21.050 244.440 2495.600 245.840 ;
        RECT 21.050 236.320 2499.575 244.440 ;
        RECT 21.050 234.920 2495.600 236.320 ;
        RECT 21.050 226.800 2499.575 234.920 ;
        RECT 21.050 225.400 2495.600 226.800 ;
        RECT 21.050 217.280 2499.575 225.400 ;
        RECT 21.050 215.880 2495.600 217.280 ;
        RECT 21.050 207.760 2499.575 215.880 ;
        RECT 21.050 206.360 2495.600 207.760 ;
        RECT 21.050 198.240 2499.575 206.360 ;
        RECT 21.050 196.840 2495.600 198.240 ;
        RECT 21.050 188.720 2499.575 196.840 ;
        RECT 21.050 187.320 2495.600 188.720 ;
        RECT 21.050 179.200 2499.575 187.320 ;
        RECT 21.050 177.800 2495.600 179.200 ;
        RECT 21.050 169.680 2499.575 177.800 ;
        RECT 21.050 168.280 2495.600 169.680 ;
        RECT 21.050 160.160 2499.575 168.280 ;
        RECT 21.050 158.760 2495.600 160.160 ;
        RECT 21.050 150.640 2499.575 158.760 ;
        RECT 21.050 149.240 2495.600 150.640 ;
        RECT 21.050 141.120 2499.575 149.240 ;
        RECT 21.050 139.720 2495.600 141.120 ;
        RECT 21.050 131.600 2499.575 139.720 ;
        RECT 21.050 130.200 2495.600 131.600 ;
        RECT 21.050 122.080 2499.575 130.200 ;
        RECT 21.050 120.680 2495.600 122.080 ;
        RECT 21.050 112.560 2499.575 120.680 ;
        RECT 21.050 111.160 2495.600 112.560 ;
        RECT 21.050 103.040 2499.575 111.160 ;
        RECT 21.050 101.640 2495.600 103.040 ;
        RECT 21.050 93.520 2499.575 101.640 ;
        RECT 21.050 92.120 2495.600 93.520 ;
        RECT 21.050 84.000 2499.575 92.120 ;
        RECT 21.050 82.600 2495.600 84.000 ;
        RECT 21.050 74.480 2499.575 82.600 ;
        RECT 21.050 73.080 2495.600 74.480 ;
        RECT 21.050 64.960 2499.575 73.080 ;
        RECT 21.050 63.560 2495.600 64.960 ;
        RECT 21.050 55.440 2499.575 63.560 ;
        RECT 21.050 54.040 2495.600 55.440 ;
        RECT 21.050 45.920 2499.575 54.040 ;
        RECT 21.050 44.520 2495.600 45.920 ;
        RECT 21.050 3.575 2499.575 44.520 ;
      LAYER met4 ;
        RECT 73.040 585.110 82.240 711.105 ;
        RECT 71.040 52.870 82.240 585.110 ;
        RECT 73.040 3.575 82.240 52.870 ;
        RECT 84.640 3.575 120.640 711.105 ;
        RECT 123.040 585.110 132.240 711.105 ;
        RECT 134.640 585.110 170.640 711.105 ;
        RECT 123.040 52.870 170.640 585.110 ;
        RECT 123.040 3.575 132.240 52.870 ;
        RECT 134.640 3.575 170.640 52.870 ;
        RECT 173.040 3.575 182.240 711.105 ;
        RECT 184.640 585.110 220.640 711.105 ;
        RECT 223.040 585.110 232.240 711.105 ;
        RECT 184.640 554.475 232.240 585.110 ;
        RECT 234.640 554.475 270.640 711.105 ;
        RECT 273.040 585.110 282.240 711.105 ;
        RECT 284.640 585.110 320.640 711.105 ;
        RECT 273.040 554.475 320.640 585.110 ;
        RECT 323.040 554.475 332.240 711.105 ;
        RECT 334.640 585.110 370.640 711.105 ;
        RECT 373.040 585.110 382.240 711.105 ;
        RECT 334.640 554.475 382.240 585.110 ;
        RECT 384.640 554.475 420.640 711.105 ;
        RECT 423.040 585.110 432.240 711.105 ;
        RECT 434.640 585.110 470.640 711.105 ;
        RECT 423.040 554.475 470.640 585.110 ;
        RECT 473.040 554.475 482.240 711.105 ;
        RECT 484.640 585.110 520.640 711.105 ;
        RECT 523.040 585.110 532.240 711.105 ;
        RECT 484.640 554.475 532.240 585.110 ;
        RECT 534.640 554.475 570.640 711.105 ;
        RECT 573.040 585.110 582.240 711.105 ;
        RECT 584.640 585.110 620.640 711.105 ;
        RECT 573.040 554.475 620.640 585.110 ;
        RECT 623.040 554.475 632.240 711.105 ;
        RECT 634.640 585.110 670.640 711.105 ;
        RECT 673.040 585.110 682.240 711.105 ;
        RECT 634.640 554.475 682.240 585.110 ;
        RECT 684.640 554.475 720.640 711.105 ;
        RECT 723.040 585.110 732.240 711.105 ;
        RECT 734.640 585.110 770.640 711.105 ;
        RECT 723.040 554.475 770.640 585.110 ;
        RECT 773.040 554.475 782.240 711.105 ;
        RECT 784.640 585.110 820.640 711.105 ;
        RECT 823.040 585.110 832.240 711.105 ;
        RECT 784.640 554.475 832.240 585.110 ;
        RECT 834.640 554.475 870.640 711.105 ;
        RECT 873.040 585.110 882.240 711.105 ;
        RECT 884.640 585.110 920.640 711.105 ;
        RECT 873.040 554.475 920.640 585.110 ;
        RECT 923.040 554.475 932.240 711.105 ;
        RECT 934.640 585.110 970.640 711.105 ;
        RECT 973.040 585.110 982.240 711.105 ;
        RECT 934.640 554.475 982.240 585.110 ;
        RECT 984.640 554.475 1020.640 711.105 ;
        RECT 1023.040 585.110 1032.240 711.105 ;
        RECT 1034.640 585.110 1070.640 711.105 ;
        RECT 1023.040 554.475 1070.640 585.110 ;
        RECT 1073.040 554.475 1082.240 711.105 ;
        RECT 1084.640 585.110 1120.640 711.105 ;
        RECT 1123.040 585.110 1132.240 711.105 ;
        RECT 1084.640 554.475 1132.240 585.110 ;
        RECT 1134.640 554.475 1170.640 711.105 ;
        RECT 1173.040 585.110 1182.240 711.105 ;
        RECT 1184.640 585.110 1220.640 711.105 ;
        RECT 1173.040 554.475 1220.640 585.110 ;
        RECT 184.640 104.585 1220.640 554.475 ;
        RECT 184.640 52.870 232.240 104.585 ;
        RECT 184.640 3.575 220.640 52.870 ;
        RECT 223.040 3.575 232.240 52.870 ;
        RECT 234.640 3.575 270.640 104.585 ;
        RECT 273.040 52.870 320.640 104.585 ;
        RECT 273.040 3.575 282.240 52.870 ;
        RECT 284.640 3.575 320.640 52.870 ;
        RECT 323.040 3.575 332.240 104.585 ;
        RECT 334.640 52.870 382.240 104.585 ;
        RECT 334.640 3.575 370.640 52.870 ;
        RECT 373.040 3.575 382.240 52.870 ;
        RECT 384.640 3.575 420.640 104.585 ;
        RECT 423.040 52.870 470.640 104.585 ;
        RECT 423.040 3.575 432.240 52.870 ;
        RECT 434.640 3.575 470.640 52.870 ;
        RECT 473.040 3.575 482.240 104.585 ;
        RECT 484.640 52.870 532.240 104.585 ;
        RECT 484.640 3.575 520.640 52.870 ;
        RECT 523.040 3.575 532.240 52.870 ;
        RECT 534.640 3.575 570.640 104.585 ;
        RECT 573.040 52.870 620.640 104.585 ;
        RECT 573.040 3.575 582.240 52.870 ;
        RECT 584.640 3.575 620.640 52.870 ;
        RECT 623.040 3.575 632.240 104.585 ;
        RECT 634.640 52.870 682.240 104.585 ;
        RECT 634.640 3.575 670.640 52.870 ;
        RECT 673.040 3.575 682.240 52.870 ;
        RECT 684.640 3.575 720.640 104.585 ;
        RECT 723.040 52.870 770.640 104.585 ;
        RECT 723.040 3.575 732.240 52.870 ;
        RECT 734.640 3.575 770.640 52.870 ;
        RECT 773.040 3.575 782.240 104.585 ;
        RECT 784.640 52.870 832.240 104.585 ;
        RECT 784.640 3.575 820.640 52.870 ;
        RECT 823.040 3.575 832.240 52.870 ;
        RECT 834.640 3.575 870.640 104.585 ;
        RECT 873.040 52.870 920.640 104.585 ;
        RECT 873.040 3.575 882.240 52.870 ;
        RECT 884.640 3.575 920.640 52.870 ;
        RECT 923.040 3.575 932.240 104.585 ;
        RECT 934.640 52.870 982.240 104.585 ;
        RECT 934.640 3.575 970.640 52.870 ;
        RECT 973.040 3.575 982.240 52.870 ;
        RECT 984.640 3.575 1020.640 104.585 ;
        RECT 1023.040 52.870 1070.640 104.585 ;
        RECT 1023.040 3.575 1032.240 52.870 ;
        RECT 1034.640 3.575 1070.640 52.870 ;
        RECT 1073.040 3.575 1082.240 104.585 ;
        RECT 1084.640 52.870 1132.240 104.585 ;
        RECT 1084.640 3.575 1120.640 52.870 ;
        RECT 1123.040 3.575 1132.240 52.870 ;
        RECT 1134.640 3.575 1170.640 104.585 ;
        RECT 1173.040 52.870 1220.640 104.585 ;
        RECT 1173.040 3.575 1182.240 52.870 ;
        RECT 1184.640 3.575 1220.640 52.870 ;
        RECT 1223.040 3.575 1232.240 711.105 ;
        RECT 1234.640 3.575 1270.640 711.105 ;
        RECT 1273.040 3.575 1282.240 711.105 ;
        RECT 1284.640 3.575 1320.640 711.105 ;
        RECT 1323.040 3.575 1332.240 711.105 ;
        RECT 1334.640 3.575 1370.640 711.105 ;
        RECT 1373.040 3.575 1382.240 711.105 ;
        RECT 1384.640 3.575 1420.640 711.105 ;
        RECT 1423.040 3.575 1432.240 711.105 ;
        RECT 1434.640 3.575 1470.640 711.105 ;
        RECT 1473.040 3.575 1482.240 711.105 ;
        RECT 1484.640 3.575 1520.640 711.105 ;
        RECT 1523.040 3.575 1532.240 711.105 ;
        RECT 1534.640 3.575 1570.640 711.105 ;
        RECT 1573.040 3.575 1582.240 711.105 ;
        RECT 1584.640 3.575 1620.640 711.105 ;
        RECT 1623.040 3.575 1632.240 711.105 ;
        RECT 1634.640 3.575 1670.640 711.105 ;
        RECT 1673.040 3.575 1682.240 711.105 ;
        RECT 1684.640 3.575 1720.640 711.105 ;
        RECT 1723.040 3.575 1732.240 711.105 ;
        RECT 1734.640 3.575 1770.640 711.105 ;
        RECT 1773.040 3.575 1782.240 711.105 ;
        RECT 1784.640 3.575 1820.640 711.105 ;
        RECT 1823.040 3.575 1832.240 711.105 ;
        RECT 1834.640 3.575 1870.640 711.105 ;
        RECT 1873.040 3.575 1882.240 711.105 ;
        RECT 1884.640 3.575 1920.640 711.105 ;
        RECT 1923.040 3.575 1932.240 711.105 ;
        RECT 1934.640 3.575 1970.640 711.105 ;
        RECT 1973.040 3.575 1982.240 711.105 ;
        RECT 1984.640 580.760 2020.640 711.105 ;
        RECT 2023.040 580.760 2032.240 711.105 ;
        RECT 2034.640 580.760 2070.640 711.105 ;
        RECT 2073.040 580.760 2082.240 711.105 ;
        RECT 2084.640 580.760 2120.640 711.105 ;
        RECT 2123.040 580.760 2132.240 711.105 ;
        RECT 2134.640 580.760 2170.640 711.105 ;
        RECT 2173.040 580.760 2182.240 711.105 ;
        RECT 2184.640 580.760 2220.640 711.105 ;
        RECT 2223.040 580.760 2232.240 711.105 ;
        RECT 2234.640 580.760 2270.640 711.105 ;
        RECT 2273.040 580.760 2282.240 711.105 ;
        RECT 2284.640 580.760 2320.640 711.105 ;
        RECT 2323.040 580.760 2332.240 711.105 ;
        RECT 2334.640 580.760 2370.640 711.105 ;
        RECT 2373.040 580.760 2382.240 711.105 ;
        RECT 2384.640 580.760 2420.640 711.105 ;
        RECT 2423.040 580.760 2432.240 711.105 ;
        RECT 2434.640 580.760 2470.640 711.105 ;
        RECT 1984.640 70.350 2470.640 580.760 ;
        RECT 1984.640 3.575 2020.640 70.350 ;
        RECT 2023.040 3.575 2032.240 70.350 ;
        RECT 2034.640 3.575 2070.640 70.350 ;
        RECT 2073.040 3.575 2082.240 70.350 ;
        RECT 2084.640 3.575 2120.640 70.350 ;
        RECT 2123.040 3.575 2132.240 70.350 ;
        RECT 2134.640 3.575 2170.640 70.350 ;
        RECT 2173.040 3.575 2182.240 70.350 ;
        RECT 2184.640 3.575 2220.640 70.350 ;
        RECT 2223.040 3.575 2232.240 70.350 ;
        RECT 2234.640 3.575 2270.640 70.350 ;
        RECT 2273.040 3.575 2282.240 70.350 ;
        RECT 2284.640 3.575 2320.640 70.350 ;
        RECT 2323.040 3.575 2332.240 70.350 ;
        RECT 2334.640 3.575 2370.640 70.350 ;
        RECT 2373.040 3.575 2382.240 70.350 ;
        RECT 2384.640 3.575 2420.640 70.350 ;
        RECT 2423.040 3.575 2432.240 70.350 ;
        RECT 2434.640 3.575 2470.640 70.350 ;
        RECT 2473.040 3.575 2482.240 711.105 ;
        RECT 2484.640 3.575 2496.090 711.105 ;
      LAYER met5 ;
        RECT 697.940 691.530 2496.300 706.300 ;
        RECT 697.940 679.930 2496.300 686.730 ;
        RECT 697.940 641.530 2496.300 675.130 ;
        RECT 697.940 629.930 2496.300 636.730 ;
        RECT 697.940 591.530 2496.300 625.130 ;
        RECT 697.940 579.930 2496.300 586.730 ;
        RECT 697.940 541.530 2496.300 575.130 ;
        RECT 697.940 529.930 2496.300 536.730 ;
        RECT 697.940 491.530 2496.300 525.130 ;
        RECT 697.940 479.930 2496.300 486.730 ;
        RECT 697.940 441.530 2496.300 475.130 ;
        RECT 697.940 429.930 2496.300 436.730 ;
        RECT 697.940 391.530 2496.300 425.130 ;
        RECT 697.940 379.930 2496.300 386.730 ;
        RECT 697.940 341.530 2496.300 375.130 ;
        RECT 697.940 329.930 2496.300 336.730 ;
        RECT 697.940 291.530 2496.300 325.130 ;
        RECT 697.940 279.930 2496.300 286.730 ;
        RECT 697.940 241.530 2496.300 275.130 ;
        RECT 697.940 229.930 2496.300 236.730 ;
        RECT 697.940 191.530 2496.300 225.130 ;
        RECT 697.940 179.930 2496.300 186.730 ;
        RECT 697.940 141.530 2496.300 175.130 ;
        RECT 697.940 129.930 2496.300 136.730 ;
        RECT 697.940 91.530 2496.300 125.130 ;
        RECT 697.940 79.930 2496.300 86.730 ;
        RECT 697.940 41.530 2496.300 75.130 ;
        RECT 697.940 29.930 2496.300 36.730 ;
        RECT 697.940 11.100 2496.300 25.130 ;
  END
END mgmt_core_wrapper
END LIBRARY

