VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_core
  CLASS BLOCK ;
  FOREIGN mgmt_core ;
  ORIGIN 0.000 0.000 ;
  SIZE 2000.000 BY 740.000 ;
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 0.020 0.780 1999.600 2.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 91.490 1999.600 93.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 221.490 1999.600 223.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 351.490 1999.600 353.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 481.490 1999.600 483.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 611.490 1999.600 613.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 737.460 1999.600 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 100.640 0.780 102.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 150.640 0.780 152.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 200.640 0.780 202.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 250.640 0.780 252.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 300.640 0.780 302.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 350.640 0.780 352.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 400.640 0.780 402.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 450.640 0.780 452.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 500.640 0.780 502.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 550.640 0.780 552.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 600.640 0.780 602.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 650.640 0.780 652.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 700.640 0.780 702.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 750.640 0.780 752.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 0.020 0.780 1.620 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 50.640 0.780 52.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 100.640 537.300 102.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 150.640 537.300 152.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 200.640 537.300 202.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 250.640 537.300 252.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 300.640 537.300 302.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 350.640 537.300 352.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 400.640 537.300 402.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 450.640 537.300 452.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 500.640 537.300 502.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 550.640 537.300 552.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 600.640 537.300 602.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 650.640 537.300 652.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 700.640 537.300 702.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 750.640 537.300 752.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 800.640 0.780 802.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 850.640 0.780 852.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 900.640 0.780 902.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 950.640 0.780 952.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1000.640 0.780 1002.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1050.640 0.780 1052.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1100.640 0.780 1102.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1150.640 0.780 1152.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1200.640 0.780 1202.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1250.640 0.780 1252.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1300.640 0.780 1302.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1350.640 0.780 1352.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1400.640 0.780 1402.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1450.640 0.780 1452.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1500.640 0.780 1502.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1550.640 0.780 1552.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1600.640 0.780 1602.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1650.640 0.780 1652.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1700.640 0.780 1702.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1750.640 0.780 1752.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1800.640 0.780 1802.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1850.640 0.780 1852.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1900.640 0.780 1902.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1950.640 0.780 1952.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1998.000 0.780 1999.600 739.060 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 3.320 4.080 1996.300 5.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 26.490 1999.600 28.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 156.490 1999.600 158.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 286.490 1999.600 288.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 416.490 1999.600 418.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 546.490 1999.600 548.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 0.020 676.490 1999.600 678.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 3.320 734.160 1996.300 735.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.640 0.780 127.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 175.640 0.780 177.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 225.640 0.780 227.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 275.640 0.780 277.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.640 0.780 327.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 375.640 0.780 377.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 425.640 0.780 427.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 475.640 0.780 477.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 525.640 0.780 527.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.640 0.780 577.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 625.640 0.780 627.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.640 0.780 677.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 725.640 0.780 727.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 775.640 0.780 777.240 101.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 3.320 4.080 4.920 735.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 1994.700 4.080 1996.300 735.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 25.640 0.780 27.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 75.640 0.780 77.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 125.640 537.300 127.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 175.640 537.300 177.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 225.640 537.300 227.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 275.640 537.300 277.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 325.640 537.300 327.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 375.640 537.300 377.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 425.640 537.300 427.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 475.640 537.300 477.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 525.640 537.300 527.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 575.640 537.300 577.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 625.640 537.300 627.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 675.640 537.300 677.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 725.640 537.300 727.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 775.640 537.300 777.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 825.640 0.780 827.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 875.640 0.780 877.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 925.640 0.780 927.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 975.640 0.780 977.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1025.640 0.780 1027.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1075.640 0.780 1077.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1125.640 0.780 1127.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1175.640 0.780 1177.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1225.640 0.780 1227.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1275.640 0.780 1277.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1325.640 0.780 1327.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1375.640 0.780 1377.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1425.640 0.780 1427.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.640 0.780 1477.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1525.640 0.780 1527.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1575.640 0.780 1577.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1625.640 0.780 1627.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1675.640 0.780 1677.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1725.640 0.780 1727.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1775.640 0.780 1777.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1825.640 0.780 1827.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1875.640 0.780 1877.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1925.640 0.780 1927.240 739.060 ;
    END
    PORT
      LAYER met4 ;
        RECT 1975.640 0.780 1977.240 739.060 ;
    END
  END VPWR
  PIN core_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 736.000 1.750 740.000 ;
    END
  END core_clk
  PIN core_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.690 736.000 4.970 740.000 ;
    END
  END core_rstn
  PIN debug_mode
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.010 0.000 1588.290 4.000 ;
    END
  END debug_mode
  PIN debug_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1605.030 0.000 1605.310 4.000 ;
    END
  END debug_oeb
  PIN debug_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1916.910 736.000 1917.190 740.000 ;
    END
  END debug_rx
  PIN debug_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.800 4.000 430.400 ;
    END
  END debug_tx
  PIN flash_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 4.000 ;
    END
  END flash_clk
  PIN flash_cs_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1688.750 0.000 1689.030 4.000 ;
    END
  END flash_cs_n
  PIN flash_io0_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END flash_io0_di
  PIN flash_io0_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END flash_io0_do
  PIN flash_io0_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END flash_io0_oeb
  PIN flash_io1_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.270 0.000 176.550 4.000 ;
    END
  END flash_io1_di
  PIN flash_io1_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.830 0.000 193.110 4.000 ;
    END
  END flash_io1_do
  PIN flash_io1_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END flash_io1_oeb
  PIN flash_io2_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END flash_io2_di
  PIN flash_io2_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 0.000 243.710 4.000 ;
    END
  END flash_io2_do
  PIN flash_io2_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END flash_io2_oeb
  PIN flash_io3_di
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END flash_io3_di
  PIN flash_io3_do
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.010 0.000 277.290 4.000 ;
    END
  END flash_io3_do
  PIN flash_io3_oeb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END flash_io3_oeb
  PIN gpio_in_pad
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.370 0.000 8.650 4.000 ;
    END
  END gpio_in_pad
  PIN gpio_inenb_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 4.000 ;
    END
  END gpio_inenb_pad
  PIN gpio_mode0_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END gpio_mode0_pad
  PIN gpio_mode1_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.510 0.000 58.790 4.000 ;
    END
  END gpio_mode1_pad
  PIN gpio_out_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END gpio_out_pad
  PIN gpio_outenb_pad
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END gpio_outenb_pad
  PIN hk_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.590 0.000 310.870 4.000 ;
    END
  END hk_ack_i
  PIN hk_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1920.130 736.000 1920.410 740.000 ;
    END
  END hk_cyc_o
  PIN hk_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END hk_dat_i[0]
  PIN hk_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.530 0.000 512.810 4.000 ;
    END
  END hk_dat_i[10]
  PIN hk_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.090 0.000 529.370 4.000 ;
    END
  END hk_dat_i[11]
  PIN hk_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 0.000 546.390 4.000 ;
    END
  END hk_dat_i[12]
  PIN hk_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.670 0.000 562.950 4.000 ;
    END
  END hk_dat_i[13]
  PIN hk_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END hk_dat_i[14]
  PIN hk_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 0.000 596.530 4.000 ;
    END
  END hk_dat_i[15]
  PIN hk_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.270 0.000 613.550 4.000 ;
    END
  END hk_dat_i[16]
  PIN hk_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.830 0.000 630.110 4.000 ;
    END
  END hk_dat_i[17]
  PIN hk_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.850 0.000 647.130 4.000 ;
    END
  END hk_dat_i[18]
  PIN hk_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END hk_dat_i[19]
  PIN hk_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 0.000 361.470 4.000 ;
    END
  END hk_dat_i[1]
  PIN hk_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.430 0.000 680.710 4.000 ;
    END
  END hk_dat_i[20]
  PIN hk_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 0.000 697.730 4.000 ;
    END
  END hk_dat_i[21]
  PIN hk_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.010 0.000 714.290 4.000 ;
    END
  END hk_dat_i[22]
  PIN hk_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 731.030 0.000 731.310 4.000 ;
    END
  END hk_dat_i[23]
  PIN hk_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.590 0.000 747.870 4.000 ;
    END
  END hk_dat_i[24]
  PIN hk_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.610 0.000 764.890 4.000 ;
    END
  END hk_dat_i[25]
  PIN hk_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.170 0.000 781.450 4.000 ;
    END
  END hk_dat_i[26]
  PIN hk_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 0.000 798.470 4.000 ;
    END
  END hk_dat_i[27]
  PIN hk_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.750 0.000 815.030 4.000 ;
    END
  END hk_dat_i[28]
  PIN hk_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 831.770 0.000 832.050 4.000 ;
    END
  END hk_dat_i[29]
  PIN hk_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END hk_dat_i[2]
  PIN hk_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 848.330 0.000 848.610 4.000 ;
    END
  END hk_dat_i[30]
  PIN hk_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.350 0.000 865.630 4.000 ;
    END
  END hk_dat_i[31]
  PIN hk_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END hk_dat_i[3]
  PIN hk_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 4.000 ;
    END
  END hk_dat_i[4]
  PIN hk_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END hk_dat_i[5]
  PIN hk_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.910 0.000 445.190 4.000 ;
    END
  END hk_dat_i[6]
  PIN hk_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.930 0.000 462.210 4.000 ;
    END
  END hk_dat_i[7]
  PIN hk_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END hk_dat_i[8]
  PIN hk_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 0.000 495.790 4.000 ;
    END
  END hk_dat_i[9]
  PIN hk_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 4.000 ;
    END
  END hk_stb_o
  PIN la_iena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.910 736.000 8.190 740.000 ;
    END
  END la_iena[0]
  PIN la_iena[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.790 736.000 1309.070 740.000 ;
    END
  END la_iena[100]
  PIN la_iena[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1321.670 736.000 1321.950 740.000 ;
    END
  END la_iena[101]
  PIN la_iena[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1334.550 736.000 1334.830 740.000 ;
    END
  END la_iena[102]
  PIN la_iena[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1347.430 736.000 1347.710 740.000 ;
    END
  END la_iena[103]
  PIN la_iena[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1360.770 736.000 1361.050 740.000 ;
    END
  END la_iena[104]
  PIN la_iena[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.650 736.000 1373.930 740.000 ;
    END
  END la_iena[105]
  PIN la_iena[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.530 736.000 1386.810 740.000 ;
    END
  END la_iena[106]
  PIN la_iena[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.870 736.000 1400.150 740.000 ;
    END
  END la_iena[107]
  PIN la_iena[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1412.750 736.000 1413.030 740.000 ;
    END
  END la_iena[108]
  PIN la_iena[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1425.630 736.000 1425.910 740.000 ;
    END
  END la_iena[109]
  PIN la_iena[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.630 736.000 137.910 740.000 ;
    END
  END la_iena[10]
  PIN la_iena[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.510 736.000 1438.790 740.000 ;
    END
  END la_iena[110]
  PIN la_iena[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1451.850 736.000 1452.130 740.000 ;
    END
  END la_iena[111]
  PIN la_iena[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1464.730 736.000 1465.010 740.000 ;
    END
  END la_iena[112]
  PIN la_iena[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1477.610 736.000 1477.890 740.000 ;
    END
  END la_iena[113]
  PIN la_iena[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1490.950 736.000 1491.230 740.000 ;
    END
  END la_iena[114]
  PIN la_iena[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.830 736.000 1504.110 740.000 ;
    END
  END la_iena[115]
  PIN la_iena[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1516.710 736.000 1516.990 740.000 ;
    END
  END la_iena[116]
  PIN la_iena[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1529.590 736.000 1529.870 740.000 ;
    END
  END la_iena[117]
  PIN la_iena[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1542.930 736.000 1543.210 740.000 ;
    END
  END la_iena[118]
  PIN la_iena[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.810 736.000 1556.090 740.000 ;
    END
  END la_iena[119]
  PIN la_iena[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 736.000 151.250 740.000 ;
    END
  END la_iena[11]
  PIN la_iena[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1568.690 736.000 1568.970 740.000 ;
    END
  END la_iena[120]
  PIN la_iena[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.570 736.000 1581.850 740.000 ;
    END
  END la_iena[121]
  PIN la_iena[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1594.910 736.000 1595.190 740.000 ;
    END
  END la_iena[122]
  PIN la_iena[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1607.790 736.000 1608.070 740.000 ;
    END
  END la_iena[123]
  PIN la_iena[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1620.670 736.000 1620.950 740.000 ;
    END
  END la_iena[124]
  PIN la_iena[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1634.010 736.000 1634.290 740.000 ;
    END
  END la_iena[125]
  PIN la_iena[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1646.890 736.000 1647.170 740.000 ;
    END
  END la_iena[126]
  PIN la_iena[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1659.770 736.000 1660.050 740.000 ;
    END
  END la_iena[127]
  PIN la_iena[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 736.000 164.130 740.000 ;
    END
  END la_iena[12]
  PIN la_iena[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.730 736.000 177.010 740.000 ;
    END
  END la_iena[13]
  PIN la_iena[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 736.000 190.350 740.000 ;
    END
  END la_iena[14]
  PIN la_iena[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 736.000 203.230 740.000 ;
    END
  END la_iena[15]
  PIN la_iena[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 736.000 216.110 740.000 ;
    END
  END la_iena[16]
  PIN la_iena[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 736.000 228.990 740.000 ;
    END
  END la_iena[17]
  PIN la_iena[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 736.000 242.330 740.000 ;
    END
  END la_iena[18]
  PIN la_iena[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 736.000 255.210 740.000 ;
    END
  END la_iena[19]
  PIN la_iena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 736.000 21.070 740.000 ;
    END
  END la_iena[1]
  PIN la_iena[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 736.000 268.090 740.000 ;
    END
  END la_iena[20]
  PIN la_iena[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 736.000 281.430 740.000 ;
    END
  END la_iena[21]
  PIN la_iena[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 736.000 294.310 740.000 ;
    END
  END la_iena[22]
  PIN la_iena[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 736.000 307.190 740.000 ;
    END
  END la_iena[23]
  PIN la_iena[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.790 736.000 320.070 740.000 ;
    END
  END la_iena[24]
  PIN la_iena[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 736.000 333.410 740.000 ;
    END
  END la_iena[25]
  PIN la_iena[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.010 736.000 346.290 740.000 ;
    END
  END la_iena[26]
  PIN la_iena[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 736.000 359.170 740.000 ;
    END
  END la_iena[27]
  PIN la_iena[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.770 736.000 372.050 740.000 ;
    END
  END la_iena[28]
  PIN la_iena[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 736.000 385.390 740.000 ;
    END
  END la_iena[29]
  PIN la_iena[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 736.000 33.950 740.000 ;
    END
  END la_iena[2]
  PIN la_iena[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.990 736.000 398.270 740.000 ;
    END
  END la_iena[30]
  PIN la_iena[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.870 736.000 411.150 740.000 ;
    END
  END la_iena[31]
  PIN la_iena[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.210 736.000 424.490 740.000 ;
    END
  END la_iena[32]
  PIN la_iena[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 736.000 437.370 740.000 ;
    END
  END la_iena[33]
  PIN la_iena[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.970 736.000 450.250 740.000 ;
    END
  END la_iena[34]
  PIN la_iena[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.850 736.000 463.130 740.000 ;
    END
  END la_iena[35]
  PIN la_iena[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.190 736.000 476.470 740.000 ;
    END
  END la_iena[36]
  PIN la_iena[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.070 736.000 489.350 740.000 ;
    END
  END la_iena[37]
  PIN la_iena[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.950 736.000 502.230 740.000 ;
    END
  END la_iena[38]
  PIN la_iena[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 736.000 515.570 740.000 ;
    END
  END la_iena[39]
  PIN la_iena[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 736.000 46.830 740.000 ;
    END
  END la_iena[3]
  PIN la_iena[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 736.000 528.450 740.000 ;
    END
  END la_iena[40]
  PIN la_iena[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 736.000 541.330 740.000 ;
    END
  END la_iena[41]
  PIN la_iena[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 736.000 554.210 740.000 ;
    END
  END la_iena[42]
  PIN la_iena[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.270 736.000 567.550 740.000 ;
    END
  END la_iena[43]
  PIN la_iena[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 580.150 736.000 580.430 740.000 ;
    END
  END la_iena[44]
  PIN la_iena[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.030 736.000 593.310 740.000 ;
    END
  END la_iena[45]
  PIN la_iena[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 736.000 606.650 740.000 ;
    END
  END la_iena[46]
  PIN la_iena[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.250 736.000 619.530 740.000 ;
    END
  END la_iena[47]
  PIN la_iena[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.130 736.000 632.410 740.000 ;
    END
  END la_iena[48]
  PIN la_iena[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.010 736.000 645.290 740.000 ;
    END
  END la_iena[49]
  PIN la_iena[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 736.000 60.170 740.000 ;
    END
  END la_iena[4]
  PIN la_iena[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.350 736.000 658.630 740.000 ;
    END
  END la_iena[50]
  PIN la_iena[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.230 736.000 671.510 740.000 ;
    END
  END la_iena[51]
  PIN la_iena[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 684.110 736.000 684.390 740.000 ;
    END
  END la_iena[52]
  PIN la_iena[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.990 736.000 697.270 740.000 ;
    END
  END la_iena[53]
  PIN la_iena[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 736.000 710.610 740.000 ;
    END
  END la_iena[54]
  PIN la_iena[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.210 736.000 723.490 740.000 ;
    END
  END la_iena[55]
  PIN la_iena[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 736.090 736.000 736.370 740.000 ;
    END
  END la_iena[56]
  PIN la_iena[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 736.000 749.710 740.000 ;
    END
  END la_iena[57]
  PIN la_iena[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.310 736.000 762.590 740.000 ;
    END
  END la_iena[58]
  PIN la_iena[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 775.190 736.000 775.470 740.000 ;
    END
  END la_iena[59]
  PIN la_iena[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.770 736.000 73.050 740.000 ;
    END
  END la_iena[5]
  PIN la_iena[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.070 736.000 788.350 740.000 ;
    END
  END la_iena[60]
  PIN la_iena[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.410 736.000 801.690 740.000 ;
    END
  END la_iena[61]
  PIN la_iena[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 814.290 736.000 814.570 740.000 ;
    END
  END la_iena[62]
  PIN la_iena[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.170 736.000 827.450 740.000 ;
    END
  END la_iena[63]
  PIN la_iena[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.510 736.000 840.790 740.000 ;
    END
  END la_iena[64]
  PIN la_iena[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 736.000 853.670 740.000 ;
    END
  END la_iena[65]
  PIN la_iena[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.270 736.000 866.550 740.000 ;
    END
  END la_iena[66]
  PIN la_iena[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 736.000 879.430 740.000 ;
    END
  END la_iena[67]
  PIN la_iena[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 892.490 736.000 892.770 740.000 ;
    END
  END la_iena[68]
  PIN la_iena[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.370 736.000 905.650 740.000 ;
    END
  END la_iena[69]
  PIN la_iena[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 736.000 85.930 740.000 ;
    END
  END la_iena[6]
  PIN la_iena[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.250 736.000 918.530 740.000 ;
    END
  END la_iena[70]
  PIN la_iena[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.130 736.000 931.410 740.000 ;
    END
  END la_iena[71]
  PIN la_iena[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.470 736.000 944.750 740.000 ;
    END
  END la_iena[72]
  PIN la_iena[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 957.350 736.000 957.630 740.000 ;
    END
  END la_iena[73]
  PIN la_iena[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.230 736.000 970.510 740.000 ;
    END
  END la_iena[74]
  PIN la_iena[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.570 736.000 983.850 740.000 ;
    END
  END la_iena[75]
  PIN la_iena[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 996.450 736.000 996.730 740.000 ;
    END
  END la_iena[76]
  PIN la_iena[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.330 736.000 1009.610 740.000 ;
    END
  END la_iena[77]
  PIN la_iena[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.210 736.000 1022.490 740.000 ;
    END
  END la_iena[78]
  PIN la_iena[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1035.550 736.000 1035.830 740.000 ;
    END
  END la_iena[79]
  PIN la_iena[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.990 736.000 99.270 740.000 ;
    END
  END la_iena[7]
  PIN la_iena[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.430 736.000 1048.710 740.000 ;
    END
  END la_iena[80]
  PIN la_iena[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.310 736.000 1061.590 740.000 ;
    END
  END la_iena[81]
  PIN la_iena[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1074.650 736.000 1074.930 740.000 ;
    END
  END la_iena[82]
  PIN la_iena[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1087.530 736.000 1087.810 740.000 ;
    END
  END la_iena[83]
  PIN la_iena[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1100.410 736.000 1100.690 740.000 ;
    END
  END la_iena[84]
  PIN la_iena[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.290 736.000 1113.570 740.000 ;
    END
  END la_iena[85]
  PIN la_iena[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1126.630 736.000 1126.910 740.000 ;
    END
  END la_iena[86]
  PIN la_iena[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1139.510 736.000 1139.790 740.000 ;
    END
  END la_iena[87]
  PIN la_iena[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.390 736.000 1152.670 740.000 ;
    END
  END la_iena[88]
  PIN la_iena[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1165.730 736.000 1166.010 740.000 ;
    END
  END la_iena[89]
  PIN la_iena[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870 736.000 112.150 740.000 ;
    END
  END la_iena[8]
  PIN la_iena[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.610 736.000 1178.890 740.000 ;
    END
  END la_iena[90]
  PIN la_iena[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.490 736.000 1191.770 740.000 ;
    END
  END la_iena[91]
  PIN la_iena[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1204.370 736.000 1204.650 740.000 ;
    END
  END la_iena[92]
  PIN la_iena[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1217.710 736.000 1217.990 740.000 ;
    END
  END la_iena[93]
  PIN la_iena[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.590 736.000 1230.870 740.000 ;
    END
  END la_iena[94]
  PIN la_iena[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.470 736.000 1243.750 740.000 ;
    END
  END la_iena[95]
  PIN la_iena[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1256.350 736.000 1256.630 740.000 ;
    END
  END la_iena[96]
  PIN la_iena[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.690 736.000 1269.970 740.000 ;
    END
  END la_iena[97]
  PIN la_iena[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1282.570 736.000 1282.850 740.000 ;
    END
  END la_iena[98]
  PIN la_iena[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1295.450 736.000 1295.730 740.000 ;
    END
  END la_iena[99]
  PIN la_iena[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 736.000 125.030 740.000 ;
    END
  END la_iena[9]
  PIN la_input[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.130 736.000 11.410 740.000 ;
    END
  END la_input[0]
  PIN la_input[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.010 736.000 1312.290 740.000 ;
    END
  END la_input[100]
  PIN la_input[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1324.890 736.000 1325.170 740.000 ;
    END
  END la_input[101]
  PIN la_input[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1337.770 736.000 1338.050 740.000 ;
    END
  END la_input[102]
  PIN la_input[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1351.110 736.000 1351.390 740.000 ;
    END
  END la_input[103]
  PIN la_input[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1363.990 736.000 1364.270 740.000 ;
    END
  END la_input[104]
  PIN la_input[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1376.870 736.000 1377.150 740.000 ;
    END
  END la_input[105]
  PIN la_input[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1389.750 736.000 1390.030 740.000 ;
    END
  END la_input[106]
  PIN la_input[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.090 736.000 1403.370 740.000 ;
    END
  END la_input[107]
  PIN la_input[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.970 736.000 1416.250 740.000 ;
    END
  END la_input[108]
  PIN la_input[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1428.850 736.000 1429.130 740.000 ;
    END
  END la_input[109]
  PIN la_input[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.310 736.000 141.590 740.000 ;
    END
  END la_input[10]
  PIN la_input[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1441.730 736.000 1442.010 740.000 ;
    END
  END la_input[110]
  PIN la_input[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1455.070 736.000 1455.350 740.000 ;
    END
  END la_input[111]
  PIN la_input[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.950 736.000 1468.230 740.000 ;
    END
  END la_input[112]
  PIN la_input[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.830 736.000 1481.110 740.000 ;
    END
  END la_input[113]
  PIN la_input[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.170 736.000 1494.450 740.000 ;
    END
  END la_input[114]
  PIN la_input[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1507.050 736.000 1507.330 740.000 ;
    END
  END la_input[115]
  PIN la_input[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.930 736.000 1520.210 740.000 ;
    END
  END la_input[116]
  PIN la_input[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1532.810 736.000 1533.090 740.000 ;
    END
  END la_input[117]
  PIN la_input[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1546.150 736.000 1546.430 740.000 ;
    END
  END la_input[118]
  PIN la_input[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1559.030 736.000 1559.310 740.000 ;
    END
  END la_input[119]
  PIN la_input[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.190 736.000 154.470 740.000 ;
    END
  END la_input[11]
  PIN la_input[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.910 736.000 1572.190 740.000 ;
    END
  END la_input[120]
  PIN la_input[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1585.250 736.000 1585.530 740.000 ;
    END
  END la_input[121]
  PIN la_input[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.130 736.000 1598.410 740.000 ;
    END
  END la_input[122]
  PIN la_input[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.010 736.000 1611.290 740.000 ;
    END
  END la_input[123]
  PIN la_input[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1623.890 736.000 1624.170 740.000 ;
    END
  END la_input[124]
  PIN la_input[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1637.230 736.000 1637.510 740.000 ;
    END
  END la_input[125]
  PIN la_input[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1650.110 736.000 1650.390 740.000 ;
    END
  END la_input[126]
  PIN la_input[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.990 736.000 1663.270 740.000 ;
    END
  END la_input[127]
  PIN la_input[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 736.000 167.350 740.000 ;
    END
  END la_input[12]
  PIN la_input[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 736.000 180.230 740.000 ;
    END
  END la_input[13]
  PIN la_input[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 736.000 193.570 740.000 ;
    END
  END la_input[14]
  PIN la_input[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 736.000 206.450 740.000 ;
    END
  END la_input[15]
  PIN la_input[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 736.000 219.330 740.000 ;
    END
  END la_input[16]
  PIN la_input[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 736.000 232.210 740.000 ;
    END
  END la_input[17]
  PIN la_input[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 245.270 736.000 245.550 740.000 ;
    END
  END la_input[18]
  PIN la_input[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 736.000 258.430 740.000 ;
    END
  END la_input[19]
  PIN la_input[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 736.000 24.290 740.000 ;
    END
  END la_input[1]
  PIN la_input[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.030 736.000 271.310 740.000 ;
    END
  END la_input[20]
  PIN la_input[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 736.000 284.650 740.000 ;
    END
  END la_input[21]
  PIN la_input[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 736.000 297.530 740.000 ;
    END
  END la_input[22]
  PIN la_input[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.130 736.000 310.410 740.000 ;
    END
  END la_input[23]
  PIN la_input[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.010 736.000 323.290 740.000 ;
    END
  END la_input[24]
  PIN la_input[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.350 736.000 336.630 740.000 ;
    END
  END la_input[25]
  PIN la_input[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.230 736.000 349.510 740.000 ;
    END
  END la_input[26]
  PIN la_input[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.110 736.000 362.390 740.000 ;
    END
  END la_input[27]
  PIN la_input[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 736.000 375.730 740.000 ;
    END
  END la_input[28]
  PIN la_input[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.330 736.000 388.610 740.000 ;
    END
  END la_input[29]
  PIN la_input[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.890 736.000 37.170 740.000 ;
    END
  END la_input[2]
  PIN la_input[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.210 736.000 401.490 740.000 ;
    END
  END la_input[30]
  PIN la_input[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 414.090 736.000 414.370 740.000 ;
    END
  END la_input[31]
  PIN la_input[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.430 736.000 427.710 740.000 ;
    END
  END la_input[32]
  PIN la_input[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.310 736.000 440.590 740.000 ;
    END
  END la_input[33]
  PIN la_input[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 453.190 736.000 453.470 740.000 ;
    END
  END la_input[34]
  PIN la_input[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 736.000 466.350 740.000 ;
    END
  END la_input[35]
  PIN la_input[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 736.000 479.690 740.000 ;
    END
  END la_input[36]
  PIN la_input[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.290 736.000 492.570 740.000 ;
    END
  END la_input[37]
  PIN la_input[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 736.000 505.450 740.000 ;
    END
  END la_input[38]
  PIN la_input[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 736.000 518.790 740.000 ;
    END
  END la_input[39]
  PIN la_input[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 736.000 50.510 740.000 ;
    END
  END la_input[3]
  PIN la_input[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 736.000 531.670 740.000 ;
    END
  END la_input[40]
  PIN la_input[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 736.000 544.550 740.000 ;
    END
  END la_input[41]
  PIN la_input[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 736.000 557.430 740.000 ;
    END
  END la_input[42]
  PIN la_input[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 736.000 570.770 740.000 ;
    END
  END la_input[43]
  PIN la_input[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.370 736.000 583.650 740.000 ;
    END
  END la_input[44]
  PIN la_input[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 596.250 736.000 596.530 740.000 ;
    END
  END la_input[45]
  PIN la_input[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 736.000 609.870 740.000 ;
    END
  END la_input[46]
  PIN la_input[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.470 736.000 622.750 740.000 ;
    END
  END la_input[47]
  PIN la_input[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.350 736.000 635.630 740.000 ;
    END
  END la_input[48]
  PIN la_input[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.230 736.000 648.510 740.000 ;
    END
  END la_input[49]
  PIN la_input[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.110 736.000 63.390 740.000 ;
    END
  END la_input[4]
  PIN la_input[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.570 736.000 661.850 740.000 ;
    END
  END la_input[50]
  PIN la_input[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 736.000 674.730 740.000 ;
    END
  END la_input[51]
  PIN la_input[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.330 736.000 687.610 740.000 ;
    END
  END la_input[52]
  PIN la_input[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.670 736.000 700.950 740.000 ;
    END
  END la_input[53]
  PIN la_input[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.550 736.000 713.830 740.000 ;
    END
  END la_input[54]
  PIN la_input[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 726.430 736.000 726.710 740.000 ;
    END
  END la_input[55]
  PIN la_input[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.310 736.000 739.590 740.000 ;
    END
  END la_input[56]
  PIN la_input[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.650 736.000 752.930 740.000 ;
    END
  END la_input[57]
  PIN la_input[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 765.530 736.000 765.810 740.000 ;
    END
  END la_input[58]
  PIN la_input[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.410 736.000 778.690 740.000 ;
    END
  END la_input[59]
  PIN la_input[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 736.000 76.270 740.000 ;
    END
  END la_input[5]
  PIN la_input[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.290 736.000 791.570 740.000 ;
    END
  END la_input[60]
  PIN la_input[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.630 736.000 804.910 740.000 ;
    END
  END la_input[61]
  PIN la_input[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.510 736.000 817.790 740.000 ;
    END
  END la_input[62]
  PIN la_input[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.390 736.000 830.670 740.000 ;
    END
  END la_input[63]
  PIN la_input[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.730 736.000 844.010 740.000 ;
    END
  END la_input[64]
  PIN la_input[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.610 736.000 856.890 740.000 ;
    END
  END la_input[65]
  PIN la_input[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 869.490 736.000 869.770 740.000 ;
    END
  END la_input[66]
  PIN la_input[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.370 736.000 882.650 740.000 ;
    END
  END la_input[67]
  PIN la_input[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.710 736.000 895.990 740.000 ;
    END
  END la_input[68]
  PIN la_input[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.590 736.000 908.870 740.000 ;
    END
  END la_input[69]
  PIN la_input[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 736.000 89.150 740.000 ;
    END
  END la_input[6]
  PIN la_input[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.470 736.000 921.750 740.000 ;
    END
  END la_input[70]
  PIN la_input[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.810 736.000 935.090 740.000 ;
    END
  END la_input[71]
  PIN la_input[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 947.690 736.000 947.970 740.000 ;
    END
  END la_input[72]
  PIN la_input[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 960.570 736.000 960.850 740.000 ;
    END
  END la_input[73]
  PIN la_input[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 973.450 736.000 973.730 740.000 ;
    END
  END la_input[74]
  PIN la_input[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 986.790 736.000 987.070 740.000 ;
    END
  END la_input[75]
  PIN la_input[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.670 736.000 999.950 740.000 ;
    END
  END la_input[76]
  PIN la_input[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.550 736.000 1012.830 740.000 ;
    END
  END la_input[77]
  PIN la_input[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.890 736.000 1026.170 740.000 ;
    END
  END la_input[78]
  PIN la_input[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1038.770 736.000 1039.050 740.000 ;
    END
  END la_input[79]
  PIN la_input[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 736.000 102.490 740.000 ;
    END
  END la_input[7]
  PIN la_input[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.650 736.000 1051.930 740.000 ;
    END
  END la_input[80]
  PIN la_input[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.530 736.000 1064.810 740.000 ;
    END
  END la_input[81]
  PIN la_input[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1077.870 736.000 1078.150 740.000 ;
    END
  END la_input[82]
  PIN la_input[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.750 736.000 1091.030 740.000 ;
    END
  END la_input[83]
  PIN la_input[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1103.630 736.000 1103.910 740.000 ;
    END
  END la_input[84]
  PIN la_input[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.510 736.000 1116.790 740.000 ;
    END
  END la_input[85]
  PIN la_input[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1129.850 736.000 1130.130 740.000 ;
    END
  END la_input[86]
  PIN la_input[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1142.730 736.000 1143.010 740.000 ;
    END
  END la_input[87]
  PIN la_input[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.610 736.000 1155.890 740.000 ;
    END
  END la_input[88]
  PIN la_input[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.950 736.000 1169.230 740.000 ;
    END
  END la_input[89]
  PIN la_input[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 736.000 115.370 740.000 ;
    END
  END la_input[8]
  PIN la_input[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1181.830 736.000 1182.110 740.000 ;
    END
  END la_input[90]
  PIN la_input[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.710 736.000 1194.990 740.000 ;
    END
  END la_input[91]
  PIN la_input[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.590 736.000 1207.870 740.000 ;
    END
  END la_input[92]
  PIN la_input[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.930 736.000 1221.210 740.000 ;
    END
  END la_input[93]
  PIN la_input[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1233.810 736.000 1234.090 740.000 ;
    END
  END la_input[94]
  PIN la_input[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.690 736.000 1246.970 740.000 ;
    END
  END la_input[95]
  PIN la_input[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.030 736.000 1260.310 740.000 ;
    END
  END la_input[96]
  PIN la_input[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1272.910 736.000 1273.190 740.000 ;
    END
  END la_input[97]
  PIN la_input[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.790 736.000 1286.070 740.000 ;
    END
  END la_input[98]
  PIN la_input[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.670 736.000 1298.950 740.000 ;
    END
  END la_input[99]
  PIN la_input[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.970 736.000 128.250 740.000 ;
    END
  END la_input[9]
  PIN la_oenb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 736.000 14.630 740.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1315.230 736.000 1315.510 740.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1328.110 736.000 1328.390 740.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.990 736.000 1341.270 740.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1354.330 736.000 1354.610 740.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.210 736.000 1367.490 740.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1380.090 736.000 1380.370 740.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1392.970 736.000 1393.250 740.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1406.310 736.000 1406.590 740.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.190 736.000 1419.470 740.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.070 736.000 1432.350 740.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.530 736.000 144.810 740.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.410 736.000 1445.690 740.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1458.290 736.000 1458.570 740.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1471.170 736.000 1471.450 740.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.050 736.000 1484.330 740.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.390 736.000 1497.670 740.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1510.270 736.000 1510.550 740.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.150 736.000 1523.430 740.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.490 736.000 1536.770 740.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1549.370 736.000 1549.650 740.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1562.250 736.000 1562.530 740.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.410 736.000 157.690 740.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1575.130 736.000 1575.410 740.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.470 736.000 1588.750 740.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1601.350 736.000 1601.630 740.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1614.230 736.000 1614.510 740.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.110 736.000 1627.390 740.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1640.450 736.000 1640.730 740.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1653.330 736.000 1653.610 740.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1666.210 736.000 1666.490 740.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.290 736.000 170.570 740.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.170 736.000 183.450 740.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 736.000 196.790 740.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.390 736.000 209.670 740.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 736.000 222.550 740.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 736.000 235.890 740.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.490 736.000 248.770 740.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 736.000 261.650 740.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 27.230 736.000 27.510 740.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 736.000 274.530 740.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.590 736.000 287.870 740.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 736.000 300.750 740.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 736.000 313.630 740.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.230 736.000 326.510 740.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.570 736.000 339.850 740.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.450 736.000 352.730 740.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 736.000 365.610 740.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.670 736.000 378.950 740.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 736.000 391.830 740.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 736.000 40.390 740.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.430 736.000 404.710 740.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 417.310 736.000 417.590 740.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.650 736.000 430.930 740.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.530 736.000 443.810 740.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 736.000 456.690 740.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.750 736.000 470.030 740.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 736.000 482.910 740.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.510 736.000 495.790 740.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 736.000 508.670 740.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 736.000 522.010 740.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 736.000 53.730 740.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 736.000 534.890 740.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 736.000 547.770 740.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.830 736.000 561.110 740.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.710 736.000 573.990 740.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 736.000 586.870 740.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.470 736.000 599.750 740.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 736.000 613.090 740.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.690 736.000 625.970 740.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 736.000 638.850 740.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 651.450 736.000 651.730 740.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 66.330 736.000 66.610 740.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.790 736.000 665.070 740.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.670 736.000 677.950 740.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.550 736.000 690.830 740.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 703.890 736.000 704.170 740.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.770 736.000 717.050 740.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 736.000 729.930 740.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.530 736.000 742.810 740.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.870 736.000 756.150 740.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.750 736.000 769.030 740.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 781.630 736.000 781.910 740.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.210 736.000 79.490 740.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.970 736.000 795.250 740.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.850 736.000 808.130 740.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.730 736.000 821.010 740.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.610 736.000 833.890 740.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.950 736.000 847.230 740.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.830 736.000 860.110 740.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.710 736.000 872.990 740.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 886.050 736.000 886.330 740.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.930 736.000 899.210 740.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 911.810 736.000 912.090 740.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 736.000 92.370 740.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.690 736.000 924.970 740.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 938.030 736.000 938.310 740.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 950.910 736.000 951.190 740.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.790 736.000 964.070 740.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.670 736.000 976.950 740.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 990.010 736.000 990.290 740.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.890 736.000 1003.170 740.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.770 736.000 1016.050 740.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1029.110 736.000 1029.390 740.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.990 736.000 1042.270 740.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.430 736.000 105.710 740.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.870 736.000 1055.150 740.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.750 736.000 1068.030 740.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.090 736.000 1081.370 740.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1093.970 736.000 1094.250 740.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1106.850 736.000 1107.130 740.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.190 736.000 1120.470 740.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.070 736.000 1133.350 740.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1145.950 736.000 1146.230 740.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.830 736.000 1159.110 740.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.170 736.000 1172.450 740.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 736.000 118.590 740.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.050 736.000 1185.330 740.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.930 736.000 1198.210 740.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1211.270 736.000 1211.550 740.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.150 736.000 1224.430 740.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.030 736.000 1237.310 740.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.910 736.000 1250.190 740.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.250 736.000 1263.530 740.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1276.130 736.000 1276.410 740.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1289.010 736.000 1289.290 740.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.890 736.000 1302.170 740.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 736.000 131.470 740.000 ;
    END
  END la_oenb[9]
  PIN la_output[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 17.570 736.000 17.850 740.000 ;
    END
  END la_output[0]
  PIN la_output[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1318.450 736.000 1318.730 740.000 ;
    END
  END la_output[100]
  PIN la_output[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1331.330 736.000 1331.610 740.000 ;
    END
  END la_output[101]
  PIN la_output[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.210 736.000 1344.490 740.000 ;
    END
  END la_output[102]
  PIN la_output[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1357.550 736.000 1357.830 740.000 ;
    END
  END la_output[103]
  PIN la_output[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.430 736.000 1370.710 740.000 ;
    END
  END la_output[104]
  PIN la_output[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1383.310 736.000 1383.590 740.000 ;
    END
  END la_output[105]
  PIN la_output[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.190 736.000 1396.470 740.000 ;
    END
  END la_output[106]
  PIN la_output[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.530 736.000 1409.810 740.000 ;
    END
  END la_output[107]
  PIN la_output[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1422.410 736.000 1422.690 740.000 ;
    END
  END la_output[108]
  PIN la_output[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1435.290 736.000 1435.570 740.000 ;
    END
  END la_output[109]
  PIN la_output[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 736.000 148.030 740.000 ;
    END
  END la_output[10]
  PIN la_output[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1448.630 736.000 1448.910 740.000 ;
    END
  END la_output[110]
  PIN la_output[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.510 736.000 1461.790 740.000 ;
    END
  END la_output[111]
  PIN la_output[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.390 736.000 1474.670 740.000 ;
    END
  END la_output[112]
  PIN la_output[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1487.270 736.000 1487.550 740.000 ;
    END
  END la_output[113]
  PIN la_output[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.610 736.000 1500.890 740.000 ;
    END
  END la_output[114]
  PIN la_output[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1513.490 736.000 1513.770 740.000 ;
    END
  END la_output[115]
  PIN la_output[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1526.370 736.000 1526.650 740.000 ;
    END
  END la_output[116]
  PIN la_output[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.710 736.000 1539.990 740.000 ;
    END
  END la_output[117]
  PIN la_output[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1552.590 736.000 1552.870 740.000 ;
    END
  END la_output[118]
  PIN la_output[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1565.470 736.000 1565.750 740.000 ;
    END
  END la_output[119]
  PIN la_output[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 736.000 160.910 740.000 ;
    END
  END la_output[11]
  PIN la_output[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1578.350 736.000 1578.630 740.000 ;
    END
  END la_output[120]
  PIN la_output[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1591.690 736.000 1591.970 740.000 ;
    END
  END la_output[121]
  PIN la_output[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.570 736.000 1604.850 740.000 ;
    END
  END la_output[122]
  PIN la_output[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1617.450 736.000 1617.730 740.000 ;
    END
  END la_output[123]
  PIN la_output[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1630.790 736.000 1631.070 740.000 ;
    END
  END la_output[124]
  PIN la_output[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.670 736.000 1643.950 740.000 ;
    END
  END la_output[125]
  PIN la_output[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1656.550 736.000 1656.830 740.000 ;
    END
  END la_output[126]
  PIN la_output[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.430 736.000 1669.710 740.000 ;
    END
  END la_output[127]
  PIN la_output[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.510 736.000 173.790 740.000 ;
    END
  END la_output[12]
  PIN la_output[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 736.000 186.670 740.000 ;
    END
  END la_output[13]
  PIN la_output[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 736.000 200.010 740.000 ;
    END
  END la_output[14]
  PIN la_output[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 736.000 212.890 740.000 ;
    END
  END la_output[15]
  PIN la_output[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 736.000 225.770 740.000 ;
    END
  END la_output[16]
  PIN la_output[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 736.000 239.110 740.000 ;
    END
  END la_output[17]
  PIN la_output[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.710 736.000 251.990 740.000 ;
    END
  END la_output[18]
  PIN la_output[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.590 736.000 264.870 740.000 ;
    END
  END la_output[19]
  PIN la_output[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 736.000 30.730 740.000 ;
    END
  END la_output[1]
  PIN la_output[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.470 736.000 277.750 740.000 ;
    END
  END la_output[20]
  PIN la_output[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 736.000 291.090 740.000 ;
    END
  END la_output[21]
  PIN la_output[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 736.000 303.970 740.000 ;
    END
  END la_output[22]
  PIN la_output[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.570 736.000 316.850 740.000 ;
    END
  END la_output[23]
  PIN la_output[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 329.910 736.000 330.190 740.000 ;
    END
  END la_output[24]
  PIN la_output[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 736.000 343.070 740.000 ;
    END
  END la_output[25]
  PIN la_output[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.670 736.000 355.950 740.000 ;
    END
  END la_output[26]
  PIN la_output[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.550 736.000 368.830 740.000 ;
    END
  END la_output[27]
  PIN la_output[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 381.890 736.000 382.170 740.000 ;
    END
  END la_output[28]
  PIN la_output[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 736.000 395.050 740.000 ;
    END
  END la_output[29]
  PIN la_output[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.330 736.000 43.610 740.000 ;
    END
  END la_output[2]
  PIN la_output[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 736.000 407.930 740.000 ;
    END
  END la_output[30]
  PIN la_output[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.990 736.000 421.270 740.000 ;
    END
  END la_output[31]
  PIN la_output[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 736.000 434.150 740.000 ;
    END
  END la_output[32]
  PIN la_output[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 736.000 447.030 740.000 ;
    END
  END la_output[33]
  PIN la_output[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.630 736.000 459.910 740.000 ;
    END
  END la_output[34]
  PIN la_output[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.970 736.000 473.250 740.000 ;
    END
  END la_output[35]
  PIN la_output[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.850 736.000 486.130 740.000 ;
    END
  END la_output[36]
  PIN la_output[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 736.000 499.010 740.000 ;
    END
  END la_output[37]
  PIN la_output[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.610 736.000 511.890 740.000 ;
    END
  END la_output[38]
  PIN la_output[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 736.000 525.230 740.000 ;
    END
  END la_output[39]
  PIN la_output[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 56.670 736.000 56.950 740.000 ;
    END
  END la_output[3]
  PIN la_output[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 736.000 538.110 740.000 ;
    END
  END la_output[40]
  PIN la_output[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 736.000 550.990 740.000 ;
    END
  END la_output[41]
  PIN la_output[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.050 736.000 564.330 740.000 ;
    END
  END la_output[42]
  PIN la_output[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.930 736.000 577.210 740.000 ;
    END
  END la_output[43]
  PIN la_output[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 736.000 590.090 740.000 ;
    END
  END la_output[44]
  PIN la_output[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.690 736.000 602.970 740.000 ;
    END
  END la_output[45]
  PIN la_output[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.030 736.000 616.310 740.000 ;
    END
  END la_output[46]
  PIN la_output[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.910 736.000 629.190 740.000 ;
    END
  END la_output[47]
  PIN la_output[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 736.000 642.070 740.000 ;
    END
  END la_output[48]
  PIN la_output[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.130 736.000 655.410 740.000 ;
    END
  END la_output[49]
  PIN la_output[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 736.000 69.830 740.000 ;
    END
  END la_output[4]
  PIN la_output[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.010 736.000 668.290 740.000 ;
    END
  END la_output[50]
  PIN la_output[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.890 736.000 681.170 740.000 ;
    END
  END la_output[51]
  PIN la_output[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 693.770 736.000 694.050 740.000 ;
    END
  END la_output[52]
  PIN la_output[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.110 736.000 707.390 740.000 ;
    END
  END la_output[53]
  PIN la_output[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.990 736.000 720.270 740.000 ;
    END
  END la_output[54]
  PIN la_output[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 732.870 736.000 733.150 740.000 ;
    END
  END la_output[55]
  PIN la_output[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.210 736.000 746.490 740.000 ;
    END
  END la_output[56]
  PIN la_output[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 736.000 759.370 740.000 ;
    END
  END la_output[57]
  PIN la_output[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.970 736.000 772.250 740.000 ;
    END
  END la_output[58]
  PIN la_output[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.850 736.000 785.130 740.000 ;
    END
  END la_output[59]
  PIN la_output[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 736.000 82.710 740.000 ;
    END
  END la_output[5]
  PIN la_output[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.190 736.000 798.470 740.000 ;
    END
  END la_output[60]
  PIN la_output[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.070 736.000 811.350 740.000 ;
    END
  END la_output[61]
  PIN la_output[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 823.950 736.000 824.230 740.000 ;
    END
  END la_output[62]
  PIN la_output[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.830 736.000 837.110 740.000 ;
    END
  END la_output[63]
  PIN la_output[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 736.000 850.450 740.000 ;
    END
  END la_output[64]
  PIN la_output[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 863.050 736.000 863.330 740.000 ;
    END
  END la_output[65]
  PIN la_output[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.930 736.000 876.210 740.000 ;
    END
  END la_output[66]
  PIN la_output[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.270 736.000 889.550 740.000 ;
    END
  END la_output[67]
  PIN la_output[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 902.150 736.000 902.430 740.000 ;
    END
  END la_output[68]
  PIN la_output[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.030 736.000 915.310 740.000 ;
    END
  END la_output[69]
  PIN la_output[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 736.000 96.050 740.000 ;
    END
  END la_output[6]
  PIN la_output[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 927.910 736.000 928.190 740.000 ;
    END
  END la_output[70]
  PIN la_output[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 941.250 736.000 941.530 740.000 ;
    END
  END la_output[71]
  PIN la_output[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.130 736.000 954.410 740.000 ;
    END
  END la_output[72]
  PIN la_output[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.010 736.000 967.290 740.000 ;
    END
  END la_output[73]
  PIN la_output[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 980.350 736.000 980.630 740.000 ;
    END
  END la_output[74]
  PIN la_output[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.230 736.000 993.510 740.000 ;
    END
  END la_output[75]
  PIN la_output[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1006.110 736.000 1006.390 740.000 ;
    END
  END la_output[76]
  PIN la_output[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1018.990 736.000 1019.270 740.000 ;
    END
  END la_output[77]
  PIN la_output[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1032.330 736.000 1032.610 740.000 ;
    END
  END la_output[78]
  PIN la_output[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1045.210 736.000 1045.490 740.000 ;
    END
  END la_output[79]
  PIN la_output[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 736.000 108.930 740.000 ;
    END
  END la_output[7]
  PIN la_output[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.090 736.000 1058.370 740.000 ;
    END
  END la_output[80]
  PIN la_output[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1071.430 736.000 1071.710 740.000 ;
    END
  END la_output[81]
  PIN la_output[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.310 736.000 1084.590 740.000 ;
    END
  END la_output[82]
  PIN la_output[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.190 736.000 1097.470 740.000 ;
    END
  END la_output[83]
  PIN la_output[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1110.070 736.000 1110.350 740.000 ;
    END
  END la_output[84]
  PIN la_output[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1123.410 736.000 1123.690 740.000 ;
    END
  END la_output[85]
  PIN la_output[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.290 736.000 1136.570 740.000 ;
    END
  END la_output[86]
  PIN la_output[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.170 736.000 1149.450 740.000 ;
    END
  END la_output[87]
  PIN la_output[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1162.050 736.000 1162.330 740.000 ;
    END
  END la_output[88]
  PIN la_output[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.390 736.000 1175.670 740.000 ;
    END
  END la_output[89]
  PIN la_output[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.530 736.000 121.810 740.000 ;
    END
  END la_output[8]
  PIN la_output[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.270 736.000 1188.550 740.000 ;
    END
  END la_output[90]
  PIN la_output[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.150 736.000 1201.430 740.000 ;
    END
  END la_output[91]
  PIN la_output[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.490 736.000 1214.770 740.000 ;
    END
  END la_output[92]
  PIN la_output[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.370 736.000 1227.650 740.000 ;
    END
  END la_output[93]
  PIN la_output[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1240.250 736.000 1240.530 740.000 ;
    END
  END la_output[94]
  PIN la_output[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1253.130 736.000 1253.410 740.000 ;
    END
  END la_output[95]
  PIN la_output[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1266.470 736.000 1266.750 740.000 ;
    END
  END la_output[96]
  PIN la_output[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.350 736.000 1279.630 740.000 ;
    END
  END la_output[97]
  PIN la_output[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1292.230 736.000 1292.510 740.000 ;
    END
  END la_output[98]
  PIN la_output[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1305.570 736.000 1305.850 740.000 ;
    END
  END la_output[99]
  PIN la_output[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 736.000 134.690 740.000 ;
    END
  END la_output[9]
  PIN mgmt_soc_dff_A[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.330 0.000 1722.610 4.000 ;
    END
  END mgmt_soc_dff_A[0]
  PIN mgmt_soc_dff_A[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 83.000 2000.000 83.600 ;
    END
  END mgmt_soc_dff_A[1]
  PIN mgmt_soc_dff_A[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1755.910 0.000 1756.190 4.000 ;
    END
  END mgmt_soc_dff_A[2]
  PIN mgmt_soc_dff_A[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.800 4.000 515.400 ;
    END
  END mgmt_soc_dff_A[3]
  PIN mgmt_soc_dff_A[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 184.320 2000.000 184.920 ;
    END
  END mgmt_soc_dff_A[4]
  PIN mgmt_soc_dff_A[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1952.330 736.000 1952.610 740.000 ;
    END
  END mgmt_soc_dff_A[5]
  PIN mgmt_soc_dff_A[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 251.640 2000.000 252.240 ;
    END
  END mgmt_soc_dff_A[6]
  PIN mgmt_soc_dff_A[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.080 4.000 563.680 ;
    END
  END mgmt_soc_dff_A[7]
  PIN mgmt_soc_dff_Di[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.790 736.000 1930.070 740.000 ;
    END
  END mgmt_soc_dff_Di[0]
  PIN mgmt_soc_dff_Di[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 352.280 2000.000 352.880 ;
    END
  END mgmt_soc_dff_Di[10]
  PIN mgmt_soc_dff_Di[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END mgmt_soc_dff_Di[11]
  PIN mgmt_soc_dff_Di[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1972.110 736.000 1972.390 740.000 ;
    END
  END mgmt_soc_dff_Di[12]
  PIN mgmt_soc_dff_Di[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.120 4.000 599.720 ;
    END
  END mgmt_soc_dff_Di[13]
  PIN mgmt_soc_dff_Di[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 419.600 2000.000 420.200 ;
    END
  END mgmt_soc_dff_Di[14]
  PIN mgmt_soc_dff_Di[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 611.360 4.000 611.960 ;
    END
  END mgmt_soc_dff_Di[15]
  PIN mgmt_soc_dff_Di[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 635.840 4.000 636.440 ;
    END
  END mgmt_soc_dff_Di[16]
  PIN mgmt_soc_dff_Di[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 452.920 2000.000 453.520 ;
    END
  END mgmt_soc_dff_Di[17]
  PIN mgmt_soc_dff_Di[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 486.920 2000.000 487.520 ;
    END
  END mgmt_soc_dff_Di[18]
  PIN mgmt_soc_dff_Di[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.690 0.000 1890.970 4.000 ;
    END
  END mgmt_soc_dff_Di[19]
  PIN mgmt_soc_dff_Di[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 117.000 2000.000 117.600 ;
    END
  END mgmt_soc_dff_Di[1]
  PIN mgmt_soc_dff_Di[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1978.550 736.000 1978.830 740.000 ;
    END
  END mgmt_soc_dff_Di[20]
  PIN mgmt_soc_dff_Di[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1924.270 0.000 1924.550 4.000 ;
    END
  END mgmt_soc_dff_Di[21]
  PIN mgmt_soc_dff_Di[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.880 4.000 672.480 ;
    END
  END mgmt_soc_dff_Di[22]
  PIN mgmt_soc_dff_Di[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END mgmt_soc_dff_Di[23]
  PIN mgmt_soc_dff_Di[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1940.830 0.000 1941.110 4.000 ;
    END
  END mgmt_soc_dff_Di[24]
  PIN mgmt_soc_dff_Di[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.210 736.000 1988.490 740.000 ;
    END
  END mgmt_soc_dff_Di[25]
  PIN mgmt_soc_dff_Di[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1957.850 0.000 1958.130 4.000 ;
    END
  END mgmt_soc_dff_Di[26]
  PIN mgmt_soc_dff_Di[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.650 736.000 1994.930 740.000 ;
    END
  END mgmt_soc_dff_Di[27]
  PIN mgmt_soc_dff_Di[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1991.430 0.000 1991.710 4.000 ;
    END
  END mgmt_soc_dff_Di[28]
  PIN mgmt_soc_dff_Di[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 688.880 2000.000 689.480 ;
    END
  END mgmt_soc_dff_Di[29]
  PIN mgmt_soc_dff_Di[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1936.230 736.000 1936.510 740.000 ;
    END
  END mgmt_soc_dff_Di[2]
  PIN mgmt_soc_dff_Di[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 696.360 4.000 696.960 ;
    END
  END mgmt_soc_dff_Di[30]
  PIN mgmt_soc_dff_Di[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END mgmt_soc_dff_Di[31]
  PIN mgmt_soc_dff_Di[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1789.950 0.000 1790.230 4.000 ;
    END
  END mgmt_soc_dff_Di[3]
  PIN mgmt_soc_dff_Di[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 217.640 2000.000 218.240 ;
    END
  END mgmt_soc_dff_Di[4]
  PIN mgmt_soc_dff_Di[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 538.600 4.000 539.200 ;
    END
  END mgmt_soc_dff_Di[5]
  PIN mgmt_soc_dff_Di[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1840.090 0.000 1840.370 4.000 ;
    END
  END mgmt_soc_dff_Di[6]
  PIN mgmt_soc_dff_Di[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.230 736.000 1959.510 740.000 ;
    END
  END mgmt_soc_dff_Di[7]
  PIN mgmt_soc_dff_Di[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.670 736.000 1965.950 740.000 ;
    END
  END mgmt_soc_dff_Di[8]
  PIN mgmt_soc_dff_Di[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 318.960 2000.000 319.560 ;
    END
  END mgmt_soc_dff_Di[9]
  PIN mgmt_soc_dff_Do[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 16.360 2000.000 16.960 ;
    END
  END mgmt_soc_dff_Do[0]
  PIN mgmt_soc_dff_Do[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1968.890 736.000 1969.170 740.000 ;
    END
  END mgmt_soc_dff_Do[10]
  PIN mgmt_soc_dff_Do[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 587.560 4.000 588.160 ;
    END
  END mgmt_soc_dff_Do[11]
  PIN mgmt_soc_dff_Do[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 386.280 2000.000 386.880 ;
    END
  END mgmt_soc_dff_Do[12]
  PIN mgmt_soc_dff_Do[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1975.330 736.000 1975.610 740.000 ;
    END
  END mgmt_soc_dff_Do[13]
  PIN mgmt_soc_dff_Do[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1873.670 0.000 1873.950 4.000 ;
    END
  END mgmt_soc_dff_Do[14]
  PIN mgmt_soc_dff_Do[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 623.600 4.000 624.200 ;
    END
  END mgmt_soc_dff_Do[15]
  PIN mgmt_soc_dff_Do[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 648.080 4.000 648.680 ;
    END
  END mgmt_soc_dff_Do[16]
  PIN mgmt_soc_dff_Do[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 660.320 4.000 660.920 ;
    END
  END mgmt_soc_dff_Do[17]
  PIN mgmt_soc_dff_Do[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 520.240 2000.000 520.840 ;
    END
  END mgmt_soc_dff_Do[18]
  PIN mgmt_soc_dff_Do[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1907.250 0.000 1907.530 4.000 ;
    END
  END mgmt_soc_dff_Do[19]
  PIN mgmt_soc_dff_Do[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1933.010 736.000 1933.290 740.000 ;
    END
  END mgmt_soc_dff_Do[1]
  PIN mgmt_soc_dff_Do[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 554.240 2000.000 554.840 ;
    END
  END mgmt_soc_dff_Do[20]
  PIN mgmt_soc_dff_Do[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 587.560 2000.000 588.160 ;
    END
  END mgmt_soc_dff_Do[21]
  PIN mgmt_soc_dff_Do[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1981.770 736.000 1982.050 740.000 ;
    END
  END mgmt_soc_dff_Do[22]
  PIN mgmt_soc_dff_Do[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 621.560 2000.000 622.160 ;
    END
  END mgmt_soc_dff_Do[23]
  PIN mgmt_soc_dff_Do[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1984.990 736.000 1985.270 740.000 ;
    END
  END mgmt_soc_dff_Do[24]
  PIN mgmt_soc_dff_Do[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1991.430 736.000 1991.710 740.000 ;
    END
  END mgmt_soc_dff_Do[25]
  PIN mgmt_soc_dff_Do[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 654.880 2000.000 655.480 ;
    END
  END mgmt_soc_dff_Do[26]
  PIN mgmt_soc_dff_Do[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1974.410 0.000 1974.690 4.000 ;
    END
  END mgmt_soc_dff_Do[27]
  PIN mgmt_soc_dff_Do[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1997.870 736.000 1998.150 740.000 ;
    END
  END mgmt_soc_dff_Do[28]
  PIN mgmt_soc_dff_Do[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 722.200 2000.000 722.800 ;
    END
  END mgmt_soc_dff_Do[29]
  PIN mgmt_soc_dff_Do[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 502.560 4.000 503.160 ;
    END
  END mgmt_soc_dff_Do[2]
  PIN mgmt_soc_dff_Do[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 708.600 4.000 709.200 ;
    END
  END mgmt_soc_dff_Do[30]
  PIN mgmt_soc_dff_Do[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 733.080 4.000 733.680 ;
    END
  END mgmt_soc_dff_Do[31]
  PIN mgmt_soc_dff_Do[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 526.360 4.000 526.960 ;
    END
  END mgmt_soc_dff_Do[3]
  PIN mgmt_soc_dff_Do[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1945.890 736.000 1946.170 740.000 ;
    END
  END mgmt_soc_dff_Do[4]
  PIN mgmt_soc_dff_Do[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1823.530 0.000 1823.810 4.000 ;
    END
  END mgmt_soc_dff_Do[5]
  PIN mgmt_soc_dff_Do[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1956.010 736.000 1956.290 740.000 ;
    END
  END mgmt_soc_dff_Do[6]
  PIN mgmt_soc_dff_Do[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1962.450 736.000 1962.730 740.000 ;
    END
  END mgmt_soc_dff_Do[7]
  PIN mgmt_soc_dff_Do[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 284.960 2000.000 285.560 ;
    END
  END mgmt_soc_dff_Do[8]
  PIN mgmt_soc_dff_Do[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1857.110 0.000 1857.390 4.000 ;
    END
  END mgmt_soc_dff_Do[9]
  PIN mgmt_soc_dff_EN
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.040 4.000 442.640 ;
    END
  END mgmt_soc_dff_EN
  PIN mgmt_soc_dff_WE[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 490.320 4.000 490.920 ;
    END
  END mgmt_soc_dff_WE[0]
  PIN mgmt_soc_dff_WE[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1739.350 0.000 1739.630 4.000 ;
    END
  END mgmt_soc_dff_WE[1]
  PIN mgmt_soc_dff_WE[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1939.450 736.000 1939.730 740.000 ;
    END
  END mgmt_soc_dff_WE[2]
  PIN mgmt_soc_dff_WE[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1806.510 0.000 1806.790 4.000 ;
    END
  END mgmt_soc_dff_WE[3]
  PIN mprj_ack_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 417.560 4.000 418.160 ;
    END
  END mprj_ack_i
  PIN mprj_adr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1682.770 736.000 1683.050 740.000 ;
    END
  END mprj_adr_o[0]
  PIN mprj_adr_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.510 736.000 1760.790 740.000 ;
    END
  END mprj_adr_o[10]
  PIN mprj_adr_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1766.950 736.000 1767.230 740.000 ;
    END
  END mprj_adr_o[11]
  PIN mprj_adr_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1773.850 736.000 1774.130 740.000 ;
    END
  END mprj_adr_o[12]
  PIN mprj_adr_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1780.290 736.000 1780.570 740.000 ;
    END
  END mprj_adr_o[13]
  PIN mprj_adr_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1786.730 736.000 1787.010 740.000 ;
    END
  END mprj_adr_o[14]
  PIN mprj_adr_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.170 736.000 1793.450 740.000 ;
    END
  END mprj_adr_o[15]
  PIN mprj_adr_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.610 736.000 1799.890 740.000 ;
    END
  END mprj_adr_o[16]
  PIN mprj_adr_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1806.050 736.000 1806.330 740.000 ;
    END
  END mprj_adr_o[17]
  PIN mprj_adr_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1812.490 736.000 1812.770 740.000 ;
    END
  END mprj_adr_o[18]
  PIN mprj_adr_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1819.390 736.000 1819.670 740.000 ;
    END
  END mprj_adr_o[19]
  PIN mprj_adr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1692.430 736.000 1692.710 740.000 ;
    END
  END mprj_adr_o[1]
  PIN mprj_adr_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1825.830 736.000 1826.110 740.000 ;
    END
  END mprj_adr_o[20]
  PIN mprj_adr_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1832.270 736.000 1832.550 740.000 ;
    END
  END mprj_adr_o[21]
  PIN mprj_adr_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1838.710 736.000 1838.990 740.000 ;
    END
  END mprj_adr_o[22]
  PIN mprj_adr_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.150 736.000 1845.430 740.000 ;
    END
  END mprj_adr_o[23]
  PIN mprj_adr_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1851.590 736.000 1851.870 740.000 ;
    END
  END mprj_adr_o[24]
  PIN mprj_adr_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.030 736.000 1858.310 740.000 ;
    END
  END mprj_adr_o[25]
  PIN mprj_adr_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.930 736.000 1865.210 740.000 ;
    END
  END mprj_adr_o[26]
  PIN mprj_adr_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1871.370 736.000 1871.650 740.000 ;
    END
  END mprj_adr_o[27]
  PIN mprj_adr_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1877.810 736.000 1878.090 740.000 ;
    END
  END mprj_adr_o[28]
  PIN mprj_adr_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1884.250 736.000 1884.530 740.000 ;
    END
  END mprj_adr_o[29]
  PIN mprj_adr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1702.090 736.000 1702.370 740.000 ;
    END
  END mprj_adr_o[2]
  PIN mprj_adr_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1890.690 736.000 1890.970 740.000 ;
    END
  END mprj_adr_o[30]
  PIN mprj_adr_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1897.130 736.000 1897.410 740.000 ;
    END
  END mprj_adr_o[31]
  PIN mprj_adr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1711.750 736.000 1712.030 740.000 ;
    END
  END mprj_adr_o[3]
  PIN mprj_adr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.410 736.000 1721.690 740.000 ;
    END
  END mprj_adr_o[4]
  PIN mprj_adr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.310 736.000 1728.590 740.000 ;
    END
  END mprj_adr_o[5]
  PIN mprj_adr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.750 736.000 1735.030 740.000 ;
    END
  END mprj_adr_o[6]
  PIN mprj_adr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1741.190 736.000 1741.470 740.000 ;
    END
  END mprj_adr_o[7]
  PIN mprj_adr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1747.630 736.000 1747.910 740.000 ;
    END
  END mprj_adr_o[8]
  PIN mprj_adr_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.070 736.000 1754.350 740.000 ;
    END
  END mprj_adr_o[9]
  PIN mprj_cyc_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1672.650 736.000 1672.930 740.000 ;
    END
  END mprj_cyc_o
  PIN mprj_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.280 4.000 29.880 ;
    END
  END mprj_dat_i[0]
  PIN mprj_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END mprj_dat_i[10]
  PIN mprj_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 162.560 4.000 163.160 ;
    END
  END mprj_dat_i[11]
  PIN mprj_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END mprj_dat_i[12]
  PIN mprj_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END mprj_dat_i[13]
  PIN mprj_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END mprj_dat_i[14]
  PIN mprj_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 211.520 4.000 212.120 ;
    END
  END mprj_dat_i[15]
  PIN mprj_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.760 4.000 224.360 ;
    END
  END mprj_dat_i[16]
  PIN mprj_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END mprj_dat_i[17]
  PIN mprj_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END mprj_dat_i[18]
  PIN mprj_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END mprj_dat_i[19]
  PIN mprj_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END mprj_dat_i[1]
  PIN mprj_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END mprj_dat_i[20]
  PIN mprj_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END mprj_dat_i[21]
  PIN mprj_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END mprj_dat_i[22]
  PIN mprj_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.080 4.000 308.680 ;
    END
  END mprj_dat_i[23]
  PIN mprj_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 320.320 4.000 320.920 ;
    END
  END mprj_dat_i[24]
  PIN mprj_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 332.560 4.000 333.160 ;
    END
  END mprj_dat_i[25]
  PIN mprj_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.800 4.000 345.400 ;
    END
  END mprj_dat_i[26]
  PIN mprj_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END mprj_dat_i[27]
  PIN mprj_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.280 4.000 369.880 ;
    END
  END mprj_dat_i[28]
  PIN mprj_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END mprj_dat_i[29]
  PIN mprj_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END mprj_dat_i[2]
  PIN mprj_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 393.080 4.000 393.680 ;
    END
  END mprj_dat_i[30]
  PIN mprj_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END mprj_dat_i[31]
  PIN mprj_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.000 4.000 66.600 ;
    END
  END mprj_dat_i[3]
  PIN mprj_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END mprj_dat_i[4]
  PIN mprj_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 89.800 4.000 90.400 ;
    END
  END mprj_dat_i[5]
  PIN mprj_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END mprj_dat_i[6]
  PIN mprj_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.280 4.000 114.880 ;
    END
  END mprj_dat_i[7]
  PIN mprj_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END mprj_dat_i[8]
  PIN mprj_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END mprj_dat_i[9]
  PIN mprj_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.990 736.000 1686.270 740.000 ;
    END
  END mprj_dat_o[0]
  PIN mprj_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1763.730 736.000 1764.010 740.000 ;
    END
  END mprj_dat_o[10]
  PIN mprj_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.630 736.000 1770.910 740.000 ;
    END
  END mprj_dat_o[11]
  PIN mprj_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1777.070 736.000 1777.350 740.000 ;
    END
  END mprj_dat_o[12]
  PIN mprj_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1783.510 736.000 1783.790 740.000 ;
    END
  END mprj_dat_o[13]
  PIN mprj_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1789.950 736.000 1790.230 740.000 ;
    END
  END mprj_dat_o[14]
  PIN mprj_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1796.390 736.000 1796.670 740.000 ;
    END
  END mprj_dat_o[15]
  PIN mprj_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1802.830 736.000 1803.110 740.000 ;
    END
  END mprj_dat_o[16]
  PIN mprj_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1809.270 736.000 1809.550 740.000 ;
    END
  END mprj_dat_o[17]
  PIN mprj_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1816.170 736.000 1816.450 740.000 ;
    END
  END mprj_dat_o[18]
  PIN mprj_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.610 736.000 1822.890 740.000 ;
    END
  END mprj_dat_o[19]
  PIN mprj_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1695.650 736.000 1695.930 740.000 ;
    END
  END mprj_dat_o[1]
  PIN mprj_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1829.050 736.000 1829.330 740.000 ;
    END
  END mprj_dat_o[20]
  PIN mprj_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1835.490 736.000 1835.770 740.000 ;
    END
  END mprj_dat_o[21]
  PIN mprj_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1841.930 736.000 1842.210 740.000 ;
    END
  END mprj_dat_o[22]
  PIN mprj_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1848.370 736.000 1848.650 740.000 ;
    END
  END mprj_dat_o[23]
  PIN mprj_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.810 736.000 1855.090 740.000 ;
    END
  END mprj_dat_o[24]
  PIN mprj_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1861.250 736.000 1861.530 740.000 ;
    END
  END mprj_dat_o[25]
  PIN mprj_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1868.150 736.000 1868.430 740.000 ;
    END
  END mprj_dat_o[26]
  PIN mprj_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1874.590 736.000 1874.870 740.000 ;
    END
  END mprj_dat_o[27]
  PIN mprj_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.030 736.000 1881.310 740.000 ;
    END
  END mprj_dat_o[28]
  PIN mprj_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.470 736.000 1887.750 740.000 ;
    END
  END mprj_dat_o[29]
  PIN mprj_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1705.310 736.000 1705.590 740.000 ;
    END
  END mprj_dat_o[2]
  PIN mprj_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1893.910 736.000 1894.190 740.000 ;
    END
  END mprj_dat_o[30]
  PIN mprj_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1900.350 736.000 1900.630 740.000 ;
    END
  END mprj_dat_o[31]
  PIN mprj_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1714.970 736.000 1715.250 740.000 ;
    END
  END mprj_dat_o[3]
  PIN mprj_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1725.090 736.000 1725.370 740.000 ;
    END
  END mprj_dat_o[4]
  PIN mprj_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1731.530 736.000 1731.810 740.000 ;
    END
  END mprj_dat_o[5]
  PIN mprj_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1737.970 736.000 1738.250 740.000 ;
    END
  END mprj_dat_o[6]
  PIN mprj_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1744.410 736.000 1744.690 740.000 ;
    END
  END mprj_dat_o[7]
  PIN mprj_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1750.850 736.000 1751.130 740.000 ;
    END
  END mprj_dat_o[8]
  PIN mprj_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1757.290 736.000 1757.570 740.000 ;
    END
  END mprj_dat_o[9]
  PIN mprj_sel_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1689.210 736.000 1689.490 740.000 ;
    END
  END mprj_sel_o[0]
  PIN mprj_sel_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1698.870 736.000 1699.150 740.000 ;
    END
  END mprj_sel_o[1]
  PIN mprj_sel_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1708.530 736.000 1708.810 740.000 ;
    END
  END mprj_sel_o[2]
  PIN mprj_sel_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1718.190 736.000 1718.470 740.000 ;
    END
  END mprj_sel_o[3]
  PIN mprj_stb_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1676.330 736.000 1676.610 740.000 ;
    END
  END mprj_stb_o
  PIN mprj_wb_iena
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.570 736.000 1903.850 740.000 ;
    END
  END mprj_wb_iena
  PIN mprj_we_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.550 736.000 1679.830 740.000 ;
    END
  END mprj_we_o
  PIN qspi_enabled
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 0.000 294.310 4.000 ;
    END
  END qspi_enabled
  PIN serial_rx
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 453.600 4.000 454.200 ;
    END
  END serial_rx
  PIN serial_tx
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END serial_tx
  PIN spi_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.350 736.000 1923.630 740.000 ;
    END
  END spi_clk
  PIN spi_cs_n
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1926.570 736.000 1926.850 740.000 ;
    END
  END spi_cs_n
  PIN spi_enabled
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.590 0.000 1621.870 4.000 ;
    END
  END spi_enabled
  PIN spi_miso
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1705.770 0.000 1706.050 4.000 ;
    END
  END spi_miso
  PIN spi_mosi
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.080 4.000 478.680 ;
    END
  END spi_mosi
  PIN spi_sdoenb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1638.610 0.000 1638.890 4.000 ;
    END
  END spi_sdoenb
  PIN sram_ro_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.950 0.000 916.230 4.000 ;
    END
  END sram_ro_addr[0]
  PIN sram_ro_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.510 0.000 932.790 4.000 ;
    END
  END sram_ro_addr[1]
  PIN sram_ro_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 949.530 0.000 949.810 4.000 ;
    END
  END sram_ro_addr[2]
  PIN sram_ro_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 966.090 0.000 966.370 4.000 ;
    END
  END sram_ro_addr[3]
  PIN sram_ro_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.110 0.000 983.390 4.000 ;
    END
  END sram_ro_addr[4]
  PIN sram_ro_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 999.670 0.000 999.950 4.000 ;
    END
  END sram_ro_addr[5]
  PIN sram_ro_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1016.690 0.000 1016.970 4.000 ;
    END
  END sram_ro_addr[6]
  PIN sram_ro_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1033.250 0.000 1033.530 4.000 ;
    END
  END sram_ro_addr[7]
  PIN sram_ro_clk
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 881.910 0.000 882.190 4.000 ;
    END
  END sram_ro_clk
  PIN sram_ro_csb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.930 0.000 899.210 4.000 ;
    END
  END sram_ro_csb
  PIN sram_ro_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.270 0.000 1050.550 4.000 ;
    END
  END sram_ro_data[0]
  PIN sram_ro_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.170 0.000 1218.450 4.000 ;
    END
  END sram_ro_data[10]
  PIN sram_ro_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1235.190 0.000 1235.470 4.000 ;
    END
  END sram_ro_data[11]
  PIN sram_ro_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1251.750 0.000 1252.030 4.000 ;
    END
  END sram_ro_data[12]
  PIN sram_ro_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.770 0.000 1269.050 4.000 ;
    END
  END sram_ro_data[13]
  PIN sram_ro_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.330 0.000 1285.610 4.000 ;
    END
  END sram_ro_data[14]
  PIN sram_ro_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1302.350 0.000 1302.630 4.000 ;
    END
  END sram_ro_data[15]
  PIN sram_ro_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1318.910 0.000 1319.190 4.000 ;
    END
  END sram_ro_data[16]
  PIN sram_ro_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.930 0.000 1336.210 4.000 ;
    END
  END sram_ro_data[17]
  PIN sram_ro_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1352.950 0.000 1353.230 4.000 ;
    END
  END sram_ro_data[18]
  PIN sram_ro_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1369.510 0.000 1369.790 4.000 ;
    END
  END sram_ro_data[19]
  PIN sram_ro_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.830 0.000 1067.110 4.000 ;
    END
  END sram_ro_data[1]
  PIN sram_ro_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1386.530 0.000 1386.810 4.000 ;
    END
  END sram_ro_data[20]
  PIN sram_ro_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.090 0.000 1403.370 4.000 ;
    END
  END sram_ro_data[21]
  PIN sram_ro_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.110 0.000 1420.390 4.000 ;
    END
  END sram_ro_data[22]
  PIN sram_ro_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.670 0.000 1436.950 4.000 ;
    END
  END sram_ro_data[23]
  PIN sram_ro_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.690 0.000 1453.970 4.000 ;
    END
  END sram_ro_data[24]
  PIN sram_ro_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1470.250 0.000 1470.530 4.000 ;
    END
  END sram_ro_data[25]
  PIN sram_ro_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1487.270 0.000 1487.550 4.000 ;
    END
  END sram_ro_data[26]
  PIN sram_ro_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.830 0.000 1504.110 4.000 ;
    END
  END sram_ro_data[27]
  PIN sram_ro_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1520.850 0.000 1521.130 4.000 ;
    END
  END sram_ro_data[28]
  PIN sram_ro_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1537.410 0.000 1537.690 4.000 ;
    END
  END sram_ro_data[29]
  PIN sram_ro_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.850 0.000 1084.130 4.000 ;
    END
  END sram_ro_data[2]
  PIN sram_ro_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1554.430 0.000 1554.710 4.000 ;
    END
  END sram_ro_data[30]
  PIN sram_ro_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1571.450 0.000 1571.730 4.000 ;
    END
  END sram_ro_data[31]
  PIN sram_ro_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1100.410 0.000 1100.690 4.000 ;
    END
  END sram_ro_data[3]
  PIN sram_ro_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1117.430 0.000 1117.710 4.000 ;
    END
  END sram_ro_data[4]
  PIN sram_ro_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1134.450 0.000 1134.730 4.000 ;
    END
  END sram_ro_data[5]
  PIN sram_ro_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1151.010 0.000 1151.290 4.000 ;
    END
  END sram_ro_data[6]
  PIN sram_ro_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1168.030 0.000 1168.310 4.000 ;
    END
  END sram_ro_data[7]
  PIN sram_ro_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.590 0.000 1184.870 4.000 ;
    END
  END sram_ro_data[8]
  PIN sram_ro_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1201.610 0.000 1201.890 4.000 ;
    END
  END sram_ro_data[9]
  PIN trap
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1655.170 0.000 1655.450 4.000 ;
    END
  END trap
  PIN uart_enabled
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1672.190 0.000 1672.470 4.000 ;
    END
  END uart_enabled
  PIN user_irq[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 49.680 2000.000 50.280 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 1996.000 150.320 2000.000 150.920 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1772.930 0.000 1773.210 4.000 ;
    END
  END user_irq[2]
  PIN user_irq[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1942.670 736.000 1942.950 740.000 ;
    END
  END user_irq[3]
  PIN user_irq[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1949.110 736.000 1949.390 740.000 ;
    END
  END user_irq[4]
  PIN user_irq[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.840 4.000 551.440 ;
    END
  END user_irq[5]
  PIN user_irq_ena[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1906.790 736.000 1907.070 740.000 ;
    END
  END user_irq_ena[0]
  PIN user_irq_ena[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1910.470 736.000 1910.750 740.000 ;
    END
  END user_irq_ena[1]
  PIN user_irq_ena[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1913.690 736.000 1913.970 740.000 ;
    END
  END user_irq_ena[2]
  OBS
      LAYER li1 ;
        RECT 10.120 10.795 1989.500 729.045 ;
      LAYER met1 ;
        RECT 1.450 6.500 1998.170 732.660 ;
      LAYER met2 ;
        RECT 2.030 735.720 4.410 736.170 ;
        RECT 5.250 735.720 7.630 736.170 ;
        RECT 8.470 735.720 10.850 736.170 ;
        RECT 11.690 735.720 14.070 736.170 ;
        RECT 14.910 735.720 17.290 736.170 ;
        RECT 18.130 735.720 20.510 736.170 ;
        RECT 21.350 735.720 23.730 736.170 ;
        RECT 24.570 735.720 26.950 736.170 ;
        RECT 27.790 735.720 30.170 736.170 ;
        RECT 31.010 735.720 33.390 736.170 ;
        RECT 34.230 735.720 36.610 736.170 ;
        RECT 37.450 735.720 39.830 736.170 ;
        RECT 40.670 735.720 43.050 736.170 ;
        RECT 43.890 735.720 46.270 736.170 ;
        RECT 47.110 735.720 49.950 736.170 ;
        RECT 50.790 735.720 53.170 736.170 ;
        RECT 54.010 735.720 56.390 736.170 ;
        RECT 57.230 735.720 59.610 736.170 ;
        RECT 60.450 735.720 62.830 736.170 ;
        RECT 63.670 735.720 66.050 736.170 ;
        RECT 66.890 735.720 69.270 736.170 ;
        RECT 70.110 735.720 72.490 736.170 ;
        RECT 73.330 735.720 75.710 736.170 ;
        RECT 76.550 735.720 78.930 736.170 ;
        RECT 79.770 735.720 82.150 736.170 ;
        RECT 82.990 735.720 85.370 736.170 ;
        RECT 86.210 735.720 88.590 736.170 ;
        RECT 89.430 735.720 91.810 736.170 ;
        RECT 92.650 735.720 95.490 736.170 ;
        RECT 96.330 735.720 98.710 736.170 ;
        RECT 99.550 735.720 101.930 736.170 ;
        RECT 102.770 735.720 105.150 736.170 ;
        RECT 105.990 735.720 108.370 736.170 ;
        RECT 109.210 735.720 111.590 736.170 ;
        RECT 112.430 735.720 114.810 736.170 ;
        RECT 115.650 735.720 118.030 736.170 ;
        RECT 118.870 735.720 121.250 736.170 ;
        RECT 122.090 735.720 124.470 736.170 ;
        RECT 125.310 735.720 127.690 736.170 ;
        RECT 128.530 735.720 130.910 736.170 ;
        RECT 131.750 735.720 134.130 736.170 ;
        RECT 134.970 735.720 137.350 736.170 ;
        RECT 138.190 735.720 141.030 736.170 ;
        RECT 141.870 735.720 144.250 736.170 ;
        RECT 145.090 735.720 147.470 736.170 ;
        RECT 148.310 735.720 150.690 736.170 ;
        RECT 151.530 735.720 153.910 736.170 ;
        RECT 154.750 735.720 157.130 736.170 ;
        RECT 157.970 735.720 160.350 736.170 ;
        RECT 161.190 735.720 163.570 736.170 ;
        RECT 164.410 735.720 166.790 736.170 ;
        RECT 167.630 735.720 170.010 736.170 ;
        RECT 170.850 735.720 173.230 736.170 ;
        RECT 174.070 735.720 176.450 736.170 ;
        RECT 177.290 735.720 179.670 736.170 ;
        RECT 180.510 735.720 182.890 736.170 ;
        RECT 183.730 735.720 186.110 736.170 ;
        RECT 186.950 735.720 189.790 736.170 ;
        RECT 190.630 735.720 193.010 736.170 ;
        RECT 193.850 735.720 196.230 736.170 ;
        RECT 197.070 735.720 199.450 736.170 ;
        RECT 200.290 735.720 202.670 736.170 ;
        RECT 203.510 735.720 205.890 736.170 ;
        RECT 206.730 735.720 209.110 736.170 ;
        RECT 209.950 735.720 212.330 736.170 ;
        RECT 213.170 735.720 215.550 736.170 ;
        RECT 216.390 735.720 218.770 736.170 ;
        RECT 219.610 735.720 221.990 736.170 ;
        RECT 222.830 735.720 225.210 736.170 ;
        RECT 226.050 735.720 228.430 736.170 ;
        RECT 229.270 735.720 231.650 736.170 ;
        RECT 232.490 735.720 235.330 736.170 ;
        RECT 236.170 735.720 238.550 736.170 ;
        RECT 239.390 735.720 241.770 736.170 ;
        RECT 242.610 735.720 244.990 736.170 ;
        RECT 245.830 735.720 248.210 736.170 ;
        RECT 249.050 735.720 251.430 736.170 ;
        RECT 252.270 735.720 254.650 736.170 ;
        RECT 255.490 735.720 257.870 736.170 ;
        RECT 258.710 735.720 261.090 736.170 ;
        RECT 261.930 735.720 264.310 736.170 ;
        RECT 265.150 735.720 267.530 736.170 ;
        RECT 268.370 735.720 270.750 736.170 ;
        RECT 271.590 735.720 273.970 736.170 ;
        RECT 274.810 735.720 277.190 736.170 ;
        RECT 278.030 735.720 280.870 736.170 ;
        RECT 281.710 735.720 284.090 736.170 ;
        RECT 284.930 735.720 287.310 736.170 ;
        RECT 288.150 735.720 290.530 736.170 ;
        RECT 291.370 735.720 293.750 736.170 ;
        RECT 294.590 735.720 296.970 736.170 ;
        RECT 297.810 735.720 300.190 736.170 ;
        RECT 301.030 735.720 303.410 736.170 ;
        RECT 304.250 735.720 306.630 736.170 ;
        RECT 307.470 735.720 309.850 736.170 ;
        RECT 310.690 735.720 313.070 736.170 ;
        RECT 313.910 735.720 316.290 736.170 ;
        RECT 317.130 735.720 319.510 736.170 ;
        RECT 320.350 735.720 322.730 736.170 ;
        RECT 323.570 735.720 325.950 736.170 ;
        RECT 326.790 735.720 329.630 736.170 ;
        RECT 330.470 735.720 332.850 736.170 ;
        RECT 333.690 735.720 336.070 736.170 ;
        RECT 336.910 735.720 339.290 736.170 ;
        RECT 340.130 735.720 342.510 736.170 ;
        RECT 343.350 735.720 345.730 736.170 ;
        RECT 346.570 735.720 348.950 736.170 ;
        RECT 349.790 735.720 352.170 736.170 ;
        RECT 353.010 735.720 355.390 736.170 ;
        RECT 356.230 735.720 358.610 736.170 ;
        RECT 359.450 735.720 361.830 736.170 ;
        RECT 362.670 735.720 365.050 736.170 ;
        RECT 365.890 735.720 368.270 736.170 ;
        RECT 369.110 735.720 371.490 736.170 ;
        RECT 372.330 735.720 375.170 736.170 ;
        RECT 376.010 735.720 378.390 736.170 ;
        RECT 379.230 735.720 381.610 736.170 ;
        RECT 382.450 735.720 384.830 736.170 ;
        RECT 385.670 735.720 388.050 736.170 ;
        RECT 388.890 735.720 391.270 736.170 ;
        RECT 392.110 735.720 394.490 736.170 ;
        RECT 395.330 735.720 397.710 736.170 ;
        RECT 398.550 735.720 400.930 736.170 ;
        RECT 401.770 735.720 404.150 736.170 ;
        RECT 404.990 735.720 407.370 736.170 ;
        RECT 408.210 735.720 410.590 736.170 ;
        RECT 411.430 735.720 413.810 736.170 ;
        RECT 414.650 735.720 417.030 736.170 ;
        RECT 417.870 735.720 420.710 736.170 ;
        RECT 421.550 735.720 423.930 736.170 ;
        RECT 424.770 735.720 427.150 736.170 ;
        RECT 427.990 735.720 430.370 736.170 ;
        RECT 431.210 735.720 433.590 736.170 ;
        RECT 434.430 735.720 436.810 736.170 ;
        RECT 437.650 735.720 440.030 736.170 ;
        RECT 440.870 735.720 443.250 736.170 ;
        RECT 444.090 735.720 446.470 736.170 ;
        RECT 447.310 735.720 449.690 736.170 ;
        RECT 450.530 735.720 452.910 736.170 ;
        RECT 453.750 735.720 456.130 736.170 ;
        RECT 456.970 735.720 459.350 736.170 ;
        RECT 460.190 735.720 462.570 736.170 ;
        RECT 463.410 735.720 465.790 736.170 ;
        RECT 466.630 735.720 469.470 736.170 ;
        RECT 470.310 735.720 472.690 736.170 ;
        RECT 473.530 735.720 475.910 736.170 ;
        RECT 476.750 735.720 479.130 736.170 ;
        RECT 479.970 735.720 482.350 736.170 ;
        RECT 483.190 735.720 485.570 736.170 ;
        RECT 486.410 735.720 488.790 736.170 ;
        RECT 489.630 735.720 492.010 736.170 ;
        RECT 492.850 735.720 495.230 736.170 ;
        RECT 496.070 735.720 498.450 736.170 ;
        RECT 499.290 735.720 501.670 736.170 ;
        RECT 502.510 735.720 504.890 736.170 ;
        RECT 505.730 735.720 508.110 736.170 ;
        RECT 508.950 735.720 511.330 736.170 ;
        RECT 512.170 735.720 515.010 736.170 ;
        RECT 515.850 735.720 518.230 736.170 ;
        RECT 519.070 735.720 521.450 736.170 ;
        RECT 522.290 735.720 524.670 736.170 ;
        RECT 525.510 735.720 527.890 736.170 ;
        RECT 528.730 735.720 531.110 736.170 ;
        RECT 531.950 735.720 534.330 736.170 ;
        RECT 535.170 735.720 537.550 736.170 ;
        RECT 538.390 735.720 540.770 736.170 ;
        RECT 541.610 735.720 543.990 736.170 ;
        RECT 544.830 735.720 547.210 736.170 ;
        RECT 548.050 735.720 550.430 736.170 ;
        RECT 551.270 735.720 553.650 736.170 ;
        RECT 554.490 735.720 556.870 736.170 ;
        RECT 557.710 735.720 560.550 736.170 ;
        RECT 561.390 735.720 563.770 736.170 ;
        RECT 564.610 735.720 566.990 736.170 ;
        RECT 567.830 735.720 570.210 736.170 ;
        RECT 571.050 735.720 573.430 736.170 ;
        RECT 574.270 735.720 576.650 736.170 ;
        RECT 577.490 735.720 579.870 736.170 ;
        RECT 580.710 735.720 583.090 736.170 ;
        RECT 583.930 735.720 586.310 736.170 ;
        RECT 587.150 735.720 589.530 736.170 ;
        RECT 590.370 735.720 592.750 736.170 ;
        RECT 593.590 735.720 595.970 736.170 ;
        RECT 596.810 735.720 599.190 736.170 ;
        RECT 600.030 735.720 602.410 736.170 ;
        RECT 603.250 735.720 606.090 736.170 ;
        RECT 606.930 735.720 609.310 736.170 ;
        RECT 610.150 735.720 612.530 736.170 ;
        RECT 613.370 735.720 615.750 736.170 ;
        RECT 616.590 735.720 618.970 736.170 ;
        RECT 619.810 735.720 622.190 736.170 ;
        RECT 623.030 735.720 625.410 736.170 ;
        RECT 626.250 735.720 628.630 736.170 ;
        RECT 629.470 735.720 631.850 736.170 ;
        RECT 632.690 735.720 635.070 736.170 ;
        RECT 635.910 735.720 638.290 736.170 ;
        RECT 639.130 735.720 641.510 736.170 ;
        RECT 642.350 735.720 644.730 736.170 ;
        RECT 645.570 735.720 647.950 736.170 ;
        RECT 648.790 735.720 651.170 736.170 ;
        RECT 652.010 735.720 654.850 736.170 ;
        RECT 655.690 735.720 658.070 736.170 ;
        RECT 658.910 735.720 661.290 736.170 ;
        RECT 662.130 735.720 664.510 736.170 ;
        RECT 665.350 735.720 667.730 736.170 ;
        RECT 668.570 735.720 670.950 736.170 ;
        RECT 671.790 735.720 674.170 736.170 ;
        RECT 675.010 735.720 677.390 736.170 ;
        RECT 678.230 735.720 680.610 736.170 ;
        RECT 681.450 735.720 683.830 736.170 ;
        RECT 684.670 735.720 687.050 736.170 ;
        RECT 687.890 735.720 690.270 736.170 ;
        RECT 691.110 735.720 693.490 736.170 ;
        RECT 694.330 735.720 696.710 736.170 ;
        RECT 697.550 735.720 700.390 736.170 ;
        RECT 701.230 735.720 703.610 736.170 ;
        RECT 704.450 735.720 706.830 736.170 ;
        RECT 707.670 735.720 710.050 736.170 ;
        RECT 710.890 735.720 713.270 736.170 ;
        RECT 714.110 735.720 716.490 736.170 ;
        RECT 717.330 735.720 719.710 736.170 ;
        RECT 720.550 735.720 722.930 736.170 ;
        RECT 723.770 735.720 726.150 736.170 ;
        RECT 726.990 735.720 729.370 736.170 ;
        RECT 730.210 735.720 732.590 736.170 ;
        RECT 733.430 735.720 735.810 736.170 ;
        RECT 736.650 735.720 739.030 736.170 ;
        RECT 739.870 735.720 742.250 736.170 ;
        RECT 743.090 735.720 745.930 736.170 ;
        RECT 746.770 735.720 749.150 736.170 ;
        RECT 749.990 735.720 752.370 736.170 ;
        RECT 753.210 735.720 755.590 736.170 ;
        RECT 756.430 735.720 758.810 736.170 ;
        RECT 759.650 735.720 762.030 736.170 ;
        RECT 762.870 735.720 765.250 736.170 ;
        RECT 766.090 735.720 768.470 736.170 ;
        RECT 769.310 735.720 771.690 736.170 ;
        RECT 772.530 735.720 774.910 736.170 ;
        RECT 775.750 735.720 778.130 736.170 ;
        RECT 778.970 735.720 781.350 736.170 ;
        RECT 782.190 735.720 784.570 736.170 ;
        RECT 785.410 735.720 787.790 736.170 ;
        RECT 788.630 735.720 791.010 736.170 ;
        RECT 791.850 735.720 794.690 736.170 ;
        RECT 795.530 735.720 797.910 736.170 ;
        RECT 798.750 735.720 801.130 736.170 ;
        RECT 801.970 735.720 804.350 736.170 ;
        RECT 805.190 735.720 807.570 736.170 ;
        RECT 808.410 735.720 810.790 736.170 ;
        RECT 811.630 735.720 814.010 736.170 ;
        RECT 814.850 735.720 817.230 736.170 ;
        RECT 818.070 735.720 820.450 736.170 ;
        RECT 821.290 735.720 823.670 736.170 ;
        RECT 824.510 735.720 826.890 736.170 ;
        RECT 827.730 735.720 830.110 736.170 ;
        RECT 830.950 735.720 833.330 736.170 ;
        RECT 834.170 735.720 836.550 736.170 ;
        RECT 837.390 735.720 840.230 736.170 ;
        RECT 841.070 735.720 843.450 736.170 ;
        RECT 844.290 735.720 846.670 736.170 ;
        RECT 847.510 735.720 849.890 736.170 ;
        RECT 850.730 735.720 853.110 736.170 ;
        RECT 853.950 735.720 856.330 736.170 ;
        RECT 857.170 735.720 859.550 736.170 ;
        RECT 860.390 735.720 862.770 736.170 ;
        RECT 863.610 735.720 865.990 736.170 ;
        RECT 866.830 735.720 869.210 736.170 ;
        RECT 870.050 735.720 872.430 736.170 ;
        RECT 873.270 735.720 875.650 736.170 ;
        RECT 876.490 735.720 878.870 736.170 ;
        RECT 879.710 735.720 882.090 736.170 ;
        RECT 882.930 735.720 885.770 736.170 ;
        RECT 886.610 735.720 888.990 736.170 ;
        RECT 889.830 735.720 892.210 736.170 ;
        RECT 893.050 735.720 895.430 736.170 ;
        RECT 896.270 735.720 898.650 736.170 ;
        RECT 899.490 735.720 901.870 736.170 ;
        RECT 902.710 735.720 905.090 736.170 ;
        RECT 905.930 735.720 908.310 736.170 ;
        RECT 909.150 735.720 911.530 736.170 ;
        RECT 912.370 735.720 914.750 736.170 ;
        RECT 915.590 735.720 917.970 736.170 ;
        RECT 918.810 735.720 921.190 736.170 ;
        RECT 922.030 735.720 924.410 736.170 ;
        RECT 925.250 735.720 927.630 736.170 ;
        RECT 928.470 735.720 930.850 736.170 ;
        RECT 931.690 735.720 934.530 736.170 ;
        RECT 935.370 735.720 937.750 736.170 ;
        RECT 938.590 735.720 940.970 736.170 ;
        RECT 941.810 735.720 944.190 736.170 ;
        RECT 945.030 735.720 947.410 736.170 ;
        RECT 948.250 735.720 950.630 736.170 ;
        RECT 951.470 735.720 953.850 736.170 ;
        RECT 954.690 735.720 957.070 736.170 ;
        RECT 957.910 735.720 960.290 736.170 ;
        RECT 961.130 735.720 963.510 736.170 ;
        RECT 964.350 735.720 966.730 736.170 ;
        RECT 967.570 735.720 969.950 736.170 ;
        RECT 970.790 735.720 973.170 736.170 ;
        RECT 974.010 735.720 976.390 736.170 ;
        RECT 977.230 735.720 980.070 736.170 ;
        RECT 980.910 735.720 983.290 736.170 ;
        RECT 984.130 735.720 986.510 736.170 ;
        RECT 987.350 735.720 989.730 736.170 ;
        RECT 990.570 735.720 992.950 736.170 ;
        RECT 993.790 735.720 996.170 736.170 ;
        RECT 997.010 735.720 999.390 736.170 ;
        RECT 1000.230 735.720 1002.610 736.170 ;
        RECT 1003.450 735.720 1005.830 736.170 ;
        RECT 1006.670 735.720 1009.050 736.170 ;
        RECT 1009.890 735.720 1012.270 736.170 ;
        RECT 1013.110 735.720 1015.490 736.170 ;
        RECT 1016.330 735.720 1018.710 736.170 ;
        RECT 1019.550 735.720 1021.930 736.170 ;
        RECT 1022.770 735.720 1025.610 736.170 ;
        RECT 1026.450 735.720 1028.830 736.170 ;
        RECT 1029.670 735.720 1032.050 736.170 ;
        RECT 1032.890 735.720 1035.270 736.170 ;
        RECT 1036.110 735.720 1038.490 736.170 ;
        RECT 1039.330 735.720 1041.710 736.170 ;
        RECT 1042.550 735.720 1044.930 736.170 ;
        RECT 1045.770 735.720 1048.150 736.170 ;
        RECT 1048.990 735.720 1051.370 736.170 ;
        RECT 1052.210 735.720 1054.590 736.170 ;
        RECT 1055.430 735.720 1057.810 736.170 ;
        RECT 1058.650 735.720 1061.030 736.170 ;
        RECT 1061.870 735.720 1064.250 736.170 ;
        RECT 1065.090 735.720 1067.470 736.170 ;
        RECT 1068.310 735.720 1071.150 736.170 ;
        RECT 1071.990 735.720 1074.370 736.170 ;
        RECT 1075.210 735.720 1077.590 736.170 ;
        RECT 1078.430 735.720 1080.810 736.170 ;
        RECT 1081.650 735.720 1084.030 736.170 ;
        RECT 1084.870 735.720 1087.250 736.170 ;
        RECT 1088.090 735.720 1090.470 736.170 ;
        RECT 1091.310 735.720 1093.690 736.170 ;
        RECT 1094.530 735.720 1096.910 736.170 ;
        RECT 1097.750 735.720 1100.130 736.170 ;
        RECT 1100.970 735.720 1103.350 736.170 ;
        RECT 1104.190 735.720 1106.570 736.170 ;
        RECT 1107.410 735.720 1109.790 736.170 ;
        RECT 1110.630 735.720 1113.010 736.170 ;
        RECT 1113.850 735.720 1116.230 736.170 ;
        RECT 1117.070 735.720 1119.910 736.170 ;
        RECT 1120.750 735.720 1123.130 736.170 ;
        RECT 1123.970 735.720 1126.350 736.170 ;
        RECT 1127.190 735.720 1129.570 736.170 ;
        RECT 1130.410 735.720 1132.790 736.170 ;
        RECT 1133.630 735.720 1136.010 736.170 ;
        RECT 1136.850 735.720 1139.230 736.170 ;
        RECT 1140.070 735.720 1142.450 736.170 ;
        RECT 1143.290 735.720 1145.670 736.170 ;
        RECT 1146.510 735.720 1148.890 736.170 ;
        RECT 1149.730 735.720 1152.110 736.170 ;
        RECT 1152.950 735.720 1155.330 736.170 ;
        RECT 1156.170 735.720 1158.550 736.170 ;
        RECT 1159.390 735.720 1161.770 736.170 ;
        RECT 1162.610 735.720 1165.450 736.170 ;
        RECT 1166.290 735.720 1168.670 736.170 ;
        RECT 1169.510 735.720 1171.890 736.170 ;
        RECT 1172.730 735.720 1175.110 736.170 ;
        RECT 1175.950 735.720 1178.330 736.170 ;
        RECT 1179.170 735.720 1181.550 736.170 ;
        RECT 1182.390 735.720 1184.770 736.170 ;
        RECT 1185.610 735.720 1187.990 736.170 ;
        RECT 1188.830 735.720 1191.210 736.170 ;
        RECT 1192.050 735.720 1194.430 736.170 ;
        RECT 1195.270 735.720 1197.650 736.170 ;
        RECT 1198.490 735.720 1200.870 736.170 ;
        RECT 1201.710 735.720 1204.090 736.170 ;
        RECT 1204.930 735.720 1207.310 736.170 ;
        RECT 1208.150 735.720 1210.990 736.170 ;
        RECT 1211.830 735.720 1214.210 736.170 ;
        RECT 1215.050 735.720 1217.430 736.170 ;
        RECT 1218.270 735.720 1220.650 736.170 ;
        RECT 1221.490 735.720 1223.870 736.170 ;
        RECT 1224.710 735.720 1227.090 736.170 ;
        RECT 1227.930 735.720 1230.310 736.170 ;
        RECT 1231.150 735.720 1233.530 736.170 ;
        RECT 1234.370 735.720 1236.750 736.170 ;
        RECT 1237.590 735.720 1239.970 736.170 ;
        RECT 1240.810 735.720 1243.190 736.170 ;
        RECT 1244.030 735.720 1246.410 736.170 ;
        RECT 1247.250 735.720 1249.630 736.170 ;
        RECT 1250.470 735.720 1252.850 736.170 ;
        RECT 1253.690 735.720 1256.070 736.170 ;
        RECT 1256.910 735.720 1259.750 736.170 ;
        RECT 1260.590 735.720 1262.970 736.170 ;
        RECT 1263.810 735.720 1266.190 736.170 ;
        RECT 1267.030 735.720 1269.410 736.170 ;
        RECT 1270.250 735.720 1272.630 736.170 ;
        RECT 1273.470 735.720 1275.850 736.170 ;
        RECT 1276.690 735.720 1279.070 736.170 ;
        RECT 1279.910 735.720 1282.290 736.170 ;
        RECT 1283.130 735.720 1285.510 736.170 ;
        RECT 1286.350 735.720 1288.730 736.170 ;
        RECT 1289.570 735.720 1291.950 736.170 ;
        RECT 1292.790 735.720 1295.170 736.170 ;
        RECT 1296.010 735.720 1298.390 736.170 ;
        RECT 1299.230 735.720 1301.610 736.170 ;
        RECT 1302.450 735.720 1305.290 736.170 ;
        RECT 1306.130 735.720 1308.510 736.170 ;
        RECT 1309.350 735.720 1311.730 736.170 ;
        RECT 1312.570 735.720 1314.950 736.170 ;
        RECT 1315.790 735.720 1318.170 736.170 ;
        RECT 1319.010 735.720 1321.390 736.170 ;
        RECT 1322.230 735.720 1324.610 736.170 ;
        RECT 1325.450 735.720 1327.830 736.170 ;
        RECT 1328.670 735.720 1331.050 736.170 ;
        RECT 1331.890 735.720 1334.270 736.170 ;
        RECT 1335.110 735.720 1337.490 736.170 ;
        RECT 1338.330 735.720 1340.710 736.170 ;
        RECT 1341.550 735.720 1343.930 736.170 ;
        RECT 1344.770 735.720 1347.150 736.170 ;
        RECT 1347.990 735.720 1350.830 736.170 ;
        RECT 1351.670 735.720 1354.050 736.170 ;
        RECT 1354.890 735.720 1357.270 736.170 ;
        RECT 1358.110 735.720 1360.490 736.170 ;
        RECT 1361.330 735.720 1363.710 736.170 ;
        RECT 1364.550 735.720 1366.930 736.170 ;
        RECT 1367.770 735.720 1370.150 736.170 ;
        RECT 1370.990 735.720 1373.370 736.170 ;
        RECT 1374.210 735.720 1376.590 736.170 ;
        RECT 1377.430 735.720 1379.810 736.170 ;
        RECT 1380.650 735.720 1383.030 736.170 ;
        RECT 1383.870 735.720 1386.250 736.170 ;
        RECT 1387.090 735.720 1389.470 736.170 ;
        RECT 1390.310 735.720 1392.690 736.170 ;
        RECT 1393.530 735.720 1395.910 736.170 ;
        RECT 1396.750 735.720 1399.590 736.170 ;
        RECT 1400.430 735.720 1402.810 736.170 ;
        RECT 1403.650 735.720 1406.030 736.170 ;
        RECT 1406.870 735.720 1409.250 736.170 ;
        RECT 1410.090 735.720 1412.470 736.170 ;
        RECT 1413.310 735.720 1415.690 736.170 ;
        RECT 1416.530 735.720 1418.910 736.170 ;
        RECT 1419.750 735.720 1422.130 736.170 ;
        RECT 1422.970 735.720 1425.350 736.170 ;
        RECT 1426.190 735.720 1428.570 736.170 ;
        RECT 1429.410 735.720 1431.790 736.170 ;
        RECT 1432.630 735.720 1435.010 736.170 ;
        RECT 1435.850 735.720 1438.230 736.170 ;
        RECT 1439.070 735.720 1441.450 736.170 ;
        RECT 1442.290 735.720 1445.130 736.170 ;
        RECT 1445.970 735.720 1448.350 736.170 ;
        RECT 1449.190 735.720 1451.570 736.170 ;
        RECT 1452.410 735.720 1454.790 736.170 ;
        RECT 1455.630 735.720 1458.010 736.170 ;
        RECT 1458.850 735.720 1461.230 736.170 ;
        RECT 1462.070 735.720 1464.450 736.170 ;
        RECT 1465.290 735.720 1467.670 736.170 ;
        RECT 1468.510 735.720 1470.890 736.170 ;
        RECT 1471.730 735.720 1474.110 736.170 ;
        RECT 1474.950 735.720 1477.330 736.170 ;
        RECT 1478.170 735.720 1480.550 736.170 ;
        RECT 1481.390 735.720 1483.770 736.170 ;
        RECT 1484.610 735.720 1486.990 736.170 ;
        RECT 1487.830 735.720 1490.670 736.170 ;
        RECT 1491.510 735.720 1493.890 736.170 ;
        RECT 1494.730 735.720 1497.110 736.170 ;
        RECT 1497.950 735.720 1500.330 736.170 ;
        RECT 1501.170 735.720 1503.550 736.170 ;
        RECT 1504.390 735.720 1506.770 736.170 ;
        RECT 1507.610 735.720 1509.990 736.170 ;
        RECT 1510.830 735.720 1513.210 736.170 ;
        RECT 1514.050 735.720 1516.430 736.170 ;
        RECT 1517.270 735.720 1519.650 736.170 ;
        RECT 1520.490 735.720 1522.870 736.170 ;
        RECT 1523.710 735.720 1526.090 736.170 ;
        RECT 1526.930 735.720 1529.310 736.170 ;
        RECT 1530.150 735.720 1532.530 736.170 ;
        RECT 1533.370 735.720 1536.210 736.170 ;
        RECT 1537.050 735.720 1539.430 736.170 ;
        RECT 1540.270 735.720 1542.650 736.170 ;
        RECT 1543.490 735.720 1545.870 736.170 ;
        RECT 1546.710 735.720 1549.090 736.170 ;
        RECT 1549.930 735.720 1552.310 736.170 ;
        RECT 1553.150 735.720 1555.530 736.170 ;
        RECT 1556.370 735.720 1558.750 736.170 ;
        RECT 1559.590 735.720 1561.970 736.170 ;
        RECT 1562.810 735.720 1565.190 736.170 ;
        RECT 1566.030 735.720 1568.410 736.170 ;
        RECT 1569.250 735.720 1571.630 736.170 ;
        RECT 1572.470 735.720 1574.850 736.170 ;
        RECT 1575.690 735.720 1578.070 736.170 ;
        RECT 1578.910 735.720 1581.290 736.170 ;
        RECT 1582.130 735.720 1584.970 736.170 ;
        RECT 1585.810 735.720 1588.190 736.170 ;
        RECT 1589.030 735.720 1591.410 736.170 ;
        RECT 1592.250 735.720 1594.630 736.170 ;
        RECT 1595.470 735.720 1597.850 736.170 ;
        RECT 1598.690 735.720 1601.070 736.170 ;
        RECT 1601.910 735.720 1604.290 736.170 ;
        RECT 1605.130 735.720 1607.510 736.170 ;
        RECT 1608.350 735.720 1610.730 736.170 ;
        RECT 1611.570 735.720 1613.950 736.170 ;
        RECT 1614.790 735.720 1617.170 736.170 ;
        RECT 1618.010 735.720 1620.390 736.170 ;
        RECT 1621.230 735.720 1623.610 736.170 ;
        RECT 1624.450 735.720 1626.830 736.170 ;
        RECT 1627.670 735.720 1630.510 736.170 ;
        RECT 1631.350 735.720 1633.730 736.170 ;
        RECT 1634.570 735.720 1636.950 736.170 ;
        RECT 1637.790 735.720 1640.170 736.170 ;
        RECT 1641.010 735.720 1643.390 736.170 ;
        RECT 1644.230 735.720 1646.610 736.170 ;
        RECT 1647.450 735.720 1649.830 736.170 ;
        RECT 1650.670 735.720 1653.050 736.170 ;
        RECT 1653.890 735.720 1656.270 736.170 ;
        RECT 1657.110 735.720 1659.490 736.170 ;
        RECT 1660.330 735.720 1662.710 736.170 ;
        RECT 1663.550 735.720 1665.930 736.170 ;
        RECT 1666.770 735.720 1669.150 736.170 ;
        RECT 1669.990 735.720 1672.370 736.170 ;
        RECT 1673.210 735.720 1676.050 736.170 ;
        RECT 1676.890 735.720 1679.270 736.170 ;
        RECT 1680.110 735.720 1682.490 736.170 ;
        RECT 1683.330 735.720 1685.710 736.170 ;
        RECT 1686.550 735.720 1688.930 736.170 ;
        RECT 1689.770 735.720 1692.150 736.170 ;
        RECT 1692.990 735.720 1695.370 736.170 ;
        RECT 1696.210 735.720 1698.590 736.170 ;
        RECT 1699.430 735.720 1701.810 736.170 ;
        RECT 1702.650 735.720 1705.030 736.170 ;
        RECT 1705.870 735.720 1708.250 736.170 ;
        RECT 1709.090 735.720 1711.470 736.170 ;
        RECT 1712.310 735.720 1714.690 736.170 ;
        RECT 1715.530 735.720 1717.910 736.170 ;
        RECT 1718.750 735.720 1721.130 736.170 ;
        RECT 1721.970 735.720 1724.810 736.170 ;
        RECT 1725.650 735.720 1728.030 736.170 ;
        RECT 1728.870 735.720 1731.250 736.170 ;
        RECT 1732.090 735.720 1734.470 736.170 ;
        RECT 1735.310 735.720 1737.690 736.170 ;
        RECT 1738.530 735.720 1740.910 736.170 ;
        RECT 1741.750 735.720 1744.130 736.170 ;
        RECT 1744.970 735.720 1747.350 736.170 ;
        RECT 1748.190 735.720 1750.570 736.170 ;
        RECT 1751.410 735.720 1753.790 736.170 ;
        RECT 1754.630 735.720 1757.010 736.170 ;
        RECT 1757.850 735.720 1760.230 736.170 ;
        RECT 1761.070 735.720 1763.450 736.170 ;
        RECT 1764.290 735.720 1766.670 736.170 ;
        RECT 1767.510 735.720 1770.350 736.170 ;
        RECT 1771.190 735.720 1773.570 736.170 ;
        RECT 1774.410 735.720 1776.790 736.170 ;
        RECT 1777.630 735.720 1780.010 736.170 ;
        RECT 1780.850 735.720 1783.230 736.170 ;
        RECT 1784.070 735.720 1786.450 736.170 ;
        RECT 1787.290 735.720 1789.670 736.170 ;
        RECT 1790.510 735.720 1792.890 736.170 ;
        RECT 1793.730 735.720 1796.110 736.170 ;
        RECT 1796.950 735.720 1799.330 736.170 ;
        RECT 1800.170 735.720 1802.550 736.170 ;
        RECT 1803.390 735.720 1805.770 736.170 ;
        RECT 1806.610 735.720 1808.990 736.170 ;
        RECT 1809.830 735.720 1812.210 736.170 ;
        RECT 1813.050 735.720 1815.890 736.170 ;
        RECT 1816.730 735.720 1819.110 736.170 ;
        RECT 1819.950 735.720 1822.330 736.170 ;
        RECT 1823.170 735.720 1825.550 736.170 ;
        RECT 1826.390 735.720 1828.770 736.170 ;
        RECT 1829.610 735.720 1831.990 736.170 ;
        RECT 1832.830 735.720 1835.210 736.170 ;
        RECT 1836.050 735.720 1838.430 736.170 ;
        RECT 1839.270 735.720 1841.650 736.170 ;
        RECT 1842.490 735.720 1844.870 736.170 ;
        RECT 1845.710 735.720 1848.090 736.170 ;
        RECT 1848.930 735.720 1851.310 736.170 ;
        RECT 1852.150 735.720 1854.530 736.170 ;
        RECT 1855.370 735.720 1857.750 736.170 ;
        RECT 1858.590 735.720 1860.970 736.170 ;
        RECT 1861.810 735.720 1864.650 736.170 ;
        RECT 1865.490 735.720 1867.870 736.170 ;
        RECT 1868.710 735.720 1871.090 736.170 ;
        RECT 1871.930 735.720 1874.310 736.170 ;
        RECT 1875.150 735.720 1877.530 736.170 ;
        RECT 1878.370 735.720 1880.750 736.170 ;
        RECT 1881.590 735.720 1883.970 736.170 ;
        RECT 1884.810 735.720 1887.190 736.170 ;
        RECT 1888.030 735.720 1890.410 736.170 ;
        RECT 1891.250 735.720 1893.630 736.170 ;
        RECT 1894.470 735.720 1896.850 736.170 ;
        RECT 1897.690 735.720 1900.070 736.170 ;
        RECT 1900.910 735.720 1903.290 736.170 ;
        RECT 1904.130 735.720 1906.510 736.170 ;
        RECT 1907.350 735.720 1910.190 736.170 ;
        RECT 1911.030 735.720 1913.410 736.170 ;
        RECT 1914.250 735.720 1916.630 736.170 ;
        RECT 1917.470 735.720 1919.850 736.170 ;
        RECT 1920.690 735.720 1923.070 736.170 ;
        RECT 1923.910 735.720 1926.290 736.170 ;
        RECT 1927.130 735.720 1929.510 736.170 ;
        RECT 1930.350 735.720 1932.730 736.170 ;
        RECT 1933.570 735.720 1935.950 736.170 ;
        RECT 1936.790 735.720 1939.170 736.170 ;
        RECT 1940.010 735.720 1942.390 736.170 ;
        RECT 1943.230 735.720 1945.610 736.170 ;
        RECT 1946.450 735.720 1948.830 736.170 ;
        RECT 1949.670 735.720 1952.050 736.170 ;
        RECT 1952.890 735.720 1955.730 736.170 ;
        RECT 1956.570 735.720 1958.950 736.170 ;
        RECT 1959.790 735.720 1962.170 736.170 ;
        RECT 1963.010 735.720 1965.390 736.170 ;
        RECT 1966.230 735.720 1968.610 736.170 ;
        RECT 1969.450 735.720 1971.830 736.170 ;
        RECT 1972.670 735.720 1975.050 736.170 ;
        RECT 1975.890 735.720 1978.270 736.170 ;
        RECT 1979.110 735.720 1981.490 736.170 ;
        RECT 1982.330 735.720 1984.710 736.170 ;
        RECT 1985.550 735.720 1987.930 736.170 ;
        RECT 1988.770 735.720 1991.150 736.170 ;
        RECT 1991.990 735.720 1994.370 736.170 ;
        RECT 1995.210 735.720 1997.590 736.170 ;
        RECT 1.480 4.280 1998.140 735.720 ;
        RECT 1.480 3.670 8.090 4.280 ;
        RECT 8.930 3.670 24.650 4.280 ;
        RECT 25.490 3.670 41.670 4.280 ;
        RECT 42.510 3.670 58.230 4.280 ;
        RECT 59.070 3.670 75.250 4.280 ;
        RECT 76.090 3.670 91.810 4.280 ;
        RECT 92.650 3.670 108.830 4.280 ;
        RECT 109.670 3.670 125.390 4.280 ;
        RECT 126.230 3.670 142.410 4.280 ;
        RECT 143.250 3.670 158.970 4.280 ;
        RECT 159.810 3.670 175.990 4.280 ;
        RECT 176.830 3.670 192.550 4.280 ;
        RECT 193.390 3.670 209.570 4.280 ;
        RECT 210.410 3.670 226.130 4.280 ;
        RECT 226.970 3.670 243.150 4.280 ;
        RECT 243.990 3.670 260.170 4.280 ;
        RECT 261.010 3.670 276.730 4.280 ;
        RECT 277.570 3.670 293.750 4.280 ;
        RECT 294.590 3.670 310.310 4.280 ;
        RECT 311.150 3.670 327.330 4.280 ;
        RECT 328.170 3.670 343.890 4.280 ;
        RECT 344.730 3.670 360.910 4.280 ;
        RECT 361.750 3.670 377.470 4.280 ;
        RECT 378.310 3.670 394.490 4.280 ;
        RECT 395.330 3.670 411.050 4.280 ;
        RECT 411.890 3.670 428.070 4.280 ;
        RECT 428.910 3.670 444.630 4.280 ;
        RECT 445.470 3.670 461.650 4.280 ;
        RECT 462.490 3.670 478.670 4.280 ;
        RECT 479.510 3.670 495.230 4.280 ;
        RECT 496.070 3.670 512.250 4.280 ;
        RECT 513.090 3.670 528.810 4.280 ;
        RECT 529.650 3.670 545.830 4.280 ;
        RECT 546.670 3.670 562.390 4.280 ;
        RECT 563.230 3.670 579.410 4.280 ;
        RECT 580.250 3.670 595.970 4.280 ;
        RECT 596.810 3.670 612.990 4.280 ;
        RECT 613.830 3.670 629.550 4.280 ;
        RECT 630.390 3.670 646.570 4.280 ;
        RECT 647.410 3.670 663.130 4.280 ;
        RECT 663.970 3.670 680.150 4.280 ;
        RECT 680.990 3.670 697.170 4.280 ;
        RECT 698.010 3.670 713.730 4.280 ;
        RECT 714.570 3.670 730.750 4.280 ;
        RECT 731.590 3.670 747.310 4.280 ;
        RECT 748.150 3.670 764.330 4.280 ;
        RECT 765.170 3.670 780.890 4.280 ;
        RECT 781.730 3.670 797.910 4.280 ;
        RECT 798.750 3.670 814.470 4.280 ;
        RECT 815.310 3.670 831.490 4.280 ;
        RECT 832.330 3.670 848.050 4.280 ;
        RECT 848.890 3.670 865.070 4.280 ;
        RECT 865.910 3.670 881.630 4.280 ;
        RECT 882.470 3.670 898.650 4.280 ;
        RECT 899.490 3.670 915.670 4.280 ;
        RECT 916.510 3.670 932.230 4.280 ;
        RECT 933.070 3.670 949.250 4.280 ;
        RECT 950.090 3.670 965.810 4.280 ;
        RECT 966.650 3.670 982.830 4.280 ;
        RECT 983.670 3.670 999.390 4.280 ;
        RECT 1000.230 3.670 1016.410 4.280 ;
        RECT 1017.250 3.670 1032.970 4.280 ;
        RECT 1033.810 3.670 1049.990 4.280 ;
        RECT 1050.830 3.670 1066.550 4.280 ;
        RECT 1067.390 3.670 1083.570 4.280 ;
        RECT 1084.410 3.670 1100.130 4.280 ;
        RECT 1100.970 3.670 1117.150 4.280 ;
        RECT 1117.990 3.670 1134.170 4.280 ;
        RECT 1135.010 3.670 1150.730 4.280 ;
        RECT 1151.570 3.670 1167.750 4.280 ;
        RECT 1168.590 3.670 1184.310 4.280 ;
        RECT 1185.150 3.670 1201.330 4.280 ;
        RECT 1202.170 3.670 1217.890 4.280 ;
        RECT 1218.730 3.670 1234.910 4.280 ;
        RECT 1235.750 3.670 1251.470 4.280 ;
        RECT 1252.310 3.670 1268.490 4.280 ;
        RECT 1269.330 3.670 1285.050 4.280 ;
        RECT 1285.890 3.670 1302.070 4.280 ;
        RECT 1302.910 3.670 1318.630 4.280 ;
        RECT 1319.470 3.670 1335.650 4.280 ;
        RECT 1336.490 3.670 1352.670 4.280 ;
        RECT 1353.510 3.670 1369.230 4.280 ;
        RECT 1370.070 3.670 1386.250 4.280 ;
        RECT 1387.090 3.670 1402.810 4.280 ;
        RECT 1403.650 3.670 1419.830 4.280 ;
        RECT 1420.670 3.670 1436.390 4.280 ;
        RECT 1437.230 3.670 1453.410 4.280 ;
        RECT 1454.250 3.670 1469.970 4.280 ;
        RECT 1470.810 3.670 1486.990 4.280 ;
        RECT 1487.830 3.670 1503.550 4.280 ;
        RECT 1504.390 3.670 1520.570 4.280 ;
        RECT 1521.410 3.670 1537.130 4.280 ;
        RECT 1537.970 3.670 1554.150 4.280 ;
        RECT 1554.990 3.670 1571.170 4.280 ;
        RECT 1572.010 3.670 1587.730 4.280 ;
        RECT 1588.570 3.670 1604.750 4.280 ;
        RECT 1605.590 3.670 1621.310 4.280 ;
        RECT 1622.150 3.670 1638.330 4.280 ;
        RECT 1639.170 3.670 1654.890 4.280 ;
        RECT 1655.730 3.670 1671.910 4.280 ;
        RECT 1672.750 3.670 1688.470 4.280 ;
        RECT 1689.310 3.670 1705.490 4.280 ;
        RECT 1706.330 3.670 1722.050 4.280 ;
        RECT 1722.890 3.670 1739.070 4.280 ;
        RECT 1739.910 3.670 1755.630 4.280 ;
        RECT 1756.470 3.670 1772.650 4.280 ;
        RECT 1773.490 3.670 1789.670 4.280 ;
        RECT 1790.510 3.670 1806.230 4.280 ;
        RECT 1807.070 3.670 1823.250 4.280 ;
        RECT 1824.090 3.670 1839.810 4.280 ;
        RECT 1840.650 3.670 1856.830 4.280 ;
        RECT 1857.670 3.670 1873.390 4.280 ;
        RECT 1874.230 3.670 1890.410 4.280 ;
        RECT 1891.250 3.670 1906.970 4.280 ;
        RECT 1907.810 3.670 1923.990 4.280 ;
        RECT 1924.830 3.670 1940.550 4.280 ;
        RECT 1941.390 3.670 1957.570 4.280 ;
        RECT 1958.410 3.670 1974.130 4.280 ;
        RECT 1974.970 3.670 1991.150 4.280 ;
        RECT 1991.990 3.670 1998.140 4.280 ;
      LAYER met3 ;
        RECT 4.400 732.680 1996.000 733.545 ;
        RECT 4.000 723.200 1996.000 732.680 ;
        RECT 4.000 721.840 1995.600 723.200 ;
        RECT 4.400 721.800 1995.600 721.840 ;
        RECT 4.400 720.440 1996.000 721.800 ;
        RECT 4.000 709.600 1996.000 720.440 ;
        RECT 4.400 708.200 1996.000 709.600 ;
        RECT 4.000 697.360 1996.000 708.200 ;
        RECT 4.400 695.960 1996.000 697.360 ;
        RECT 4.000 689.880 1996.000 695.960 ;
        RECT 4.000 688.480 1995.600 689.880 ;
        RECT 4.000 685.120 1996.000 688.480 ;
        RECT 4.400 683.720 1996.000 685.120 ;
        RECT 4.000 672.880 1996.000 683.720 ;
        RECT 4.400 671.480 1996.000 672.880 ;
        RECT 4.000 661.320 1996.000 671.480 ;
        RECT 4.400 659.920 1996.000 661.320 ;
        RECT 4.000 655.880 1996.000 659.920 ;
        RECT 4.000 654.480 1995.600 655.880 ;
        RECT 4.000 649.080 1996.000 654.480 ;
        RECT 4.400 647.680 1996.000 649.080 ;
        RECT 4.000 636.840 1996.000 647.680 ;
        RECT 4.400 635.440 1996.000 636.840 ;
        RECT 4.000 624.600 1996.000 635.440 ;
        RECT 4.400 623.200 1996.000 624.600 ;
        RECT 4.000 622.560 1996.000 623.200 ;
        RECT 4.000 621.160 1995.600 622.560 ;
        RECT 4.000 612.360 1996.000 621.160 ;
        RECT 4.400 610.960 1996.000 612.360 ;
        RECT 4.000 600.120 1996.000 610.960 ;
        RECT 4.400 598.720 1996.000 600.120 ;
        RECT 4.000 588.560 1996.000 598.720 ;
        RECT 4.400 587.160 1995.600 588.560 ;
        RECT 4.000 576.320 1996.000 587.160 ;
        RECT 4.400 574.920 1996.000 576.320 ;
        RECT 4.000 564.080 1996.000 574.920 ;
        RECT 4.400 562.680 1996.000 564.080 ;
        RECT 4.000 555.240 1996.000 562.680 ;
        RECT 4.000 553.840 1995.600 555.240 ;
        RECT 4.000 551.840 1996.000 553.840 ;
        RECT 4.400 550.440 1996.000 551.840 ;
        RECT 4.000 539.600 1996.000 550.440 ;
        RECT 4.400 538.200 1996.000 539.600 ;
        RECT 4.000 527.360 1996.000 538.200 ;
        RECT 4.400 525.960 1996.000 527.360 ;
        RECT 4.000 521.240 1996.000 525.960 ;
        RECT 4.000 519.840 1995.600 521.240 ;
        RECT 4.000 515.800 1996.000 519.840 ;
        RECT 4.400 514.400 1996.000 515.800 ;
        RECT 4.000 503.560 1996.000 514.400 ;
        RECT 4.400 502.160 1996.000 503.560 ;
        RECT 4.000 491.320 1996.000 502.160 ;
        RECT 4.400 489.920 1996.000 491.320 ;
        RECT 4.000 487.920 1996.000 489.920 ;
        RECT 4.000 486.520 1995.600 487.920 ;
        RECT 4.000 479.080 1996.000 486.520 ;
        RECT 4.400 477.680 1996.000 479.080 ;
        RECT 4.000 466.840 1996.000 477.680 ;
        RECT 4.400 465.440 1996.000 466.840 ;
        RECT 4.000 454.600 1996.000 465.440 ;
        RECT 4.400 453.920 1996.000 454.600 ;
        RECT 4.400 453.200 1995.600 453.920 ;
        RECT 4.000 452.520 1995.600 453.200 ;
        RECT 4.000 443.040 1996.000 452.520 ;
        RECT 4.400 441.640 1996.000 443.040 ;
        RECT 4.000 430.800 1996.000 441.640 ;
        RECT 4.400 429.400 1996.000 430.800 ;
        RECT 4.000 420.600 1996.000 429.400 ;
        RECT 4.000 419.200 1995.600 420.600 ;
        RECT 4.000 418.560 1996.000 419.200 ;
        RECT 4.400 417.160 1996.000 418.560 ;
        RECT 4.000 406.320 1996.000 417.160 ;
        RECT 4.400 404.920 1996.000 406.320 ;
        RECT 4.000 394.080 1996.000 404.920 ;
        RECT 4.400 392.680 1996.000 394.080 ;
        RECT 4.000 387.280 1996.000 392.680 ;
        RECT 4.000 385.880 1995.600 387.280 ;
        RECT 4.000 381.840 1996.000 385.880 ;
        RECT 4.400 380.440 1996.000 381.840 ;
        RECT 4.000 370.280 1996.000 380.440 ;
        RECT 4.400 368.880 1996.000 370.280 ;
        RECT 4.000 358.040 1996.000 368.880 ;
        RECT 4.400 356.640 1996.000 358.040 ;
        RECT 4.000 353.280 1996.000 356.640 ;
        RECT 4.000 351.880 1995.600 353.280 ;
        RECT 4.000 345.800 1996.000 351.880 ;
        RECT 4.400 344.400 1996.000 345.800 ;
        RECT 4.000 333.560 1996.000 344.400 ;
        RECT 4.400 332.160 1996.000 333.560 ;
        RECT 4.000 321.320 1996.000 332.160 ;
        RECT 4.400 319.960 1996.000 321.320 ;
        RECT 4.400 319.920 1995.600 319.960 ;
        RECT 4.000 318.560 1995.600 319.920 ;
        RECT 4.000 309.080 1996.000 318.560 ;
        RECT 4.400 307.680 1996.000 309.080 ;
        RECT 4.000 297.520 1996.000 307.680 ;
        RECT 4.400 296.120 1996.000 297.520 ;
        RECT 4.000 285.960 1996.000 296.120 ;
        RECT 4.000 285.280 1995.600 285.960 ;
        RECT 4.400 284.560 1995.600 285.280 ;
        RECT 4.400 283.880 1996.000 284.560 ;
        RECT 4.000 273.040 1996.000 283.880 ;
        RECT 4.400 271.640 1996.000 273.040 ;
        RECT 4.000 260.800 1996.000 271.640 ;
        RECT 4.400 259.400 1996.000 260.800 ;
        RECT 4.000 252.640 1996.000 259.400 ;
        RECT 4.000 251.240 1995.600 252.640 ;
        RECT 4.000 248.560 1996.000 251.240 ;
        RECT 4.400 247.160 1996.000 248.560 ;
        RECT 4.000 236.320 1996.000 247.160 ;
        RECT 4.400 234.920 1996.000 236.320 ;
        RECT 4.000 224.760 1996.000 234.920 ;
        RECT 4.400 223.360 1996.000 224.760 ;
        RECT 4.000 218.640 1996.000 223.360 ;
        RECT 4.000 217.240 1995.600 218.640 ;
        RECT 4.000 212.520 1996.000 217.240 ;
        RECT 4.400 211.120 1996.000 212.520 ;
        RECT 4.000 200.280 1996.000 211.120 ;
        RECT 4.400 198.880 1996.000 200.280 ;
        RECT 4.000 188.040 1996.000 198.880 ;
        RECT 4.400 186.640 1996.000 188.040 ;
        RECT 4.000 185.320 1996.000 186.640 ;
        RECT 4.000 183.920 1995.600 185.320 ;
        RECT 4.000 175.800 1996.000 183.920 ;
        RECT 4.400 174.400 1996.000 175.800 ;
        RECT 4.000 163.560 1996.000 174.400 ;
        RECT 4.400 162.160 1996.000 163.560 ;
        RECT 4.000 152.000 1996.000 162.160 ;
        RECT 4.400 151.320 1996.000 152.000 ;
        RECT 4.400 150.600 1995.600 151.320 ;
        RECT 4.000 149.920 1995.600 150.600 ;
        RECT 4.000 139.760 1996.000 149.920 ;
        RECT 4.400 138.360 1996.000 139.760 ;
        RECT 4.000 127.520 1996.000 138.360 ;
        RECT 4.400 126.120 1996.000 127.520 ;
        RECT 4.000 118.000 1996.000 126.120 ;
        RECT 4.000 116.600 1995.600 118.000 ;
        RECT 4.000 115.280 1996.000 116.600 ;
        RECT 4.400 113.880 1996.000 115.280 ;
        RECT 4.000 103.040 1996.000 113.880 ;
        RECT 4.400 101.640 1996.000 103.040 ;
        RECT 4.000 90.800 1996.000 101.640 ;
        RECT 4.400 89.400 1996.000 90.800 ;
        RECT 4.000 84.000 1996.000 89.400 ;
        RECT 4.000 82.600 1995.600 84.000 ;
        RECT 4.000 79.240 1996.000 82.600 ;
        RECT 4.400 77.840 1996.000 79.240 ;
        RECT 4.000 67.000 1996.000 77.840 ;
        RECT 4.400 65.600 1996.000 67.000 ;
        RECT 4.000 54.760 1996.000 65.600 ;
        RECT 4.400 53.360 1996.000 54.760 ;
        RECT 4.000 50.680 1996.000 53.360 ;
        RECT 4.000 49.280 1995.600 50.680 ;
        RECT 4.000 42.520 1996.000 49.280 ;
        RECT 4.400 41.120 1996.000 42.520 ;
        RECT 4.000 30.280 1996.000 41.120 ;
        RECT 4.400 28.880 1996.000 30.280 ;
        RECT 4.000 18.040 1996.000 28.880 ;
        RECT 4.400 17.360 1996.000 18.040 ;
        RECT 4.400 16.640 1995.600 17.360 ;
        RECT 4.000 15.960 1995.600 16.640 ;
        RECT 4.000 6.480 1996.000 15.960 ;
        RECT 4.400 5.615 1996.000 6.480 ;
      LAYER met4 ;
        RECT 18.270 11.735 25.240 723.345 ;
        RECT 27.640 11.735 50.240 723.345 ;
        RECT 52.640 11.735 75.240 723.345 ;
        RECT 77.640 536.900 100.240 723.345 ;
        RECT 102.640 536.900 125.240 723.345 ;
        RECT 127.640 536.900 150.240 723.345 ;
        RECT 152.640 536.900 175.240 723.345 ;
        RECT 177.640 536.900 200.240 723.345 ;
        RECT 202.640 536.900 225.240 723.345 ;
        RECT 227.640 536.900 250.240 723.345 ;
        RECT 252.640 536.900 275.240 723.345 ;
        RECT 277.640 536.900 300.240 723.345 ;
        RECT 302.640 536.900 325.240 723.345 ;
        RECT 327.640 536.900 350.240 723.345 ;
        RECT 352.640 536.900 375.240 723.345 ;
        RECT 377.640 536.900 400.240 723.345 ;
        RECT 402.640 536.900 425.240 723.345 ;
        RECT 427.640 536.900 450.240 723.345 ;
        RECT 452.640 536.900 475.240 723.345 ;
        RECT 477.640 536.900 500.240 723.345 ;
        RECT 502.640 536.900 525.240 723.345 ;
        RECT 527.640 536.900 550.240 723.345 ;
        RECT 552.640 536.900 575.240 723.345 ;
        RECT 577.640 536.900 600.240 723.345 ;
        RECT 602.640 536.900 625.240 723.345 ;
        RECT 627.640 536.900 650.240 723.345 ;
        RECT 652.640 536.900 675.240 723.345 ;
        RECT 677.640 536.900 700.240 723.345 ;
        RECT 702.640 536.900 725.240 723.345 ;
        RECT 727.640 536.900 750.240 723.345 ;
        RECT 752.640 536.900 775.240 723.345 ;
        RECT 777.640 536.900 800.240 723.345 ;
        RECT 77.640 101.640 800.240 536.900 ;
        RECT 77.640 11.735 100.240 101.640 ;
        RECT 102.640 11.735 125.240 101.640 ;
        RECT 127.640 11.735 150.240 101.640 ;
        RECT 152.640 11.735 175.240 101.640 ;
        RECT 177.640 11.735 200.240 101.640 ;
        RECT 202.640 11.735 225.240 101.640 ;
        RECT 227.640 11.735 250.240 101.640 ;
        RECT 252.640 11.735 275.240 101.640 ;
        RECT 277.640 11.735 300.240 101.640 ;
        RECT 302.640 11.735 325.240 101.640 ;
        RECT 327.640 11.735 350.240 101.640 ;
        RECT 352.640 11.735 375.240 101.640 ;
        RECT 377.640 11.735 400.240 101.640 ;
        RECT 402.640 11.735 425.240 101.640 ;
        RECT 427.640 11.735 450.240 101.640 ;
        RECT 452.640 11.735 475.240 101.640 ;
        RECT 477.640 11.735 500.240 101.640 ;
        RECT 502.640 11.735 525.240 101.640 ;
        RECT 527.640 11.735 550.240 101.640 ;
        RECT 552.640 11.735 575.240 101.640 ;
        RECT 577.640 11.735 600.240 101.640 ;
        RECT 602.640 11.735 625.240 101.640 ;
        RECT 627.640 11.735 650.240 101.640 ;
        RECT 652.640 11.735 675.240 101.640 ;
        RECT 677.640 11.735 700.240 101.640 ;
        RECT 702.640 11.735 725.240 101.640 ;
        RECT 727.640 11.735 750.240 101.640 ;
        RECT 752.640 11.735 775.240 101.640 ;
        RECT 777.640 11.735 800.240 101.640 ;
        RECT 802.640 11.735 825.240 723.345 ;
        RECT 827.640 11.735 850.240 723.345 ;
        RECT 852.640 11.735 875.240 723.345 ;
        RECT 877.640 11.735 900.240 723.345 ;
        RECT 902.640 11.735 925.240 723.345 ;
        RECT 927.640 11.735 950.240 723.345 ;
        RECT 952.640 11.735 975.240 723.345 ;
        RECT 977.640 11.735 1000.240 723.345 ;
        RECT 1002.640 11.735 1025.240 723.345 ;
        RECT 1027.640 11.735 1050.240 723.345 ;
        RECT 1052.640 11.735 1075.240 723.345 ;
        RECT 1077.640 11.735 1100.240 723.345 ;
        RECT 1102.640 11.735 1125.240 723.345 ;
        RECT 1127.640 11.735 1150.240 723.345 ;
        RECT 1152.640 11.735 1175.240 723.345 ;
        RECT 1177.640 11.735 1200.240 723.345 ;
        RECT 1202.640 11.735 1225.240 723.345 ;
        RECT 1227.640 11.735 1250.240 723.345 ;
        RECT 1252.640 11.735 1275.240 723.345 ;
        RECT 1277.640 11.735 1300.240 723.345 ;
        RECT 1302.640 11.735 1325.240 723.345 ;
        RECT 1327.640 11.735 1350.240 723.345 ;
        RECT 1352.640 11.735 1375.240 723.345 ;
        RECT 1377.640 11.735 1400.240 723.345 ;
        RECT 1402.640 11.735 1425.240 723.345 ;
        RECT 1427.640 11.735 1450.240 723.345 ;
        RECT 1452.640 11.735 1475.240 723.345 ;
        RECT 1477.640 11.735 1500.240 723.345 ;
        RECT 1502.640 11.735 1525.240 723.345 ;
        RECT 1527.640 11.735 1550.240 723.345 ;
        RECT 1552.640 11.735 1575.240 723.345 ;
        RECT 1577.640 11.735 1600.240 723.345 ;
        RECT 1602.640 11.735 1625.240 723.345 ;
        RECT 1627.640 11.735 1650.240 723.345 ;
        RECT 1652.640 11.735 1675.240 723.345 ;
        RECT 1677.640 11.735 1700.240 723.345 ;
        RECT 1702.640 11.735 1725.240 723.345 ;
        RECT 1727.640 11.735 1750.240 723.345 ;
        RECT 1752.640 11.735 1775.240 723.345 ;
        RECT 1777.640 11.735 1780.825 723.345 ;
      LAYER met5 ;
        RECT 18.060 679.690 1362.860 716.500 ;
        RECT 18.060 614.690 1362.860 674.890 ;
        RECT 18.060 549.690 1362.860 609.890 ;
        RECT 18.060 484.690 1362.860 544.890 ;
        RECT 18.060 419.690 1362.860 479.890 ;
        RECT 18.060 354.690 1362.860 414.890 ;
        RECT 18.060 289.690 1362.860 349.890 ;
        RECT 18.060 224.690 1362.860 284.890 ;
        RECT 18.060 159.690 1362.860 219.890 ;
        RECT 18.060 109.700 1362.860 154.890 ;
  END
END mgmt_core
END LIBRARY

