magic
tech sky130A
magscale 1 2
timestamp 1638138710
<< locali >>
rect 173081 157267 173115 157301
rect 172931 157233 173115 157267
rect 173449 156587 173483 157233
rect 173725 156587 173759 157165
rect 175933 156587 175967 157029
rect 182005 156451 182039 157301
rect 185535 157165 185627 157199
rect 185593 157063 185627 157165
rect 185501 156315 185535 157029
rect 185685 156383 185719 157301
rect 185777 156315 185811 157233
rect 185593 156281 185811 156315
rect 185409 156247 185443 156281
rect 185593 156247 185627 156281
rect 185409 156213 185627 156247
rect 195161 156247 195195 156485
rect 204913 156451 204947 156689
rect 195253 156247 195287 156349
rect 195345 156179 195379 156349
rect 194919 156145 195379 156179
rect 205005 156179 205039 156485
rect 213745 156451 213779 156757
rect 113281 155839 113315 156077
rect 118065 155635 118099 155805
rect 117973 155295 118007 155601
rect 117881 154751 117915 155261
rect 124781 155091 124815 155193
rect 127541 155091 127575 155805
rect 127449 153867 127483 155057
rect 127633 154683 127667 155805
rect 133889 155363 133923 155465
rect 137109 155431 137143 155669
rect 137235 155329 137511 155363
rect 128829 155091 128863 155329
rect 133153 155227 133187 155261
rect 132911 155193 133187 155227
rect 137109 155261 137385 155295
rect 137109 155227 137143 155261
rect 127725 154683 127759 155057
rect 137385 154819 137419 155125
rect 137477 154819 137511 155329
rect 138029 155295 138063 155465
rect 143733 155431 143767 155533
rect 145423 155397 145757 155431
rect 146861 155159 146895 155329
rect 143641 154955 143675 155125
rect 146953 155159 146987 155873
rect 153393 155567 153427 155737
rect 143549 154887 143583 154921
rect 143733 154887 143767 155125
rect 143549 154853 143767 154887
rect 147137 154139 147171 155465
rect 156153 155023 156187 155533
rect 156429 154955 156463 155873
rect 169861 155771 169895 155873
rect 158821 155363 158855 155737
rect 172897 155703 172931 155873
rect 185685 155159 185719 155873
rect 171149 154887 171183 154989
rect 190469 154887 190503 155873
rect 195253 154615 195287 154989
rect 197461 154887 197495 155873
rect 202061 155431 202095 155873
rect 202153 155227 202187 155397
rect 197553 154683 197587 154853
rect 202981 154683 203015 155057
rect 203073 154683 203107 155261
rect 204821 154819 204855 155873
rect 205925 155261 206143 155295
rect 205925 154683 205959 155261
rect 206109 155227 206143 155261
rect 204947 154649 205189 154683
rect 206017 154615 206051 155193
rect 209881 155091 209915 155397
rect 213193 155295 213227 155805
rect 213837 154615 213871 156757
rect 220737 156451 220771 156757
rect 214297 155975 214331 156009
rect 214147 155941 214331 155975
rect 229235 155737 229419 155771
rect 214481 155091 214515 155261
rect 214573 154683 214607 155057
rect 214665 154683 214699 155329
rect 221565 155295 221599 155601
rect 221657 155499 221691 155601
rect 219357 154615 219391 155261
rect 223589 155295 223623 155397
rect 224141 155363 224175 155601
rect 224233 155363 224267 155533
rect 229385 155363 229419 155737
rect 233801 155737 234111 155771
rect 233801 155363 233835 155737
rect 234077 155703 234111 155737
rect 219449 154615 219483 155261
rect 233893 154615 233927 155329
rect 233985 154615 234019 155669
rect 241069 154887 241103 155737
rect 241989 154955 242023 155125
rect 242081 154955 242115 155873
rect 243553 155023 243587 155669
rect 248981 155499 249015 155873
rect 262815 155805 262907 155839
rect 244933 154887 244967 155057
rect 248889 154887 248923 155465
rect 249073 155193 249257 155227
rect 249073 155091 249107 155193
rect 258641 155091 258675 155329
rect 258641 155057 259469 155091
rect 244323 154853 244599 154887
rect 244473 154751 244507 154785
rect 244323 154717 244507 154751
rect 244565 154751 244599 154853
rect 163823 154377 164157 154411
rect 159741 154275 159775 154377
rect 166917 154207 166951 154513
rect 248797 154479 248831 154853
rect 252695 154717 252845 154751
rect 254777 154683 254811 154785
rect 256559 154717 256709 154751
rect 261309 154615 261343 154649
rect 261309 154581 261493 154615
rect 169711 154309 170263 154343
rect 140823 154105 141099 154139
rect 141065 154071 141099 154105
rect 137235 154037 137477 154071
rect 144745 154003 144779 154105
rect 146953 153935 146987 154037
rect 149345 154003 149379 154105
rect 108313 153323 108347 153425
rect 113557 153255 113591 153425
rect 113649 153323 113683 153425
rect 120181 153391 120215 153493
rect 120123 153357 120215 153391
rect 114937 153323 114971 153357
rect 166273 153323 166307 154173
rect 168113 154139 168147 154309
rect 170229 154139 170263 154309
rect 175933 153459 175967 153697
rect 262689 153391 262723 155057
rect 262781 154887 262815 155057
rect 262873 154751 262907 155805
rect 262965 155227 262999 155873
rect 286977 155703 287011 156009
rect 296729 155941 296821 155975
rect 277409 155669 277593 155703
rect 264161 155227 264195 155329
rect 262873 154717 262965 154751
rect 268301 154479 268335 154989
rect 272441 154479 272475 154989
rect 272533 154751 272567 154989
rect 272625 154751 272659 155193
rect 272717 154887 272751 155329
rect 277409 155159 277443 155669
rect 277501 155023 277535 155125
rect 277443 154989 277535 155023
rect 276213 154819 276247 154921
rect 276121 154615 276155 154785
rect 280077 154751 280111 155601
rect 282009 155499 282043 155669
rect 287897 155567 287931 155805
rect 281825 154275 281859 154717
rect 282009 154207 282043 154785
rect 282101 154683 282135 155057
rect 282193 154955 282227 155125
rect 282285 154819 282319 154921
rect 285781 154819 285815 154989
rect 282101 154649 282285 154683
rect 287805 154615 287839 155533
rect 288909 155363 288943 155533
rect 288725 155159 288759 155329
rect 288633 154887 288667 155125
rect 288541 154615 288575 154853
rect 289829 154683 289863 155873
rect 292865 155091 292899 155533
rect 296729 155431 296763 155941
rect 296821 155295 296855 155397
rect 296763 155261 296855 155295
rect 298661 155159 298695 155397
rect 291853 154615 291887 155057
rect 296671 154853 296729 154887
rect 288541 154581 288633 154615
rect 296913 154479 296947 154921
rect 300593 154751 300627 155737
rect 302341 155703 302375 156009
rect 302525 155635 302559 155941
rect 302283 155601 302375 155635
rect 301363 155329 301547 155363
rect 301513 155159 301547 155329
rect 301421 154411 301455 155125
rect 302341 155091 302375 155601
rect 303261 155567 303295 155805
rect 306849 155703 306883 155941
rect 302525 154955 302559 155397
rect 303445 154819 303479 155465
rect 304457 154615 304491 155601
rect 306941 155159 306975 155669
rect 307033 155567 307067 155873
rect 306941 154819 306975 154989
rect 307033 154683 307067 154853
rect 307125 154683 307159 155261
rect 307217 155159 307251 155737
rect 308137 155499 308171 156009
rect 313381 155567 313415 155873
rect 407957 155703 407991 155873
rect 412465 155635 412499 155941
rect 319085 154819 319119 155533
rect 412557 155499 412591 155737
rect 412407 155465 412591 155499
rect 402253 154819 402287 154989
rect 409889 154955 409923 155125
rect 417341 154751 417375 155737
rect 417433 154819 417467 155533
rect 420837 154751 420871 154921
rect 317187 154581 317429 154615
rect 433349 154479 433383 154649
rect 395537 154207 395571 154377
rect 324973 153459 325007 153629
rect 114937 153289 115121 153323
rect 124873 153289 125057 153323
rect 113741 153255 113775 153289
rect 113557 153221 113775 153255
rect 124873 153255 124907 153289
rect 127483 152677 127633 152711
rect 158453 152439 158487 153017
rect 195253 151963 195287 152677
rect 214573 151963 214607 152541
rect 491033 152167 491067 152473
rect 40141 150943 40175 151385
rect 41337 151079 41371 151793
rect 75193 151079 75227 151861
rect 78137 151011 78171 151861
rect 88349 150467 88383 151861
rect 91937 150535 91971 151861
rect 95157 151147 95191 151861
rect 99297 151215 99331 151861
rect 105645 150603 105679 151793
rect 127541 151521 127725 151555
rect 127541 151487 127575 151521
rect 506949 151283 506983 151589
rect 508881 151079 508915 151317
rect 578249 52411 578283 155533
rect 12173 4471 12207 4777
rect 62681 4403 62715 4845
rect 79333 4403 79367 4981
rect 95985 4335 96019 5049
rect 444389 4675 444423 5117
rect 463341 4675 463375 5117
rect 130669 2975 130703 3349
rect 407715 3349 407899 3383
rect 404829 3179 404863 3349
rect 407865 3247 407899 3349
rect 417433 3179 417467 3281
rect 407405 3043 407439 3145
rect 417525 3043 417559 3145
rect 108313 1887 108347 2125
rect 115489 1853 115765 1887
rect 115489 1819 115523 1853
<< viali >>
rect 173081 157301 173115 157335
rect 182005 157301 182039 157335
rect 172897 157233 172931 157267
rect 173449 157233 173483 157267
rect 173449 156553 173483 156587
rect 173725 157165 173759 157199
rect 173725 156553 173759 156587
rect 175933 157029 175967 157063
rect 175933 156553 175967 156587
rect 185685 157301 185719 157335
rect 185501 157165 185535 157199
rect 182005 156417 182039 156451
rect 185501 157029 185535 157063
rect 185593 157029 185627 157063
rect 185685 156349 185719 156383
rect 185777 157233 185811 157267
rect 213745 156757 213779 156791
rect 204913 156689 204947 156723
rect 185409 156281 185443 156315
rect 185501 156281 185535 156315
rect 195161 156485 195195 156519
rect 204913 156417 204947 156451
rect 205005 156485 205039 156519
rect 195161 156213 195195 156247
rect 195253 156349 195287 156383
rect 195253 156213 195287 156247
rect 195345 156349 195379 156383
rect 194885 156145 194919 156179
rect 213745 156417 213779 156451
rect 213837 156757 213871 156791
rect 205005 156145 205039 156179
rect 113281 156077 113315 156111
rect 146953 155873 146987 155907
rect 113281 155805 113315 155839
rect 118065 155805 118099 155839
rect 117973 155601 118007 155635
rect 118065 155601 118099 155635
rect 127541 155805 127575 155839
rect 117881 155261 117915 155295
rect 117973 155261 118007 155295
rect 124781 155193 124815 155227
rect 124781 155057 124815 155091
rect 127449 155057 127483 155091
rect 127541 155057 127575 155091
rect 127633 155805 127667 155839
rect 117881 154717 117915 154751
rect 137109 155669 137143 155703
rect 133889 155465 133923 155499
rect 143733 155533 143767 155567
rect 137109 155397 137143 155431
rect 138029 155465 138063 155499
rect 128829 155329 128863 155363
rect 133889 155329 133923 155363
rect 137201 155329 137235 155363
rect 133153 155261 133187 155295
rect 132877 155193 132911 155227
rect 137385 155261 137419 155295
rect 137109 155193 137143 155227
rect 127633 154649 127667 154683
rect 127725 155057 127759 155091
rect 128829 155057 128863 155091
rect 137385 155125 137419 155159
rect 137385 154785 137419 154819
rect 143733 155397 143767 155431
rect 145389 155397 145423 155431
rect 145757 155397 145791 155431
rect 138029 155261 138063 155295
rect 146861 155329 146895 155363
rect 143641 155125 143675 155159
rect 143549 154921 143583 154955
rect 143641 154921 143675 154955
rect 143733 155125 143767 155159
rect 146861 155125 146895 155159
rect 156429 155873 156463 155907
rect 153393 155737 153427 155771
rect 153393 155533 153427 155567
rect 156153 155533 156187 155567
rect 146953 155125 146987 155159
rect 147137 155465 147171 155499
rect 137477 154785 137511 154819
rect 127725 154649 127759 154683
rect 156153 154989 156187 155023
rect 169861 155873 169895 155907
rect 158821 155737 158855 155771
rect 169861 155737 169895 155771
rect 172897 155873 172931 155907
rect 172897 155669 172931 155703
rect 185685 155873 185719 155907
rect 158821 155329 158855 155363
rect 185685 155125 185719 155159
rect 190469 155873 190503 155907
rect 156429 154921 156463 154955
rect 171149 154989 171183 155023
rect 171149 154853 171183 154887
rect 197461 155873 197495 155907
rect 190469 154853 190503 154887
rect 195253 154989 195287 155023
rect 202061 155873 202095 155907
rect 204821 155873 204855 155907
rect 202061 155397 202095 155431
rect 202153 155397 202187 155431
rect 202153 155193 202187 155227
rect 203073 155261 203107 155295
rect 202981 155057 203015 155091
rect 197461 154853 197495 154887
rect 197553 154853 197587 154887
rect 197553 154649 197587 154683
rect 202981 154649 203015 154683
rect 213193 155805 213227 155839
rect 209881 155397 209915 155431
rect 204821 154785 204855 154819
rect 203073 154649 203107 154683
rect 204913 154649 204947 154683
rect 205189 154649 205223 154683
rect 205925 154649 205959 154683
rect 206017 155193 206051 155227
rect 206109 155193 206143 155227
rect 195253 154581 195287 154615
rect 213193 155261 213227 155295
rect 209881 155057 209915 155091
rect 206017 154581 206051 154615
rect 220737 156757 220771 156791
rect 220737 156417 220771 156451
rect 214297 156009 214331 156043
rect 214113 155941 214147 155975
rect 286977 156009 287011 156043
rect 242081 155873 242115 155907
rect 229201 155737 229235 155771
rect 221565 155601 221599 155635
rect 214665 155329 214699 155363
rect 214481 155261 214515 155295
rect 214481 155057 214515 155091
rect 214573 155057 214607 155091
rect 214573 154649 214607 154683
rect 221657 155601 221691 155635
rect 221657 155465 221691 155499
rect 224141 155601 224175 155635
rect 214665 154649 214699 154683
rect 219357 155261 219391 155295
rect 213837 154581 213871 154615
rect 219357 154581 219391 154615
rect 219449 155261 219483 155295
rect 221565 155261 221599 155295
rect 223589 155397 223623 155431
rect 224141 155329 224175 155363
rect 224233 155533 224267 155567
rect 224233 155329 224267 155363
rect 229385 155329 229419 155363
rect 233985 155669 234019 155703
rect 234077 155669 234111 155703
rect 241069 155737 241103 155771
rect 233801 155329 233835 155363
rect 233893 155329 233927 155363
rect 223589 155261 223623 155295
rect 219449 154581 219483 154615
rect 233893 154581 233927 154615
rect 241989 155125 242023 155159
rect 241989 154921 242023 154955
rect 248981 155873 249015 155907
rect 243553 155669 243587 155703
rect 262965 155873 262999 155907
rect 262781 155805 262815 155839
rect 248889 155465 248923 155499
rect 248981 155465 249015 155499
rect 243553 154989 243587 155023
rect 244933 155057 244967 155091
rect 242081 154921 242115 154955
rect 258641 155329 258675 155363
rect 249257 155193 249291 155227
rect 249073 155057 249107 155091
rect 259469 155057 259503 155091
rect 262689 155057 262723 155091
rect 241069 154853 241103 154887
rect 244289 154853 244323 154887
rect 244933 154853 244967 154887
rect 248797 154853 248831 154887
rect 248889 154853 248923 154887
rect 244473 154785 244507 154819
rect 244289 154717 244323 154751
rect 244565 154717 244599 154751
rect 233985 154581 234019 154615
rect 166917 154513 166951 154547
rect 159741 154377 159775 154411
rect 163789 154377 163823 154411
rect 164157 154377 164191 154411
rect 159741 154241 159775 154275
rect 254777 154785 254811 154819
rect 252661 154717 252695 154751
rect 252845 154717 252879 154751
rect 256525 154717 256559 154751
rect 256709 154717 256743 154751
rect 254777 154649 254811 154683
rect 261309 154649 261343 154683
rect 261493 154581 261527 154615
rect 248797 154445 248831 154479
rect 166273 154173 166307 154207
rect 166917 154173 166951 154207
rect 168113 154309 168147 154343
rect 169677 154309 169711 154343
rect 140789 154105 140823 154139
rect 137201 154037 137235 154071
rect 137477 154037 137511 154071
rect 141065 154037 141099 154071
rect 144745 154105 144779 154139
rect 147137 154105 147171 154139
rect 149345 154105 149379 154139
rect 144745 153969 144779 154003
rect 146953 154037 146987 154071
rect 149345 153969 149379 154003
rect 146953 153901 146987 153935
rect 127449 153833 127483 153867
rect 120181 153493 120215 153527
rect 108313 153425 108347 153459
rect 108313 153289 108347 153323
rect 113557 153425 113591 153459
rect 113649 153425 113683 153459
rect 114937 153357 114971 153391
rect 120089 153357 120123 153391
rect 168113 154105 168147 154139
rect 170229 154105 170263 154139
rect 175933 153697 175967 153731
rect 175933 153425 175967 153459
rect 262781 155057 262815 155091
rect 262781 154853 262815 154887
rect 302341 156009 302375 156043
rect 296821 155941 296855 155975
rect 289829 155873 289863 155907
rect 277593 155669 277627 155703
rect 282009 155669 282043 155703
rect 286977 155669 287011 155703
rect 287897 155805 287931 155839
rect 262965 155193 262999 155227
rect 264161 155329 264195 155363
rect 272717 155329 272751 155363
rect 264161 155193 264195 155227
rect 272625 155193 272659 155227
rect 268301 154989 268335 155023
rect 262965 154717 262999 154751
rect 268301 154445 268335 154479
rect 272441 154989 272475 155023
rect 272533 154989 272567 155023
rect 272533 154717 272567 154751
rect 280077 155601 280111 155635
rect 277409 155125 277443 155159
rect 277501 155125 277535 155159
rect 277409 154989 277443 155023
rect 272717 154853 272751 154887
rect 276213 154921 276247 154955
rect 272625 154717 272659 154751
rect 276121 154785 276155 154819
rect 276213 154785 276247 154819
rect 282009 155465 282043 155499
rect 287805 155533 287839 155567
rect 287897 155533 287931 155567
rect 288909 155533 288943 155567
rect 282193 155125 282227 155159
rect 282101 155057 282135 155091
rect 282009 154785 282043 154819
rect 280077 154717 280111 154751
rect 281825 154717 281859 154751
rect 276121 154581 276155 154615
rect 272441 154445 272475 154479
rect 281825 154241 281859 154275
rect 285781 154989 285815 155023
rect 282193 154921 282227 154955
rect 282285 154921 282319 154955
rect 282285 154785 282319 154819
rect 285781 154785 285815 154819
rect 282285 154649 282319 154683
rect 288725 155329 288759 155363
rect 288909 155329 288943 155363
rect 288633 155125 288667 155159
rect 288725 155125 288759 155159
rect 287805 154581 287839 154615
rect 288541 154853 288575 154887
rect 288633 154853 288667 154887
rect 292865 155533 292899 155567
rect 300593 155737 300627 155771
rect 296729 155397 296763 155431
rect 296821 155397 296855 155431
rect 296729 155261 296763 155295
rect 298661 155397 298695 155431
rect 298661 155125 298695 155159
rect 289829 154649 289863 154683
rect 291853 155057 291887 155091
rect 292865 155057 292899 155091
rect 296913 154921 296947 154955
rect 296637 154853 296671 154887
rect 296729 154853 296763 154887
rect 288633 154581 288667 154615
rect 291853 154581 291887 154615
rect 308137 156009 308171 156043
rect 302341 155669 302375 155703
rect 302525 155941 302559 155975
rect 306849 155941 306883 155975
rect 302249 155601 302283 155635
rect 302525 155601 302559 155635
rect 303261 155805 303295 155839
rect 301329 155329 301363 155363
rect 300593 154717 300627 154751
rect 301421 155125 301455 155159
rect 301513 155125 301547 155159
rect 296913 154445 296947 154479
rect 307033 155873 307067 155907
rect 306849 155669 306883 155703
rect 306941 155669 306975 155703
rect 303261 155533 303295 155567
rect 304457 155601 304491 155635
rect 303445 155465 303479 155499
rect 302341 155057 302375 155091
rect 302525 155397 302559 155431
rect 302525 154921 302559 154955
rect 303445 154785 303479 154819
rect 307033 155533 307067 155567
rect 307217 155737 307251 155771
rect 306941 155125 306975 155159
rect 307125 155261 307159 155295
rect 306941 154989 306975 155023
rect 306941 154785 306975 154819
rect 307033 154853 307067 154887
rect 307033 154649 307067 154683
rect 412465 155941 412499 155975
rect 313381 155873 313415 155907
rect 407957 155873 407991 155907
rect 407957 155669 407991 155703
rect 412465 155601 412499 155635
rect 412557 155737 412591 155771
rect 313381 155533 313415 155567
rect 319085 155533 319119 155567
rect 308137 155465 308171 155499
rect 307217 155125 307251 155159
rect 412373 155465 412407 155499
rect 417341 155737 417375 155771
rect 409889 155125 409923 155159
rect 319085 154785 319119 154819
rect 402253 154989 402287 155023
rect 409889 154921 409923 154955
rect 402253 154785 402287 154819
rect 417433 155533 417467 155567
rect 578249 155533 578283 155567
rect 417433 154785 417467 154819
rect 420837 154921 420871 154955
rect 417341 154717 417375 154751
rect 420837 154717 420871 154751
rect 307125 154649 307159 154683
rect 433349 154649 433383 154683
rect 304457 154581 304491 154615
rect 317153 154581 317187 154615
rect 317429 154581 317463 154615
rect 433349 154445 433383 154479
rect 301421 154377 301455 154411
rect 395537 154377 395571 154411
rect 282009 154173 282043 154207
rect 395537 154173 395571 154207
rect 324973 153629 325007 153663
rect 324973 153425 325007 153459
rect 262689 153357 262723 153391
rect 113649 153289 113683 153323
rect 113741 153289 113775 153323
rect 115121 153289 115155 153323
rect 125057 153289 125091 153323
rect 166273 153289 166307 153323
rect 124873 153221 124907 153255
rect 158453 153017 158487 153051
rect 127449 152677 127483 152711
rect 127633 152677 127667 152711
rect 158453 152405 158487 152439
rect 195253 152677 195287 152711
rect 195253 151929 195287 151963
rect 214573 152541 214607 152575
rect 491033 152473 491067 152507
rect 491033 152133 491067 152167
rect 214573 151929 214607 151963
rect 75193 151861 75227 151895
rect 41337 151793 41371 151827
rect 40141 151385 40175 151419
rect 41337 151045 41371 151079
rect 75193 151045 75227 151079
rect 78137 151861 78171 151895
rect 78137 150977 78171 151011
rect 88349 151861 88383 151895
rect 40141 150909 40175 150943
rect 91937 151861 91971 151895
rect 95157 151861 95191 151895
rect 99297 151861 99331 151895
rect 99297 151181 99331 151215
rect 105645 151793 105679 151827
rect 95157 151113 95191 151147
rect 506949 151589 506983 151623
rect 127725 151521 127759 151555
rect 127541 151453 127575 151487
rect 506949 151249 506983 151283
rect 508881 151317 508915 151351
rect 508881 151045 508915 151079
rect 105645 150569 105679 150603
rect 91937 150501 91971 150535
rect 88349 150433 88383 150467
rect 578249 52377 578283 52411
rect 444389 5117 444423 5151
rect 95985 5049 96019 5083
rect 79333 4981 79367 5015
rect 62681 4845 62715 4879
rect 12173 4777 12207 4811
rect 12173 4437 12207 4471
rect 62681 4369 62715 4403
rect 79333 4369 79367 4403
rect 444389 4641 444423 4675
rect 463341 5117 463375 5151
rect 463341 4641 463375 4675
rect 95985 4301 96019 4335
rect 130669 3349 130703 3383
rect 404829 3349 404863 3383
rect 407681 3349 407715 3383
rect 407865 3213 407899 3247
rect 417433 3281 417467 3315
rect 404829 3145 404863 3179
rect 407405 3145 407439 3179
rect 417433 3145 417467 3179
rect 417525 3145 417559 3179
rect 407405 3009 407439 3043
rect 417525 3009 417559 3043
rect 130669 2941 130703 2975
rect 108313 2125 108347 2159
rect 108313 1853 108347 1887
rect 115765 1853 115799 1887
rect 115489 1785 115523 1819
<< metal1 >>
rect 38470 158924 38476 158976
rect 38528 158964 38534 158976
rect 145282 158964 145288 158976
rect 38528 158936 145288 158964
rect 38528 158924 38534 158936
rect 145282 158924 145288 158936
rect 145340 158924 145346 158976
rect 34514 158856 34520 158908
rect 34572 158896 34578 158908
rect 142798 158896 142804 158908
rect 34572 158868 142804 158896
rect 34572 158856 34578 158868
rect 142798 158856 142804 158868
rect 142856 158856 142862 158908
rect 30650 158788 30656 158840
rect 30708 158828 30714 158840
rect 140130 158828 140136 158840
rect 30708 158800 140136 158828
rect 30708 158788 30714 158800
rect 140130 158788 140136 158800
rect 140188 158788 140194 158840
rect 26786 158720 26792 158772
rect 26844 158760 26850 158772
rect 137462 158760 137468 158772
rect 26844 158732 137468 158760
rect 26844 158720 26850 158732
rect 137462 158720 137468 158732
rect 137520 158720 137526 158772
rect 11146 158652 11152 158704
rect 11204 158692 11210 158704
rect 127066 158692 127072 158704
rect 11204 158664 127072 158692
rect 11204 158652 11210 158664
rect 127066 158652 127072 158664
rect 127124 158652 127130 158704
rect 22830 158584 22836 158636
rect 22888 158624 22894 158636
rect 134886 158624 134892 158636
rect 22888 158596 134892 158624
rect 22888 158584 22894 158596
rect 134886 158584 134892 158596
rect 134944 158584 134950 158636
rect 70578 158516 70584 158568
rect 70636 158556 70642 158568
rect 167270 158556 167276 158568
rect 70636 158528 167276 158556
rect 70636 158516 70642 158528
rect 167270 158516 167276 158528
rect 167328 158516 167334 158568
rect 66714 158448 66720 158500
rect 66772 158488 66778 158500
rect 164234 158488 164240 158500
rect 66772 158460 164240 158488
rect 66772 158448 66778 158460
rect 164234 158448 164240 158460
rect 164292 158448 164298 158500
rect 62850 158380 62856 158432
rect 62908 158420 62914 158432
rect 161658 158420 161664 158432
rect 62908 158392 161664 158420
rect 62908 158380 62914 158392
rect 161658 158380 161664 158392
rect 161716 158380 161722 158432
rect 55214 158312 55220 158364
rect 55272 158352 55278 158364
rect 156322 158352 156328 158364
rect 55272 158324 156328 158352
rect 55272 158312 55278 158324
rect 156322 158312 156328 158324
rect 156380 158312 156386 158364
rect 18966 158244 18972 158296
rect 19024 158284 19030 158296
rect 132586 158284 132592 158296
rect 19024 158256 132592 158284
rect 19024 158244 19030 158256
rect 132586 158244 132592 158256
rect 132644 158244 132650 158296
rect 104710 158176 104716 158228
rect 104768 158216 104774 158228
rect 189626 158216 189632 158228
rect 104768 158188 189632 158216
rect 104768 158176 104774 158188
rect 189626 158176 189632 158188
rect 189684 158176 189690 158228
rect 90082 158108 90088 158160
rect 90140 158148 90146 158160
rect 179874 158148 179880 158160
rect 90140 158120 179880 158148
rect 90140 158108 90146 158120
rect 179874 158108 179880 158120
rect 179932 158108 179938 158160
rect 58894 158040 58900 158092
rect 58952 158080 58958 158092
rect 158990 158080 158996 158092
rect 58952 158052 158996 158080
rect 58952 158040 58958 158052
rect 158990 158040 158996 158052
rect 159048 158040 159054 158092
rect 51074 157972 51080 158024
rect 51132 158012 51138 158024
rect 153746 158012 153752 158024
rect 51132 157984 153752 158012
rect 51132 157972 51138 157984
rect 153746 157972 153752 157984
rect 153804 157972 153810 158024
rect 47210 157904 47216 157956
rect 47268 157944 47274 157956
rect 151170 157944 151176 157956
rect 47268 157916 151176 157944
rect 47268 157904 47274 157916
rect 151170 157904 151176 157916
rect 151228 157904 151234 157956
rect 43346 157836 43352 157888
rect 43404 157876 43410 157888
rect 148502 157876 148508 157888
rect 43404 157848 148508 157876
rect 43404 157836 43410 157848
rect 148502 157836 148508 157848
rect 148560 157836 148566 157888
rect 148594 157836 148600 157888
rect 148652 157876 148658 157888
rect 218882 157876 218888 157888
rect 148652 157848 218888 157876
rect 148652 157836 148658 157848
rect 218882 157836 218888 157848
rect 218940 157836 218946 157888
rect 15010 157768 15016 157820
rect 15068 157808 15074 157820
rect 129734 157808 129740 157820
rect 15068 157780 129740 157808
rect 15068 157768 15074 157780
rect 129734 157768 129740 157780
rect 129792 157768 129798 157820
rect 132034 157768 132040 157820
rect 132092 157808 132098 157820
rect 207750 157808 207756 157820
rect 132092 157780 207756 157808
rect 132092 157768 132098 157780
rect 207750 157768 207756 157780
rect 207808 157768 207814 157820
rect 144730 157700 144736 157752
rect 144788 157740 144794 157752
rect 216214 157740 216220 157752
rect 144788 157712 216220 157740
rect 144788 157700 144794 157712
rect 216214 157700 216220 157712
rect 216272 157700 216278 157752
rect 129090 157632 129096 157684
rect 129148 157672 129154 157684
rect 205818 157672 205824 157684
rect 129148 157644 205824 157672
rect 129148 157632 129154 157644
rect 205818 157632 205824 157644
rect 205876 157632 205882 157684
rect 117406 157564 117412 157616
rect 117464 157604 117470 157616
rect 197998 157604 198004 157616
rect 117464 157576 198004 157604
rect 117464 157564 117470 157576
rect 197998 157564 198004 157576
rect 198056 157564 198062 157616
rect 108666 157496 108672 157548
rect 108724 157536 108730 157548
rect 192110 157536 192116 157548
rect 108724 157508 192116 157536
rect 108724 157496 108730 157508
rect 192110 157496 192116 157508
rect 192168 157496 192174 157548
rect 100846 157428 100852 157480
rect 100904 157468 100910 157480
rect 186958 157468 186964 157480
rect 100904 157440 186964 157468
rect 100904 157428 100910 157440
rect 186958 157428 186964 157440
rect 187016 157428 187022 157480
rect 119430 157360 119436 157412
rect 119488 157400 119494 157412
rect 510154 157400 510160 157412
rect 119488 157372 510160 157400
rect 119488 157360 119494 157372
rect 510154 157360 510160 157372
rect 510212 157360 510218 157412
rect 84286 157292 84292 157344
rect 84344 157332 84350 157344
rect 173069 157335 173127 157341
rect 84344 157304 173020 157332
rect 84344 157292 84350 157304
rect 82262 157224 82268 157276
rect 82320 157264 82326 157276
rect 172885 157267 172943 157273
rect 172885 157264 172897 157267
rect 82320 157236 172897 157264
rect 82320 157224 82326 157236
rect 172885 157233 172897 157236
rect 172931 157233 172943 157267
rect 172885 157227 172943 157233
rect 77478 157156 77484 157208
rect 77536 157196 77542 157208
rect 171410 157196 171416 157208
rect 77536 157168 171416 157196
rect 77536 157156 77542 157168
rect 171410 157156 171416 157168
rect 171468 157156 171474 157208
rect 172992 157196 173020 157304
rect 173069 157301 173081 157335
rect 173115 157332 173127 157335
rect 174538 157332 174544 157344
rect 173115 157304 174544 157332
rect 173115 157301 173127 157304
rect 173069 157295 173127 157301
rect 174538 157292 174544 157304
rect 174596 157292 174602 157344
rect 181993 157335 182051 157341
rect 181993 157301 182005 157335
rect 182039 157332 182051 157335
rect 185673 157335 185731 157341
rect 182039 157304 185624 157332
rect 182039 157301 182051 157304
rect 181993 157295 182051 157301
rect 173437 157267 173495 157273
rect 173437 157233 173449 157267
rect 173483 157264 173495 157267
rect 181070 157264 181076 157276
rect 173483 157236 181076 157264
rect 173483 157233 173495 157236
rect 173437 157227 173495 157233
rect 181070 157224 181076 157236
rect 181128 157224 181134 157276
rect 173713 157199 173771 157205
rect 173713 157196 173725 157199
rect 172992 157168 173725 157196
rect 173713 157165 173725 157168
rect 173759 157165 173771 157199
rect 173713 157159 173771 157165
rect 173894 157156 173900 157208
rect 173952 157196 173958 157208
rect 185489 157199 185547 157205
rect 185489 157196 185501 157199
rect 173952 157168 185501 157196
rect 173952 157156 173958 157168
rect 185489 157165 185501 157168
rect 185535 157165 185547 157199
rect 185596 157196 185624 157304
rect 185673 157301 185685 157335
rect 185719 157332 185731 157335
rect 190454 157332 190460 157344
rect 185719 157304 190460 157332
rect 185719 157301 185731 157304
rect 185673 157295 185731 157301
rect 190454 157292 190460 157304
rect 190512 157292 190518 157344
rect 201218 157292 201224 157344
rect 201276 157332 201282 157344
rect 253934 157332 253940 157344
rect 201276 157304 253940 157332
rect 201276 157292 201282 157304
rect 253934 157292 253940 157304
rect 253992 157292 253998 157344
rect 426250 157292 426256 157344
rect 426308 157332 426314 157344
rect 458542 157332 458548 157344
rect 426308 157304 458548 157332
rect 426308 157292 426314 157304
rect 458542 157292 458548 157304
rect 458600 157292 458606 157344
rect 472434 157292 472440 157344
rect 472492 157332 472498 157344
rect 527726 157332 527732 157344
rect 472492 157304 527732 157332
rect 472492 157292 472498 157304
rect 527726 157292 527732 157304
rect 527784 157292 527790 157344
rect 185765 157267 185823 157273
rect 185765 157233 185777 157267
rect 185811 157264 185823 157267
rect 191558 157264 191564 157276
rect 185811 157236 191564 157264
rect 185811 157233 185823 157236
rect 185765 157227 185823 157233
rect 191558 157224 191564 157236
rect 191616 157224 191622 157276
rect 193398 157224 193404 157276
rect 193456 157264 193462 157276
rect 248690 157264 248696 157276
rect 193456 157236 248696 157264
rect 193456 157224 193462 157236
rect 248690 157224 248696 157236
rect 248748 157224 248754 157276
rect 428918 157224 428924 157276
rect 428976 157264 428982 157276
rect 462498 157264 462504 157276
rect 428976 157236 462504 157264
rect 428976 157224 428982 157236
rect 462498 157224 462504 157236
rect 462556 157224 462562 157276
rect 473722 157224 473728 157276
rect 473780 157264 473786 157276
rect 529750 157264 529756 157276
rect 473780 157236 529756 157264
rect 473780 157224 473786 157236
rect 529750 157224 529756 157236
rect 529808 157224 529814 157276
rect 189074 157196 189080 157208
rect 185596 157168 189080 157196
rect 185489 157159 185547 157165
rect 189074 157156 189080 157168
rect 189132 157156 189138 157208
rect 189534 157156 189540 157208
rect 189592 157196 189598 157208
rect 246114 157196 246120 157208
rect 189592 157168 246120 157196
rect 189592 157156 189598 157168
rect 246114 157156 246120 157168
rect 246172 157156 246178 157208
rect 442534 157156 442540 157208
rect 442592 157196 442598 157208
rect 482922 157196 482928 157208
rect 442592 157168 482928 157196
rect 442592 157156 442598 157168
rect 482922 157156 482928 157168
rect 482980 157156 482986 157208
rect 484946 157156 484952 157208
rect 485004 157196 485010 157208
rect 540422 157196 540428 157208
rect 485004 157168 540428 157196
rect 485004 157156 485010 157168
rect 540422 157156 540428 157168
rect 540480 157156 540486 157208
rect 76466 157088 76472 157140
rect 76524 157128 76530 157140
rect 170674 157128 170680 157140
rect 76524 157100 170680 157128
rect 76524 157088 76530 157100
rect 170674 157088 170680 157100
rect 170732 157088 170738 157140
rect 173802 157088 173808 157140
rect 173860 157128 173866 157140
rect 173860 157100 176056 157128
rect 173860 157088 173866 157100
rect 69658 157020 69664 157072
rect 69716 157060 69722 157072
rect 166074 157060 166080 157072
rect 69716 157032 166080 157060
rect 69716 157020 69722 157032
rect 166074 157020 166080 157032
rect 166132 157020 166138 157072
rect 169754 157020 169760 157072
rect 169812 157060 169818 157072
rect 175921 157063 175979 157069
rect 175921 157060 175933 157063
rect 169812 157032 175933 157060
rect 169812 157020 169818 157032
rect 175921 157029 175933 157032
rect 175967 157029 175979 157063
rect 176028 157060 176056 157100
rect 177850 157088 177856 157140
rect 177908 157128 177914 157140
rect 238386 157128 238392 157140
rect 177908 157100 238392 157128
rect 177908 157088 177914 157100
rect 238386 157088 238392 157100
rect 238444 157088 238450 157140
rect 251910 157088 251916 157140
rect 251968 157128 251974 157140
rect 287790 157128 287796 157140
rect 251968 157100 287796 157128
rect 251968 157088 251974 157100
rect 287790 157088 287796 157100
rect 287848 157088 287854 157140
rect 434622 157088 434628 157140
rect 434680 157128 434686 157140
rect 471238 157128 471244 157140
rect 434680 157100 471244 157128
rect 434680 157088 434686 157100
rect 471238 157088 471244 157100
rect 471296 157088 471302 157140
rect 474458 157088 474464 157140
rect 474516 157128 474522 157140
rect 530670 157128 530676 157140
rect 474516 157100 530676 157128
rect 474516 157088 474522 157100
rect 530670 157088 530676 157100
rect 530728 157088 530734 157140
rect 185489 157063 185547 157069
rect 185489 157060 185501 157063
rect 176028 157032 185501 157060
rect 175921 157023 175979 157029
rect 185489 157029 185501 157032
rect 185535 157029 185547 157063
rect 185489 157023 185547 157029
rect 185581 157063 185639 157069
rect 185581 157029 185593 157063
rect 185627 157060 185639 157063
rect 235994 157060 236000 157072
rect 185627 157032 236000 157060
rect 185627 157029 185639 157032
rect 185581 157023 185639 157029
rect 235994 157020 236000 157032
rect 236052 157020 236058 157072
rect 244090 157020 244096 157072
rect 244148 157060 244154 157072
rect 282546 157060 282552 157072
rect 244148 157032 282552 157060
rect 244148 157020 244154 157032
rect 282546 157020 282552 157032
rect 282604 157020 282610 157072
rect 436646 157020 436652 157072
rect 436704 157060 436710 157072
rect 474182 157060 474188 157072
rect 436704 157032 474188 157060
rect 436704 157020 436710 157032
rect 474182 157020 474188 157032
rect 474240 157020 474246 157072
rect 476022 157020 476028 157072
rect 476080 157060 476086 157072
rect 533614 157060 533620 157072
rect 476080 157032 533620 157060
rect 476080 157020 476086 157032
rect 533614 157020 533620 157032
rect 533672 157020 533678 157072
rect 68646 156952 68652 157004
rect 68704 156992 68710 157004
rect 165614 156992 165620 157004
rect 68704 156964 165620 156992
rect 68704 156952 68710 156964
rect 165614 156952 165620 156964
rect 165672 156952 165678 157004
rect 168098 156952 168104 157004
rect 168156 156992 168162 157004
rect 231854 156992 231860 157004
rect 168156 156964 231860 156992
rect 168156 156952 168162 156964
rect 231854 156952 231860 156964
rect 231912 156952 231918 157004
rect 240226 156952 240232 157004
rect 240284 156992 240290 157004
rect 280246 156992 280252 157004
rect 240284 156964 280252 156992
rect 240284 156952 240290 156964
rect 280246 156952 280252 156964
rect 280304 156952 280310 157004
rect 437382 156952 437388 157004
rect 437440 156992 437446 157004
rect 475102 156992 475108 157004
rect 437440 156964 475108 156992
rect 437440 156952 437446 156964
rect 475102 156952 475108 156964
rect 475160 156952 475166 157004
rect 476942 156952 476948 157004
rect 477000 156992 477006 157004
rect 534626 156992 534632 157004
rect 477000 156964 534632 156992
rect 477000 156952 477006 156964
rect 534626 156952 534632 156964
rect 534684 156952 534690 157004
rect 54018 156884 54024 156936
rect 54076 156924 54082 156936
rect 155954 156924 155960 156936
rect 54076 156896 155960 156924
rect 54076 156884 54082 156896
rect 155954 156884 155960 156896
rect 156012 156884 156018 156936
rect 166166 156884 166172 156936
rect 166224 156924 166230 156936
rect 230566 156924 230572 156936
rect 166224 156896 230572 156924
rect 166224 156884 166230 156896
rect 230566 156884 230572 156896
rect 230624 156884 230630 156936
rect 236270 156884 236276 156936
rect 236328 156924 236334 156936
rect 277578 156924 277584 156936
rect 236328 156896 277584 156924
rect 236328 156884 236334 156896
rect 277578 156884 277584 156896
rect 277636 156884 277642 156936
rect 439958 156884 439964 156936
rect 440016 156924 440022 156936
rect 479058 156924 479064 156936
rect 440016 156896 479064 156924
rect 440016 156884 440022 156896
rect 479058 156884 479064 156896
rect 479116 156884 479122 156936
rect 480070 156884 480076 156936
rect 480128 156924 480134 156936
rect 539502 156924 539508 156936
rect 480128 156896 539508 156924
rect 480128 156884 480134 156896
rect 539502 156884 539508 156896
rect 539560 156884 539566 156936
rect 46198 156816 46204 156868
rect 46256 156856 46262 156868
rect 150618 156856 150624 156868
rect 46256 156828 150624 156856
rect 46256 156816 46262 156828
rect 150618 156816 150624 156828
rect 150676 156816 150682 156868
rect 158346 156816 158352 156868
rect 158404 156856 158410 156868
rect 225322 156856 225328 156868
rect 158404 156828 225328 156856
rect 158404 156816 158410 156828
rect 225322 156816 225328 156828
rect 225380 156816 225386 156868
rect 233418 156816 233424 156868
rect 233476 156856 233482 156868
rect 275370 156856 275376 156868
rect 233476 156828 275376 156856
rect 233476 156816 233482 156828
rect 275370 156816 275376 156828
rect 275428 156816 275434 156868
rect 441522 156816 441528 156868
rect 441580 156856 441586 156868
rect 481910 156856 481916 156868
rect 441580 156828 481916 156856
rect 441580 156816 441586 156828
rect 481910 156816 481916 156828
rect 481968 156816 481974 156868
rect 484210 156816 484216 156868
rect 484268 156856 484274 156868
rect 545298 156856 545304 156868
rect 484268 156828 545304 156856
rect 484268 156816 484274 156828
rect 545298 156816 545304 156828
rect 545356 156816 545362 156868
rect 33594 156748 33600 156800
rect 33652 156788 33658 156800
rect 142246 156788 142252 156800
rect 33652 156760 142252 156788
rect 33652 156748 33658 156760
rect 142246 156748 142252 156760
rect 142304 156748 142310 156800
rect 146662 156748 146668 156800
rect 146720 156788 146726 156800
rect 213733 156791 213791 156797
rect 213733 156788 213745 156791
rect 146720 156760 213745 156788
rect 146720 156748 146726 156760
rect 213733 156757 213745 156760
rect 213779 156757 213791 156791
rect 213733 156751 213791 156757
rect 213825 156791 213883 156797
rect 213825 156757 213837 156791
rect 213871 156788 213883 156791
rect 220725 156791 220783 156797
rect 220725 156788 220737 156791
rect 213871 156760 220737 156788
rect 213871 156757 213883 156760
rect 213825 156751 213883 156757
rect 220725 156757 220737 156760
rect 220771 156757 220783 156791
rect 220725 156751 220783 156757
rect 228542 156748 228548 156800
rect 228600 156788 228606 156800
rect 272150 156788 272156 156800
rect 228600 156760 272156 156788
rect 228600 156748 228606 156760
rect 272150 156748 272156 156760
rect 272208 156748 272214 156800
rect 442810 156748 442816 156800
rect 442868 156788 442874 156800
rect 483934 156788 483940 156800
rect 442868 156760 483940 156788
rect 442868 156748 442874 156760
rect 483934 156748 483940 156760
rect 483992 156748 483998 156800
rect 486694 156748 486700 156800
rect 486752 156788 486758 156800
rect 549162 156788 549168 156800
rect 486752 156760 549168 156788
rect 486752 156748 486758 156760
rect 549162 156748 549168 156760
rect 549220 156748 549226 156800
rect 17954 156680 17960 156732
rect 18012 156720 18018 156732
rect 131666 156720 131672 156732
rect 18012 156692 131672 156720
rect 18012 156680 18018 156692
rect 131666 156680 131672 156692
rect 131724 156680 131730 156732
rect 134978 156680 134984 156732
rect 135036 156720 135042 156732
rect 204901 156723 204959 156729
rect 204901 156720 204913 156723
rect 135036 156692 204913 156720
rect 135036 156680 135042 156692
rect 204901 156689 204913 156692
rect 204947 156689 204959 156723
rect 204901 156683 204959 156689
rect 212902 156680 212908 156732
rect 212960 156720 212966 156732
rect 261754 156720 261760 156732
rect 212960 156692 261760 156720
rect 212960 156680 212966 156692
rect 261754 156680 261760 156692
rect 261812 156680 261818 156732
rect 447042 156680 447048 156732
rect 447100 156720 447106 156732
rect 489730 156720 489736 156732
rect 447100 156692 489736 156720
rect 447100 156680 447106 156692
rect 489730 156680 489736 156692
rect 489788 156680 489794 156732
rect 490650 156680 490656 156732
rect 490708 156720 490714 156732
rect 555050 156720 555056 156732
rect 490708 156692 555056 156720
rect 490708 156680 490714 156692
rect 555050 156680 555056 156692
rect 555108 156680 555114 156732
rect 6270 156612 6276 156664
rect 6328 156652 6334 156664
rect 123846 156652 123852 156664
rect 6328 156624 123852 156652
rect 6328 156612 6334 156624
rect 123846 156612 123852 156624
rect 123904 156612 123910 156664
rect 131022 156612 131028 156664
rect 131080 156652 131086 156664
rect 207014 156652 207020 156664
rect 131080 156624 207020 156652
rect 131080 156612 131086 156624
rect 207014 156612 207020 156624
rect 207072 156612 207078 156664
rect 207106 156612 207112 156664
rect 207164 156652 207170 156664
rect 258074 156652 258080 156664
rect 207164 156624 258080 156652
rect 207164 156612 207170 156624
rect 258074 156612 258080 156624
rect 258132 156612 258138 156664
rect 263594 156612 263600 156664
rect 263652 156652 263658 156664
rect 295518 156652 295524 156664
rect 263652 156624 295524 156652
rect 263652 156612 263658 156624
rect 295518 156612 295524 156624
rect 295576 156612 295582 156664
rect 415854 156612 415860 156664
rect 415912 156652 415918 156664
rect 442994 156652 443000 156664
rect 415912 156624 443000 156652
rect 415912 156612 415918 156624
rect 442994 156612 443000 156624
rect 443052 156612 443058 156664
rect 448422 156612 448428 156664
rect 448480 156652 448486 156664
rect 491662 156652 491668 156664
rect 448480 156624 491668 156652
rect 448480 156612 448486 156624
rect 491662 156612 491668 156624
rect 491720 156612 491726 156664
rect 491938 156612 491944 156664
rect 491996 156652 492002 156664
rect 556982 156652 556988 156664
rect 491996 156624 556988 156652
rect 491996 156612 492002 156624
rect 556982 156612 556988 156624
rect 557040 156612 557046 156664
rect 92014 156544 92020 156596
rect 92072 156584 92078 156596
rect 173437 156587 173495 156593
rect 173437 156584 173449 156587
rect 92072 156556 173449 156584
rect 92072 156544 92078 156556
rect 173437 156553 173449 156556
rect 173483 156553 173495 156587
rect 173437 156547 173495 156553
rect 173713 156587 173771 156593
rect 173713 156553 173725 156587
rect 173759 156584 173771 156587
rect 175734 156584 175740 156596
rect 173759 156556 175740 156584
rect 173759 156553 173771 156556
rect 173713 156547 173771 156553
rect 175734 156544 175740 156556
rect 175792 156544 175798 156596
rect 175921 156587 175979 156593
rect 175921 156553 175933 156587
rect 175967 156584 175979 156587
rect 225966 156584 225972 156596
rect 175967 156556 225972 156584
rect 175967 156553 175979 156556
rect 175921 156547 175979 156553
rect 225966 156544 225972 156556
rect 226024 156544 226030 156596
rect 420730 156544 420736 156596
rect 420788 156584 420794 156596
rect 450722 156584 450728 156596
rect 420788 156556 450728 156584
rect 420788 156544 420794 156556
rect 450722 156544 450728 156556
rect 450780 156544 450786 156596
rect 469858 156544 469864 156596
rect 469916 156584 469922 156596
rect 523862 156584 523868 156596
rect 469916 156556 523868 156584
rect 469916 156544 469922 156556
rect 523862 156544 523868 156556
rect 523920 156544 523926 156596
rect 99834 156476 99840 156528
rect 99892 156516 99898 156528
rect 186406 156516 186412 156528
rect 99892 156488 186412 156516
rect 99892 156476 99898 156488
rect 186406 156476 186412 156488
rect 186464 156476 186470 156528
rect 195149 156519 195207 156525
rect 195149 156485 195161 156519
rect 195195 156516 195207 156519
rect 196710 156516 196716 156528
rect 195195 156488 196716 156516
rect 195195 156485 195207 156488
rect 195149 156479 195207 156485
rect 196710 156476 196716 156488
rect 196768 156476 196774 156528
rect 197354 156476 197360 156528
rect 197412 156516 197418 156528
rect 204993 156519 205051 156525
rect 204993 156516 205005 156519
rect 197412 156488 205005 156516
rect 197412 156476 197418 156488
rect 204993 156485 205005 156488
rect 205039 156485 205051 156519
rect 204993 156479 205051 156485
rect 205082 156476 205088 156528
rect 205140 156516 205146 156528
rect 256694 156516 256700 156528
rect 205140 156488 256700 156516
rect 205140 156476 205146 156488
rect 256694 156476 256700 156488
rect 256752 156476 256758 156528
rect 467190 156476 467196 156528
rect 467248 156516 467254 156528
rect 519998 156516 520004 156528
rect 467248 156488 520004 156516
rect 467248 156476 467254 156488
rect 519998 156476 520004 156488
rect 520056 156476 520062 156528
rect 103790 156408 103796 156460
rect 103848 156448 103854 156460
rect 181993 156451 182051 156457
rect 181993 156448 182005 156451
rect 103848 156420 182005 156448
rect 103848 156408 103854 156420
rect 181993 156417 182005 156420
rect 182039 156417 182051 156451
rect 181993 156411 182051 156417
rect 182082 156408 182088 156460
rect 182140 156448 182146 156460
rect 182140 156420 185808 156448
rect 182140 156408 182146 156420
rect 105722 156340 105728 156392
rect 105780 156380 105786 156392
rect 185673 156383 185731 156389
rect 185673 156380 185685 156383
rect 105780 156352 185685 156380
rect 105780 156340 105786 156352
rect 185673 156349 185685 156352
rect 185719 156349 185731 156383
rect 185780 156380 185808 156420
rect 186314 156408 186320 156460
rect 186372 156448 186378 156460
rect 204901 156451 204959 156457
rect 186372 156420 200114 156448
rect 186372 156408 186378 156420
rect 195241 156383 195299 156389
rect 195241 156380 195253 156383
rect 185780 156352 195253 156380
rect 185673 156343 185731 156349
rect 195241 156349 195253 156352
rect 195287 156349 195299 156383
rect 195241 156343 195299 156349
rect 195333 156383 195391 156389
rect 195333 156349 195345 156383
rect 195379 156380 195391 156383
rect 199378 156380 199384 156392
rect 195379 156352 199384 156380
rect 195379 156349 195391 156352
rect 195333 156343 195391 156349
rect 199378 156340 199384 156352
rect 199436 156340 199442 156392
rect 200086 156380 200114 156420
rect 204901 156417 204913 156451
rect 204947 156448 204959 156451
rect 209866 156448 209872 156460
rect 204947 156420 209872 156448
rect 204947 156417 204959 156420
rect 204901 156411 204959 156417
rect 209866 156408 209872 156420
rect 209924 156408 209930 156460
rect 213733 156451 213791 156457
rect 213733 156417 213745 156451
rect 213779 156448 213791 156451
rect 217502 156448 217508 156460
rect 213779 156420 217508 156448
rect 213779 156417 213791 156420
rect 213733 156411 213791 156417
rect 217502 156408 217508 156420
rect 217560 156408 217566 156460
rect 220725 156451 220783 156457
rect 220725 156417 220737 156451
rect 220771 156448 220783 156451
rect 254578 156448 254584 156460
rect 220771 156420 254584 156448
rect 220771 156417 220783 156420
rect 220725 156411 220783 156417
rect 254578 156408 254584 156420
rect 254636 156408 254642 156460
rect 462682 156408 462688 156460
rect 462740 156448 462746 156460
rect 513098 156448 513104 156460
rect 462740 156420 513104 156448
rect 462740 156408 462746 156420
rect 513098 156408 513104 156420
rect 513156 156408 513162 156460
rect 239030 156380 239036 156392
rect 200086 156352 239036 156380
rect 239030 156340 239036 156352
rect 239088 156340 239094 156392
rect 456518 156340 456524 156392
rect 456576 156380 456582 156392
rect 504358 156380 504364 156392
rect 456576 156352 504364 156380
rect 456576 156340 456582 156352
rect 504358 156340 504364 156352
rect 504416 156340 504422 156392
rect 107654 156272 107660 156324
rect 107712 156312 107718 156324
rect 185397 156315 185455 156321
rect 185397 156312 185409 156315
rect 107712 156284 185409 156312
rect 107712 156272 107718 156284
rect 185397 156281 185409 156284
rect 185443 156281 185455 156315
rect 185397 156275 185455 156281
rect 185489 156315 185547 156321
rect 185489 156281 185501 156315
rect 185535 156312 185547 156315
rect 228542 156312 228548 156324
rect 185535 156284 228548 156312
rect 185535 156281 185547 156284
rect 185489 156275 185547 156281
rect 228542 156272 228548 156284
rect 228600 156272 228606 156324
rect 452562 156272 452568 156324
rect 452620 156312 452626 156324
rect 498562 156312 498568 156324
rect 452620 156284 498568 156312
rect 452620 156272 452626 156284
rect 498562 156272 498568 156284
rect 498620 156272 498626 156324
rect 115474 156204 115480 156256
rect 115532 156244 115538 156256
rect 195149 156247 195207 156253
rect 195149 156244 195161 156247
rect 115532 156216 195161 156244
rect 115532 156204 115538 156216
rect 195149 156213 195161 156216
rect 195195 156213 195207 156247
rect 195149 156207 195207 156213
rect 195241 156247 195299 156253
rect 195241 156213 195253 156247
rect 195287 156244 195299 156247
rect 233786 156244 233792 156256
rect 195287 156216 233792 156244
rect 195287 156213 195299 156216
rect 195241 156207 195299 156213
rect 233786 156204 233792 156216
rect 233844 156204 233850 156256
rect 449066 156204 449072 156256
rect 449124 156244 449130 156256
rect 492674 156244 492680 156256
rect 449124 156216 492680 156244
rect 449124 156204 449130 156216
rect 492674 156204 492680 156216
rect 492732 156204 492738 156256
rect 119338 156136 119344 156188
rect 119396 156176 119402 156188
rect 194873 156179 194931 156185
rect 194873 156176 194885 156179
rect 119396 156148 194885 156176
rect 119396 156136 119402 156148
rect 194873 156145 194885 156148
rect 194919 156145 194931 156179
rect 194873 156139 194931 156145
rect 194962 156136 194968 156188
rect 195020 156176 195026 156188
rect 204993 156179 205051 156185
rect 195020 156148 204944 156176
rect 195020 156136 195026 156148
rect 112530 156068 112536 156120
rect 112588 156108 112594 156120
rect 113269 156111 113327 156117
rect 113269 156108 113281 156111
rect 112588 156080 113281 156108
rect 112588 156068 112594 156080
rect 113269 156077 113281 156080
rect 113315 156077 113327 156111
rect 113269 156071 113327 156077
rect 128078 156068 128084 156120
rect 128136 156108 128142 156120
rect 204806 156108 204812 156120
rect 128136 156080 204812 156108
rect 128136 156068 128142 156080
rect 204806 156068 204812 156080
rect 204864 156068 204870 156120
rect 204916 156108 204944 156148
rect 204993 156145 205005 156179
rect 205039 156176 205051 156179
rect 247218 156176 247224 156188
rect 205039 156148 247224 156176
rect 205039 156145 205051 156148
rect 204993 156139 205051 156145
rect 247218 156136 247224 156148
rect 247276 156136 247282 156188
rect 453574 156136 453580 156188
rect 453632 156176 453638 156188
rect 499482 156176 499488 156188
rect 453632 156148 499488 156176
rect 453632 156136 453638 156148
rect 499482 156136 499488 156148
rect 499540 156136 499546 156188
rect 241606 156108 241612 156120
rect 204916 156080 241612 156108
rect 241606 156068 241612 156080
rect 241664 156068 241670 156120
rect 450354 156068 450360 156120
rect 450412 156108 450418 156120
rect 494606 156108 494612 156120
rect 450412 156080 494612 156108
rect 450412 156068 450418 156080
rect 494606 156068 494612 156080
rect 494664 156068 494670 156120
rect 96890 156000 96896 156052
rect 96948 156040 96954 156052
rect 155862 156040 155868 156052
rect 96948 156012 155868 156040
rect 96948 156000 96954 156012
rect 155862 156000 155868 156012
rect 155920 156000 155926 156052
rect 158714 156000 158720 156052
rect 158772 156040 158778 156052
rect 214285 156043 214343 156049
rect 158772 156012 214236 156040
rect 158772 156000 158778 156012
rect 128998 155972 129004 155984
rect 16546 155944 129004 155972
rect 14090 155864 14096 155916
rect 14148 155904 14154 155916
rect 16546 155904 16574 155944
rect 128998 155932 129004 155944
rect 129056 155932 129062 155984
rect 151740 155944 151860 155972
rect 14148 155876 16574 155904
rect 14148 155864 14154 155876
rect 44266 155864 44272 155916
rect 44324 155904 44330 155916
rect 140682 155904 140688 155916
rect 44324 155876 140688 155904
rect 44324 155864 44330 155876
rect 140682 155864 140688 155876
rect 140740 155864 140746 155916
rect 140774 155864 140780 155916
rect 140832 155904 140838 155916
rect 146941 155907 146999 155913
rect 146941 155904 146953 155907
rect 140832 155876 146953 155904
rect 140832 155864 140838 155876
rect 146941 155873 146953 155876
rect 146987 155873 146999 155907
rect 146941 155867 146999 155873
rect 149606 155864 149612 155916
rect 149664 155904 149670 155916
rect 151740 155904 151768 155944
rect 149664 155876 151768 155904
rect 151832 155904 151860 155944
rect 155402 155932 155408 155984
rect 155460 155972 155466 155984
rect 155460 155944 156552 155972
rect 155460 155932 155466 155944
rect 156417 155907 156475 155913
rect 156417 155904 156429 155907
rect 151832 155876 156429 155904
rect 149664 155864 149670 155876
rect 156417 155873 156429 155876
rect 156463 155873 156475 155907
rect 156524 155904 156552 155944
rect 156598 155932 156604 155984
rect 156656 155972 156662 155984
rect 214101 155975 214159 155981
rect 214101 155972 214113 155975
rect 156656 155944 214113 155972
rect 156656 155932 156662 155944
rect 214101 155941 214113 155944
rect 214147 155941 214159 155975
rect 214208 155972 214236 156012
rect 214285 156009 214297 156043
rect 214331 156040 214343 156043
rect 218146 156040 218152 156052
rect 214331 156012 218152 156040
rect 214331 156009 214343 156012
rect 214285 156003 214343 156009
rect 218146 156000 218152 156012
rect 218204 156000 218210 156052
rect 220630 156000 220636 156052
rect 220688 156040 220694 156052
rect 259822 156040 259828 156052
rect 220688 156012 259828 156040
rect 220688 156000 220694 156012
rect 259822 156000 259828 156012
rect 259880 156000 259886 156052
rect 286962 156040 286968 156052
rect 286923 156012 286968 156040
rect 286962 156000 286968 156012
rect 287020 156000 287026 156052
rect 302329 156043 302387 156049
rect 302329 156009 302341 156043
rect 302375 156040 302387 156043
rect 308125 156043 308183 156049
rect 308125 156040 308137 156043
rect 302375 156012 308137 156040
rect 302375 156009 302387 156012
rect 302329 156003 302387 156009
rect 308125 156009 308137 156012
rect 308171 156009 308183 156043
rect 308125 156003 308183 156009
rect 445110 156000 445116 156052
rect 445168 156040 445174 156052
rect 486786 156040 486792 156052
rect 445168 156012 486792 156040
rect 445168 156000 445174 156012
rect 486786 156000 486792 156012
rect 486844 156000 486850 156052
rect 220814 155972 220820 155984
rect 214208 155944 220820 155972
rect 214101 155935 214159 155941
rect 220814 155932 220820 155944
rect 220872 155932 220878 155984
rect 222102 155932 222108 155984
rect 222160 155972 222166 155984
rect 265066 155972 265072 155984
rect 222160 155944 265072 155972
rect 222160 155932 222166 155944
rect 265066 155932 265072 155944
rect 265124 155932 265130 155984
rect 287054 155972 287060 155984
rect 286888 155944 287060 155972
rect 158898 155904 158904 155916
rect 156524 155876 158904 155904
rect 156417 155867 156475 155873
rect 158898 155864 158904 155876
rect 158956 155864 158962 155916
rect 163222 155864 163228 155916
rect 163280 155904 163286 155916
rect 169849 155907 169907 155913
rect 169849 155904 169861 155907
rect 163280 155876 169861 155904
rect 163280 155864 163286 155876
rect 169849 155873 169861 155876
rect 169895 155873 169907 155907
rect 169849 155867 169907 155873
rect 172885 155907 172943 155913
rect 172885 155873 172897 155907
rect 172931 155904 172943 155907
rect 179414 155904 179420 155916
rect 172931 155876 179420 155904
rect 172931 155873 172943 155876
rect 172885 155867 172943 155873
rect 179414 155864 179420 155876
rect 179472 155864 179478 155916
rect 180794 155864 180800 155916
rect 180852 155904 180858 155916
rect 185673 155907 185731 155913
rect 185673 155904 185685 155907
rect 180852 155876 185685 155904
rect 180852 155864 180858 155876
rect 185673 155873 185685 155876
rect 185719 155873 185731 155907
rect 185673 155867 185731 155873
rect 186590 155864 186596 155916
rect 186648 155904 186654 155916
rect 190457 155907 190515 155913
rect 190457 155904 190469 155907
rect 186648 155876 190469 155904
rect 186648 155864 186654 155876
rect 190457 155873 190469 155876
rect 190503 155873 190515 155907
rect 190457 155867 190515 155873
rect 190546 155864 190552 155916
rect 190604 155904 190610 155916
rect 197354 155904 197360 155916
rect 190604 155876 197360 155904
rect 190604 155864 190610 155876
rect 197354 155864 197360 155876
rect 197412 155864 197418 155916
rect 197449 155907 197507 155913
rect 197449 155873 197461 155907
rect 197495 155904 197507 155907
rect 201954 155904 201960 155916
rect 197495 155876 201960 155904
rect 197495 155873 197507 155876
rect 197449 155867 197507 155873
rect 201954 155864 201960 155876
rect 202012 155864 202018 155916
rect 202049 155907 202107 155913
rect 202049 155873 202061 155907
rect 202095 155904 202107 155907
rect 204809 155907 204867 155913
rect 202095 155876 202920 155904
rect 202095 155873 202107 155876
rect 202049 155867 202107 155873
rect 5258 155796 5264 155848
rect 5316 155836 5322 155848
rect 102134 155836 102140 155848
rect 5316 155808 102140 155836
rect 5316 155796 5322 155808
rect 102134 155796 102140 155808
rect 102192 155796 102198 155848
rect 110598 155796 110604 155848
rect 110656 155836 110662 155848
rect 113174 155836 113180 155848
rect 110656 155808 113180 155836
rect 110656 155796 110662 155808
rect 113174 155796 113180 155808
rect 113232 155796 113238 155848
rect 113269 155839 113327 155845
rect 113269 155805 113281 155839
rect 113315 155836 113327 155839
rect 118053 155839 118111 155845
rect 118053 155836 118065 155839
rect 113315 155808 118065 155836
rect 113315 155805 113327 155808
rect 113269 155799 113327 155805
rect 118053 155805 118065 155808
rect 118099 155805 118111 155839
rect 118053 155799 118111 155805
rect 118326 155796 118332 155848
rect 118384 155836 118390 155848
rect 127529 155839 127587 155845
rect 127529 155836 127541 155839
rect 118384 155808 127541 155836
rect 118384 155796 118390 155808
rect 127529 155805 127541 155808
rect 127575 155805 127587 155839
rect 127529 155799 127587 155805
rect 127621 155839 127679 155845
rect 127621 155805 127633 155839
rect 127667 155836 127679 155839
rect 200022 155836 200028 155848
rect 127667 155808 200028 155836
rect 127667 155805 127679 155808
rect 127621 155799 127679 155805
rect 200022 155796 200028 155808
rect 200080 155796 200086 155848
rect 200206 155796 200212 155848
rect 200264 155836 200270 155848
rect 202782 155836 202788 155848
rect 200264 155808 202788 155836
rect 200264 155796 200270 155808
rect 202782 155796 202788 155808
rect 202840 155796 202846 155848
rect 202892 155836 202920 155876
rect 204809 155873 204821 155907
rect 204855 155904 204867 155907
rect 242069 155907 242127 155913
rect 242069 155904 242081 155907
rect 204855 155876 242081 155904
rect 204855 155873 204867 155876
rect 204809 155867 204867 155873
rect 242069 155873 242081 155876
rect 242115 155873 242127 155907
rect 242069 155867 242127 155873
rect 242158 155864 242164 155916
rect 242216 155904 242222 155916
rect 248969 155907 249027 155913
rect 248969 155904 248981 155907
rect 242216 155876 248981 155904
rect 242216 155864 242222 155876
rect 248969 155873 248981 155876
rect 249015 155873 249027 155907
rect 255406 155904 255412 155916
rect 248969 155867 249027 155873
rect 249076 155876 255412 155904
rect 208486 155836 208492 155848
rect 202892 155808 208492 155836
rect 208486 155796 208492 155808
rect 208544 155796 208550 155848
rect 213181 155839 213239 155845
rect 213181 155805 213193 155839
rect 213227 155836 213239 155839
rect 249076 155836 249104 155876
rect 255406 155864 255412 155876
rect 255464 155864 255470 155916
rect 257798 155864 257804 155916
rect 257856 155904 257862 155916
rect 262953 155907 263011 155913
rect 257856 155876 262904 155904
rect 257856 155864 257862 155876
rect 213227 155808 249104 155836
rect 213227 155805 213239 155808
rect 213181 155799 213239 155805
rect 252922 155796 252928 155848
rect 252980 155836 252986 155848
rect 262769 155839 262827 155845
rect 262769 155836 262781 155839
rect 252980 155808 262781 155836
rect 252980 155796 252986 155808
rect 262769 155805 262781 155808
rect 262815 155805 262827 155839
rect 262876 155836 262904 155876
rect 262953 155873 262965 155907
rect 262999 155904 263011 155907
rect 286888 155904 286916 155944
rect 287054 155932 287060 155944
rect 287112 155932 287118 155984
rect 296809 155975 296867 155981
rect 296548 155944 296714 155972
rect 262999 155876 286916 155904
rect 262999 155873 263011 155876
rect 262953 155867 263011 155873
rect 286962 155864 286968 155916
rect 287020 155904 287026 155916
rect 289817 155907 289875 155913
rect 289817 155904 289829 155907
rect 287020 155876 289829 155904
rect 287020 155864 287026 155876
rect 289817 155873 289829 155876
rect 289863 155873 289875 155907
rect 289817 155867 289875 155873
rect 289906 155864 289912 155916
rect 289964 155904 289970 155916
rect 296548 155904 296576 155944
rect 289964 155876 296576 155904
rect 296686 155904 296714 155944
rect 296809 155941 296821 155975
rect 296855 155972 296867 155975
rect 302513 155975 302571 155981
rect 302513 155972 302525 155975
rect 296855 155944 302525 155972
rect 296855 155941 296867 155944
rect 296809 155935 296867 155941
rect 302513 155941 302525 155944
rect 302559 155941 302571 155975
rect 302513 155935 302571 155941
rect 306837 155975 306895 155981
rect 306837 155941 306849 155975
rect 306883 155972 306895 155975
rect 412453 155975 412511 155981
rect 306883 155944 307156 155972
rect 306883 155941 306895 155944
rect 306837 155935 306895 155941
rect 307021 155907 307079 155913
rect 307021 155904 307033 155907
rect 296686 155876 307033 155904
rect 289964 155864 289970 155876
rect 307021 155873 307033 155876
rect 307067 155873 307079 155907
rect 307128 155904 307156 155944
rect 412453 155941 412465 155975
rect 412499 155972 412511 155975
rect 412499 155944 412772 155972
rect 412499 155941 412511 155944
rect 412453 155935 412511 155941
rect 309134 155904 309140 155916
rect 307128 155876 309140 155904
rect 307021 155867 307079 155873
rect 309134 155864 309140 155876
rect 309192 155864 309198 155916
rect 309410 155864 309416 155916
rect 309468 155904 309474 155916
rect 313369 155907 313427 155913
rect 313369 155904 313381 155907
rect 309468 155876 313381 155904
rect 309468 155864 309474 155876
rect 313369 155873 313381 155876
rect 313415 155873 313427 155907
rect 313369 155867 313427 155873
rect 315298 155864 315304 155916
rect 315356 155904 315362 155916
rect 329742 155904 329748 155916
rect 315356 155876 329748 155904
rect 315356 155864 315362 155876
rect 329742 155864 329748 155876
rect 329800 155864 329806 155916
rect 329926 155864 329932 155916
rect 329984 155904 329990 155916
rect 336458 155904 336464 155916
rect 329984 155876 336464 155904
rect 329984 155864 329990 155876
rect 336458 155864 336464 155876
rect 336516 155864 336522 155916
rect 338666 155864 338672 155916
rect 338724 155904 338730 155916
rect 344186 155904 344192 155916
rect 338724 155876 344192 155904
rect 338724 155864 338730 155876
rect 344186 155864 344192 155876
rect 344244 155864 344250 155916
rect 354214 155864 354220 155916
rect 354272 155904 354278 155916
rect 355962 155904 355968 155916
rect 354272 155876 355968 155904
rect 354272 155864 354278 155876
rect 355962 155864 355968 155876
rect 356020 155864 356026 155916
rect 388162 155864 388168 155916
rect 388220 155904 388226 155916
rect 393222 155904 393228 155916
rect 388220 155876 393228 155904
rect 388220 155864 388226 155876
rect 393222 155864 393228 155876
rect 393280 155864 393286 155916
rect 401686 155864 401692 155916
rect 401744 155904 401750 155916
rect 403986 155904 403992 155916
rect 401744 155876 403992 155904
rect 401744 155864 401750 155876
rect 403986 155864 403992 155876
rect 404044 155864 404050 155916
rect 404814 155864 404820 155916
rect 404872 155904 404878 155916
rect 407850 155904 407856 155916
rect 404872 155876 407856 155904
rect 404872 155864 404878 155876
rect 407850 155864 407856 155876
rect 407908 155864 407914 155916
rect 407945 155907 408003 155913
rect 407945 155873 407957 155907
rect 407991 155904 408003 155907
rect 407991 155876 412496 155904
rect 407991 155873 408003 155876
rect 407945 155867 408003 155873
rect 287885 155839 287943 155845
rect 287885 155836 287897 155839
rect 262876 155808 287897 155836
rect 262769 155799 262827 155805
rect 287885 155805 287897 155808
rect 287931 155805 287943 155839
rect 287885 155799 287943 155805
rect 287974 155796 287980 155848
rect 288032 155836 288038 155848
rect 293034 155836 293040 155848
rect 288032 155808 293040 155836
rect 288032 155796 288038 155808
rect 293034 155796 293040 155808
rect 293092 155796 293098 155848
rect 294782 155796 294788 155848
rect 294840 155836 294846 155848
rect 303249 155839 303307 155845
rect 294840 155808 303200 155836
rect 294840 155796 294846 155808
rect 55950 155728 55956 155780
rect 56008 155768 56014 155780
rect 153381 155771 153439 155777
rect 153381 155768 153393 155771
rect 56008 155740 153393 155768
rect 56008 155728 56014 155740
rect 153381 155737 153393 155740
rect 153427 155737 153439 155771
rect 153381 155731 153439 155737
rect 153470 155728 153476 155780
rect 153528 155768 153534 155780
rect 158809 155771 158867 155777
rect 158809 155768 158821 155771
rect 153528 155740 158821 155768
rect 153528 155728 153534 155740
rect 158809 155737 158821 155740
rect 158855 155737 158867 155771
rect 158809 155731 158867 155737
rect 159266 155728 159272 155780
rect 159324 155768 159330 155780
rect 169754 155768 169760 155780
rect 159324 155740 169760 155768
rect 159324 155728 159330 155740
rect 169754 155728 169760 155740
rect 169812 155728 169818 155780
rect 169849 155771 169907 155777
rect 169849 155737 169861 155771
rect 169895 155768 169907 155771
rect 173802 155768 173808 155780
rect 169895 155740 173808 155768
rect 169895 155737 169907 155740
rect 169849 155731 169907 155737
rect 173802 155728 173808 155740
rect 173860 155728 173866 155780
rect 175918 155728 175924 155780
rect 175976 155768 175982 155780
rect 229189 155771 229247 155777
rect 229189 155768 229201 155771
rect 175976 155740 229201 155768
rect 175976 155728 175982 155740
rect 229189 155737 229201 155740
rect 229235 155737 229247 155771
rect 235074 155768 235080 155780
rect 229189 155731 229247 155737
rect 229296 155740 235080 155768
rect 40402 155660 40408 155712
rect 40460 155700 40466 155712
rect 137097 155703 137155 155709
rect 137097 155700 137109 155703
rect 40460 155672 137109 155700
rect 40460 155660 40466 155672
rect 137097 155669 137109 155672
rect 137143 155669 137155 155703
rect 137097 155663 137155 155669
rect 137186 155660 137192 155712
rect 137244 155700 137250 155712
rect 172885 155703 172943 155709
rect 172885 155700 172897 155703
rect 137244 155672 172897 155700
rect 137244 155660 137250 155672
rect 172885 155669 172897 155672
rect 172931 155669 172943 155703
rect 172885 155663 172943 155669
rect 172974 155660 172980 155712
rect 173032 155700 173038 155712
rect 229296 155700 229324 155740
rect 235074 155728 235080 155740
rect 235132 155728 235138 155780
rect 241057 155771 241115 155777
rect 241057 155737 241069 155771
rect 241103 155768 241115 155771
rect 241103 155740 244274 155768
rect 241103 155737 241115 155740
rect 241057 155731 241115 155737
rect 173032 155672 229324 155700
rect 173032 155660 173038 155672
rect 229370 155660 229376 155712
rect 229428 155700 229434 155712
rect 233973 155703 234031 155709
rect 233973 155700 233985 155703
rect 229428 155672 233985 155700
rect 229428 155660 229434 155672
rect 233973 155669 233985 155672
rect 234019 155669 234031 155703
rect 233973 155663 234031 155669
rect 234065 155703 234123 155709
rect 234065 155669 234077 155703
rect 234111 155700 234123 155703
rect 237006 155700 237012 155712
rect 234111 155672 237012 155700
rect 234111 155669 234123 155672
rect 234065 155663 234123 155669
rect 237006 155660 237012 155672
rect 237064 155660 237070 155712
rect 237282 155660 237288 155712
rect 237340 155700 237346 155712
rect 243541 155703 243599 155709
rect 243541 155700 243553 155703
rect 237340 155672 243553 155700
rect 237340 155660 237346 155672
rect 243541 155669 243553 155672
rect 243587 155669 243599 155703
rect 244246 155700 244274 155740
rect 246022 155728 246028 155780
rect 246080 155768 246086 155780
rect 280706 155768 280712 155780
rect 246080 155740 280712 155768
rect 246080 155728 246086 155740
rect 280706 155728 280712 155740
rect 280764 155728 280770 155780
rect 281166 155728 281172 155780
rect 281224 155768 281230 155780
rect 286686 155768 286692 155780
rect 281224 155740 286692 155768
rect 281224 155728 281230 155740
rect 286686 155728 286692 155740
rect 286744 155728 286750 155780
rect 300581 155771 300639 155777
rect 300581 155768 300593 155771
rect 286796 155740 300593 155768
rect 246942 155700 246948 155712
rect 244246 155672 246948 155700
rect 243541 155663 243599 155669
rect 246942 155660 246948 155672
rect 247000 155660 247006 155712
rect 247034 155660 247040 155712
rect 247092 155700 247098 155712
rect 277581 155703 277639 155709
rect 247092 155672 277532 155700
rect 247092 155660 247098 155672
rect 31662 155592 31668 155644
rect 31720 155632 31726 155644
rect 117961 155635 118019 155641
rect 117961 155632 117973 155635
rect 31720 155604 117973 155632
rect 31720 155592 31726 155604
rect 117961 155601 117973 155604
rect 118007 155601 118019 155635
rect 117961 155595 118019 155601
rect 118053 155635 118111 155641
rect 118053 155601 118065 155635
rect 118099 155632 118111 155635
rect 156506 155632 156512 155644
rect 118099 155604 156512 155632
rect 118099 155601 118111 155604
rect 118053 155595 118111 155601
rect 156506 155592 156512 155604
rect 156564 155592 156570 155644
rect 160278 155592 160284 155644
rect 160336 155632 160342 155644
rect 221553 155635 221611 155641
rect 221553 155632 221565 155635
rect 160336 155604 221565 155632
rect 160336 155592 160342 155604
rect 221553 155601 221565 155604
rect 221599 155601 221611 155635
rect 221553 155595 221611 155601
rect 221645 155635 221703 155641
rect 221645 155601 221657 155635
rect 221691 155632 221703 155635
rect 224034 155632 224040 155644
rect 221691 155604 224040 155632
rect 221691 155601 221703 155604
rect 221645 155595 221703 155601
rect 224034 155592 224040 155604
rect 224092 155592 224098 155644
rect 224129 155635 224187 155641
rect 224129 155601 224141 155635
rect 224175 155632 224187 155635
rect 249058 155632 249064 155644
rect 224175 155604 249064 155632
rect 224175 155601 224187 155604
rect 224129 155595 224187 155601
rect 249058 155592 249064 155604
rect 249116 155592 249122 155644
rect 250898 155592 250904 155644
rect 250956 155632 250962 155644
rect 277394 155632 277400 155644
rect 250956 155604 277400 155632
rect 250956 155592 250962 155604
rect 277394 155592 277400 155604
rect 277452 155592 277458 155644
rect 277504 155632 277532 155672
rect 277581 155669 277593 155703
rect 277627 155700 277639 155703
rect 281997 155703 282055 155709
rect 281997 155700 282009 155703
rect 277627 155672 282009 155700
rect 277627 155669 277639 155672
rect 277581 155663 277639 155669
rect 281997 155669 282009 155672
rect 282043 155669 282055 155703
rect 281997 155663 282055 155669
rect 282086 155660 282092 155712
rect 282144 155700 282150 155712
rect 286796 155700 286824 155740
rect 300581 155737 300593 155740
rect 300627 155737 300639 155771
rect 300581 155731 300639 155737
rect 300670 155728 300676 155780
rect 300728 155768 300734 155780
rect 303172 155768 303200 155808
rect 303249 155805 303261 155839
rect 303295 155836 303307 155839
rect 316034 155836 316040 155848
rect 303295 155808 316040 155836
rect 303295 155805 303307 155808
rect 303249 155799 303307 155805
rect 316034 155796 316040 155808
rect 316092 155796 316098 155848
rect 320174 155796 320180 155848
rect 320232 155836 320238 155848
rect 320232 155808 328868 155836
rect 320232 155796 320238 155808
rect 307205 155771 307263 155777
rect 307205 155768 307217 155771
rect 300728 155740 302556 155768
rect 303172 155740 307217 155768
rect 300728 155728 300734 155740
rect 282144 155672 286824 155700
rect 286965 155703 287023 155709
rect 282144 155660 282150 155672
rect 286965 155669 286977 155703
rect 287011 155700 287023 155703
rect 302329 155703 302387 155709
rect 302329 155700 302341 155703
rect 287011 155672 302341 155700
rect 287011 155669 287023 155672
rect 286965 155663 287023 155669
rect 302329 155669 302341 155672
rect 302375 155669 302387 155703
rect 302528 155700 302556 155740
rect 307205 155737 307217 155740
rect 307251 155737 307263 155771
rect 307205 155731 307263 155737
rect 307294 155728 307300 155780
rect 307352 155768 307358 155780
rect 309226 155768 309232 155780
rect 307352 155740 309232 155768
rect 307352 155728 307358 155740
rect 309226 155728 309232 155740
rect 309284 155728 309290 155780
rect 312354 155728 312360 155780
rect 312412 155768 312418 155780
rect 326798 155768 326804 155780
rect 312412 155740 326804 155768
rect 312412 155728 312418 155740
rect 326798 155728 326804 155740
rect 326856 155728 326862 155780
rect 328840 155768 328868 155808
rect 328914 155796 328920 155848
rect 328972 155836 328978 155848
rect 334434 155836 334440 155848
rect 328972 155808 334440 155836
rect 328972 155796 328978 155808
rect 334434 155796 334440 155808
rect 334492 155796 334498 155848
rect 334802 155796 334808 155848
rect 334860 155836 334866 155848
rect 340782 155836 340788 155848
rect 334860 155808 340788 155836
rect 334860 155796 334866 155808
rect 340782 155796 340788 155808
rect 340840 155796 340846 155848
rect 353294 155796 353300 155848
rect 353352 155836 353358 155848
rect 355410 155836 355416 155848
rect 353352 155808 355416 155836
rect 353352 155796 353358 155808
rect 355410 155796 355416 155808
rect 355468 155796 355474 155848
rect 365070 155796 365076 155848
rect 365128 155836 365134 155848
rect 365990 155836 365996 155848
rect 365128 155808 365996 155836
rect 365128 155796 365134 155808
rect 365990 155796 365996 155808
rect 366048 155796 366054 155848
rect 403434 155796 403440 155848
rect 403492 155836 403498 155848
rect 406930 155836 406936 155848
rect 403492 155808 406936 155836
rect 403492 155796 403498 155808
rect 406930 155796 406936 155808
rect 406988 155796 406994 155848
rect 412468 155836 412496 155876
rect 412542 155864 412548 155916
rect 412600 155904 412606 155916
rect 412634 155904 412640 155916
rect 412600 155876 412640 155904
rect 412600 155864 412606 155876
rect 412634 155864 412640 155876
rect 412692 155864 412698 155916
rect 412744 155904 412772 155944
rect 506934 155932 506940 155984
rect 506992 155972 506998 155984
rect 506992 155944 572760 155972
rect 506992 155932 506998 155944
rect 428366 155904 428372 155916
rect 412744 155876 428372 155904
rect 428366 155864 428372 155876
rect 428424 155864 428430 155916
rect 430206 155864 430212 155916
rect 430264 155904 430270 155916
rect 464430 155904 464436 155916
rect 430264 155876 464436 155904
rect 430264 155864 430270 155876
rect 464430 155864 464436 155876
rect 464488 155864 464494 155916
rect 464982 155864 464988 155916
rect 465040 155904 465046 155916
rect 517054 155904 517060 155916
rect 465040 155876 517060 155904
rect 465040 155864 465046 155876
rect 517054 155864 517060 155876
rect 517112 155864 517118 155916
rect 572732 155904 572760 155944
rect 574554 155904 574560 155916
rect 572732 155876 574560 155904
rect 574554 155864 574560 155876
rect 574612 155864 574618 155916
rect 425422 155836 425428 155848
rect 412468 155808 425428 155836
rect 425422 155796 425428 155808
rect 425480 155796 425486 155848
rect 427630 155796 427636 155848
rect 427688 155836 427694 155848
rect 460474 155836 460480 155848
rect 427688 155808 460480 155836
rect 427688 155796 427694 155808
rect 460474 155796 460480 155808
rect 460532 155796 460538 155848
rect 467742 155796 467748 155848
rect 467800 155836 467806 155848
rect 520918 155836 520924 155848
rect 467800 155808 520924 155836
rect 467800 155796 467806 155808
rect 520918 155796 520924 155808
rect 520976 155796 520982 155848
rect 333238 155768 333244 155780
rect 328840 155740 333244 155768
rect 333238 155728 333244 155740
rect 333296 155728 333302 155780
rect 380894 155728 380900 155780
rect 380952 155768 380958 155780
rect 384482 155768 384488 155780
rect 380952 155740 384488 155768
rect 380952 155728 380958 155740
rect 384482 155728 384488 155740
rect 384540 155728 384546 155780
rect 412545 155771 412603 155777
rect 412545 155737 412557 155771
rect 412591 155768 412603 155771
rect 414658 155768 414664 155780
rect 412591 155740 414664 155768
rect 412591 155737 412603 155740
rect 412545 155731 412603 155737
rect 414658 155728 414664 155740
rect 414716 155728 414722 155780
rect 417329 155771 417387 155777
rect 417329 155737 417341 155771
rect 417375 155768 417387 155771
rect 429286 155768 429292 155780
rect 417375 155740 429292 155768
rect 417375 155737 417387 155740
rect 417329 155731 417387 155737
rect 429286 155728 429292 155740
rect 429344 155728 429350 155780
rect 430482 155728 430488 155780
rect 430540 155768 430546 155780
rect 465350 155768 465356 155780
rect 430540 155740 465356 155768
rect 430540 155728 430546 155740
rect 465350 155728 465356 155740
rect 465408 155728 465414 155780
rect 473078 155728 473084 155780
rect 473136 155768 473142 155780
rect 528738 155768 528744 155780
rect 473136 155740 528744 155768
rect 473136 155728 473142 155740
rect 528738 155728 528744 155740
rect 528796 155728 528802 155780
rect 306837 155703 306895 155709
rect 306837 155700 306849 155703
rect 302528 155672 306849 155700
rect 302329 155663 302387 155669
rect 306837 155669 306849 155672
rect 306883 155669 306895 155703
rect 306837 155663 306895 155669
rect 306929 155703 306987 155709
rect 306929 155669 306941 155703
rect 306975 155700 306987 155703
rect 313734 155700 313740 155712
rect 306975 155672 313740 155700
rect 306975 155669 306987 155672
rect 306929 155663 306987 155669
rect 313734 155660 313740 155672
rect 313792 155660 313798 155712
rect 314286 155660 314292 155712
rect 314344 155700 314350 155712
rect 328178 155700 328184 155712
rect 314344 155672 328184 155700
rect 314344 155660 314350 155672
rect 328178 155660 328184 155672
rect 328236 155660 328242 155712
rect 333790 155660 333796 155712
rect 333848 155700 333854 155712
rect 339402 155700 339408 155712
rect 333848 155672 339408 155700
rect 333848 155660 333854 155672
rect 339402 155660 339408 155672
rect 339460 155660 339466 155712
rect 342530 155660 342536 155712
rect 342588 155700 342594 155712
rect 348234 155700 348240 155712
rect 342588 155672 348240 155700
rect 342588 155660 342594 155672
rect 348234 155660 348240 155672
rect 348292 155660 348298 155712
rect 404170 155660 404176 155712
rect 404228 155700 404234 155712
rect 407945 155703 408003 155709
rect 407945 155700 407957 155703
rect 404228 155672 407957 155700
rect 404228 155660 404234 155672
rect 407945 155669 407957 155672
rect 407991 155669 408003 155703
rect 407945 155663 408003 155669
rect 409690 155660 409696 155712
rect 409748 155700 409754 155712
rect 434162 155700 434168 155712
rect 409748 155672 434168 155700
rect 409748 155660 409754 155672
rect 434162 155660 434168 155672
rect 434220 155660 434226 155712
rect 435358 155660 435364 155712
rect 435416 155700 435422 155712
rect 472158 155700 472164 155712
rect 435416 155672 472164 155700
rect 435416 155660 435422 155672
rect 472158 155660 472164 155672
rect 472216 155660 472222 155712
rect 478322 155660 478328 155712
rect 478380 155700 478386 155712
rect 536558 155700 536564 155712
rect 478380 155672 536564 155700
rect 478380 155660 478386 155672
rect 536558 155660 536564 155672
rect 536616 155660 536622 155712
rect 280065 155635 280123 155641
rect 280065 155632 280077 155635
rect 277504 155604 280077 155632
rect 280065 155601 280077 155604
rect 280111 155601 280123 155635
rect 280065 155595 280123 155601
rect 280154 155592 280160 155644
rect 280212 155632 280218 155644
rect 291746 155632 291752 155644
rect 280212 155604 291752 155632
rect 280212 155592 280218 155604
rect 291746 155592 291752 155604
rect 291804 155592 291810 155644
rect 291838 155592 291844 155644
rect 291896 155632 291902 155644
rect 302237 155635 302295 155641
rect 302237 155632 302249 155635
rect 291896 155604 302249 155632
rect 291896 155592 291902 155604
rect 302237 155601 302249 155604
rect 302283 155601 302295 155635
rect 302237 155595 302295 155601
rect 302513 155635 302571 155641
rect 302513 155601 302525 155635
rect 302559 155632 302571 155635
rect 304445 155635 304503 155641
rect 304445 155632 304457 155635
rect 302559 155604 304457 155632
rect 302559 155601 302571 155604
rect 302513 155595 302571 155601
rect 304445 155601 304457 155604
rect 304491 155601 304503 155635
rect 304445 155595 304503 155601
rect 304534 155592 304540 155644
rect 304592 155632 304598 155644
rect 311986 155632 311992 155644
rect 304592 155604 311992 155632
rect 304592 155592 304598 155604
rect 311986 155592 311992 155604
rect 312044 155592 312050 155644
rect 321646 155632 321652 155644
rect 313200 155604 321652 155632
rect 35526 155524 35532 155576
rect 35584 155564 35590 155576
rect 140774 155564 140780 155576
rect 35584 155536 140780 155564
rect 35584 155524 35590 155536
rect 140774 155524 140780 155536
rect 140832 155524 140838 155576
rect 141786 155524 141792 155576
rect 141844 155564 141850 155576
rect 143721 155567 143779 155573
rect 143721 155564 143733 155567
rect 141844 155536 143733 155564
rect 141844 155524 141850 155536
rect 143721 155533 143733 155536
rect 143767 155533 143779 155567
rect 143721 155527 143779 155533
rect 143810 155524 143816 155576
rect 143868 155564 143874 155576
rect 153102 155564 153108 155576
rect 143868 155536 153108 155564
rect 143868 155524 143874 155536
rect 153102 155524 153108 155536
rect 153160 155524 153166 155576
rect 153381 155567 153439 155573
rect 153381 155533 153393 155567
rect 153427 155564 153439 155567
rect 155310 155564 155316 155576
rect 153427 155536 155316 155564
rect 153427 155533 153439 155536
rect 153381 155527 153439 155533
rect 155310 155524 155316 155536
rect 155368 155524 155374 155576
rect 156141 155567 156199 155573
rect 156141 155533 156153 155567
rect 156187 155564 156199 155567
rect 162762 155564 162768 155576
rect 156187 155536 162768 155564
rect 156187 155533 156199 155536
rect 156141 155527 156199 155533
rect 162762 155524 162768 155536
rect 162820 155524 162826 155576
rect 164142 155524 164148 155576
rect 164200 155564 164206 155576
rect 224221 155567 224279 155573
rect 224221 155564 224233 155567
rect 164200 155536 224233 155564
rect 164200 155524 164206 155536
rect 224221 155533 224233 155536
rect 224267 155533 224279 155567
rect 224221 155527 224279 155533
rect 225598 155524 225604 155576
rect 225656 155564 225662 155576
rect 229370 155564 229376 155576
rect 225656 155536 229376 155564
rect 225656 155524 225662 155536
rect 229370 155524 229376 155536
rect 229428 155524 229434 155576
rect 229462 155524 229468 155576
rect 229520 155564 229526 155576
rect 264974 155564 264980 155576
rect 229520 155536 264980 155564
rect 229520 155524 229526 155536
rect 264974 155524 264980 155536
rect 265032 155524 265038 155576
rect 266538 155524 266544 155576
rect 266596 155564 266602 155576
rect 287793 155567 287851 155573
rect 287793 155564 287805 155567
rect 266596 155536 287805 155564
rect 266596 155524 266602 155536
rect 287793 155533 287805 155536
rect 287839 155533 287851 155567
rect 287793 155527 287851 155533
rect 287885 155567 287943 155573
rect 287885 155533 287897 155567
rect 287931 155564 287943 155567
rect 288897 155567 288955 155573
rect 288897 155564 288909 155567
rect 287931 155536 288909 155564
rect 287931 155533 287943 155536
rect 287885 155527 287943 155533
rect 288897 155533 288909 155536
rect 288943 155533 288955 155567
rect 288897 155527 288955 155533
rect 288986 155524 288992 155576
rect 289044 155564 289050 155576
rect 292853 155567 292911 155573
rect 292853 155564 292865 155567
rect 289044 155536 292865 155564
rect 289044 155524 289050 155536
rect 292853 155533 292865 155536
rect 292899 155533 292911 155567
rect 292853 155527 292911 155533
rect 293862 155524 293868 155576
rect 293920 155564 293926 155576
rect 303249 155567 303307 155573
rect 303249 155564 303261 155567
rect 293920 155536 303261 155564
rect 293920 155524 293926 155536
rect 303249 155533 303261 155536
rect 303295 155533 303307 155567
rect 306926 155564 306932 155576
rect 303249 155527 303307 155533
rect 303356 155536 306932 155564
rect 29638 155456 29644 155508
rect 29696 155496 29702 155508
rect 31662 155496 31668 155508
rect 29696 155468 31668 155496
rect 29696 155456 29702 155468
rect 31662 155456 31668 155468
rect 31720 155456 31726 155508
rect 32582 155456 32588 155508
rect 32640 155496 32646 155508
rect 132770 155496 132776 155508
rect 32640 155468 132776 155496
rect 32640 155456 32646 155468
rect 132770 155456 132776 155468
rect 132828 155456 132834 155508
rect 133877 155499 133935 155505
rect 133877 155496 133889 155499
rect 132880 155468 133889 155496
rect 12158 155388 12164 155440
rect 12216 155428 12222 155440
rect 25498 155428 25504 155440
rect 12216 155400 25504 155428
rect 12216 155388 12222 155400
rect 25498 155388 25504 155400
rect 25556 155388 25562 155440
rect 27706 155388 27712 155440
rect 27764 155428 27770 155440
rect 132880 155428 132908 155468
rect 133877 155465 133889 155468
rect 133923 155465 133935 155499
rect 133877 155459 133935 155465
rect 133966 155456 133972 155508
rect 134024 155496 134030 155508
rect 138017 155499 138075 155505
rect 138017 155496 138029 155499
rect 134024 155468 138029 155496
rect 134024 155456 134030 155468
rect 138017 155465 138029 155468
rect 138063 155465 138075 155499
rect 138017 155459 138075 155465
rect 139854 155456 139860 155508
rect 139912 155496 139918 155508
rect 139912 155468 145604 155496
rect 139912 155456 139918 155468
rect 27764 155400 132908 155428
rect 27764 155388 27770 155400
rect 132954 155388 132960 155440
rect 133012 155428 133018 155440
rect 137097 155431 137155 155437
rect 133012 155400 137048 155428
rect 133012 155388 133018 155400
rect 23842 155320 23848 155372
rect 23900 155360 23906 155372
rect 23900 155332 124996 155360
rect 23900 155320 23906 155332
rect 9214 155252 9220 155304
rect 9272 155292 9278 155304
rect 117869 155295 117927 155301
rect 117869 155292 117881 155295
rect 9272 155264 117881 155292
rect 9272 155252 9278 155264
rect 117869 155261 117881 155264
rect 117915 155261 117927 155295
rect 117869 155255 117927 155261
rect 117961 155295 118019 155301
rect 117961 155261 117973 155295
rect 118007 155292 118019 155295
rect 124968 155292 124996 155332
rect 125226 155320 125232 155372
rect 125284 155360 125290 155372
rect 128817 155363 128875 155369
rect 128817 155360 128829 155363
rect 125284 155332 128829 155360
rect 125284 155320 125290 155332
rect 128817 155329 128829 155332
rect 128863 155329 128875 155363
rect 128817 155323 128875 155329
rect 130102 155320 130108 155372
rect 130160 155360 130166 155372
rect 133877 155363 133935 155369
rect 130160 155332 133092 155360
rect 130160 155320 130166 155332
rect 132954 155292 132960 155304
rect 118007 155264 124904 155292
rect 124968 155264 132960 155292
rect 118007 155261 118019 155264
rect 117961 155255 118019 155261
rect 4338 155184 4344 155236
rect 4396 155224 4402 155236
rect 11514 155224 11520 155236
rect 4396 155196 11520 155224
rect 4396 155184 4402 155196
rect 11514 155184 11520 155196
rect 11572 155184 11578 155236
rect 16022 155184 16028 155236
rect 16080 155224 16086 155236
rect 124769 155227 124827 155233
rect 124769 155224 124781 155227
rect 16080 155196 124781 155224
rect 16080 155184 16086 155196
rect 124769 155193 124781 155196
rect 124815 155193 124827 155227
rect 124876 155224 124904 155264
rect 132954 155252 132960 155264
rect 133012 155252 133018 155304
rect 132865 155227 132923 155233
rect 132865 155224 132877 155227
rect 124876 155196 132877 155224
rect 124769 155187 124827 155193
rect 132865 155193 132877 155196
rect 132911 155193 132923 155227
rect 133064 155224 133092 155332
rect 133877 155329 133889 155363
rect 133923 155360 133935 155363
rect 136542 155360 136548 155372
rect 133923 155332 136548 155360
rect 133923 155329 133935 155332
rect 133877 155323 133935 155329
rect 136542 155320 136548 155332
rect 136600 155320 136606 155372
rect 137020 155360 137048 155400
rect 137097 155397 137109 155431
rect 137143 155428 137155 155431
rect 143626 155428 143632 155440
rect 137143 155400 143632 155428
rect 137143 155397 137155 155400
rect 137097 155391 137155 155397
rect 143626 155388 143632 155400
rect 143684 155388 143690 155440
rect 143721 155431 143779 155437
rect 143721 155397 143733 155431
rect 143767 155428 143779 155431
rect 145377 155431 145435 155437
rect 145377 155428 145389 155431
rect 143767 155400 145389 155428
rect 143767 155397 143779 155400
rect 143721 155391 143779 155397
rect 145377 155397 145389 155400
rect 145423 155397 145435 155431
rect 145377 155391 145435 155397
rect 137189 155363 137247 155369
rect 137189 155360 137201 155363
rect 137020 155332 137201 155360
rect 137189 155329 137201 155332
rect 137235 155329 137247 155363
rect 144822 155360 144828 155372
rect 137189 155323 137247 155329
rect 137296 155332 144828 155360
rect 133141 155295 133199 155301
rect 133141 155261 133153 155295
rect 133187 155292 133199 155295
rect 135162 155292 135168 155304
rect 133187 155264 135168 155292
rect 133187 155261 133199 155264
rect 133141 155255 133199 155261
rect 135162 155252 135168 155264
rect 135220 155252 135226 155304
rect 137097 155227 137155 155233
rect 137097 155224 137109 155227
rect 133064 155196 137109 155224
rect 132865 155187 132923 155193
rect 137097 155193 137109 155196
rect 137143 155193 137155 155227
rect 137097 155187 137155 155193
rect 52086 155116 52092 155168
rect 52144 155156 52150 155168
rect 137296 155156 137324 155332
rect 144822 155320 144828 155332
rect 144880 155320 144886 155372
rect 145576 155360 145604 155468
rect 145650 155456 145656 155508
rect 145708 155496 145714 155508
rect 147125 155499 147183 155505
rect 147125 155496 147137 155499
rect 145708 155468 147137 155496
rect 145708 155456 145714 155468
rect 147125 155465 147137 155468
rect 147171 155465 147183 155499
rect 147125 155459 147183 155465
rect 147582 155456 147588 155508
rect 147640 155496 147646 155508
rect 156598 155496 156604 155508
rect 147640 155468 156604 155496
rect 147640 155456 147646 155468
rect 156598 155456 156604 155468
rect 156656 155456 156662 155508
rect 156690 155456 156696 155508
rect 156748 155496 156754 155508
rect 221645 155499 221703 155505
rect 221645 155496 221657 155499
rect 156748 155468 221657 155496
rect 156748 155456 156754 155468
rect 221645 155465 221657 155468
rect 221691 155465 221703 155499
rect 221645 155459 221703 155465
rect 221734 155456 221740 155508
rect 221792 155496 221798 155508
rect 248877 155499 248935 155505
rect 248877 155496 248889 155499
rect 221792 155468 248889 155496
rect 221792 155456 221798 155468
rect 248877 155465 248889 155468
rect 248923 155465 248935 155499
rect 248877 155459 248935 155465
rect 248969 155499 249027 155505
rect 248969 155465 248981 155499
rect 249015 155496 249027 155499
rect 281534 155496 281540 155508
rect 249015 155468 281540 155496
rect 249015 155465 249027 155468
rect 248969 155459 249027 155465
rect 281534 155456 281540 155468
rect 281592 155456 281598 155508
rect 281997 155499 282055 155505
rect 281997 155465 282009 155499
rect 282043 155496 282055 155499
rect 284018 155496 284024 155508
rect 282043 155468 284024 155496
rect 282043 155465 282055 155468
rect 281997 155459 282055 155465
rect 284018 155456 284024 155468
rect 284076 155456 284082 155508
rect 284110 155456 284116 155508
rect 284168 155496 284174 155508
rect 303356 155496 303384 155536
rect 306926 155524 306932 155536
rect 306984 155524 306990 155576
rect 307021 155567 307079 155573
rect 307021 155533 307033 155567
rect 307067 155564 307079 155567
rect 313090 155564 313096 155576
rect 307067 155536 313096 155564
rect 307067 155533 307079 155536
rect 307021 155527 307079 155533
rect 313090 155524 313096 155536
rect 313148 155524 313154 155576
rect 284168 155468 303384 155496
rect 303433 155499 303491 155505
rect 284168 155456 284174 155468
rect 303433 155465 303445 155499
rect 303479 155496 303491 155499
rect 308030 155496 308036 155508
rect 303479 155468 308036 155496
rect 303479 155465 303491 155468
rect 303433 155459 303491 155465
rect 308030 155456 308036 155468
rect 308088 155456 308094 155508
rect 308125 155499 308183 155505
rect 308125 155465 308137 155499
rect 308171 155496 308183 155499
rect 308171 155468 310376 155496
rect 308171 155465 308183 155468
rect 308125 155459 308183 155465
rect 145745 155431 145803 155437
rect 145745 155397 145757 155431
rect 145791 155428 145803 155431
rect 202049 155431 202107 155437
rect 202049 155428 202061 155431
rect 145791 155400 202061 155428
rect 145791 155397 145803 155400
rect 145745 155391 145803 155397
rect 202049 155397 202061 155400
rect 202095 155397 202107 155431
rect 202049 155391 202107 155397
rect 202141 155431 202199 155437
rect 202141 155397 202153 155431
rect 202187 155428 202199 155431
rect 206462 155428 206468 155440
rect 202187 155400 206468 155428
rect 202187 155397 202199 155400
rect 202141 155391 202199 155397
rect 206462 155388 206468 155400
rect 206520 155388 206526 155440
rect 209869 155431 209927 155437
rect 209869 155397 209881 155431
rect 209915 155428 209927 155431
rect 211890 155428 211896 155440
rect 209915 155400 211896 155428
rect 209915 155397 209927 155400
rect 209869 155391 209927 155397
rect 211890 155388 211896 155400
rect 211948 155388 211954 155440
rect 211982 155388 211988 155440
rect 212040 155428 212046 155440
rect 212040 155400 215708 155428
rect 212040 155388 212046 155400
rect 146478 155360 146484 155372
rect 145576 155332 146484 155360
rect 146478 155320 146484 155332
rect 146536 155320 146542 155372
rect 146849 155363 146907 155369
rect 146849 155329 146861 155363
rect 146895 155360 146907 155363
rect 149054 155360 149060 155372
rect 146895 155332 149060 155360
rect 146895 155329 146907 155332
rect 146849 155323 146907 155329
rect 149054 155320 149060 155332
rect 149112 155320 149118 155372
rect 151538 155320 151544 155372
rect 151596 155360 151602 155372
rect 158714 155360 158720 155372
rect 151596 155332 158720 155360
rect 151596 155320 151602 155332
rect 158714 155320 158720 155332
rect 158772 155320 158778 155372
rect 158809 155363 158867 155369
rect 158809 155329 158821 155363
rect 158855 155360 158867 155363
rect 214653 155363 214711 155369
rect 214653 155360 214665 155363
rect 158855 155332 214665 155360
rect 158855 155329 158867 155332
rect 158809 155323 158867 155329
rect 214653 155329 214665 155332
rect 214699 155329 214711 155363
rect 215680 155360 215708 155400
rect 217778 155388 217784 155440
rect 217836 155428 217842 155440
rect 222102 155428 222108 155440
rect 217836 155400 222108 155428
rect 217836 155388 217842 155400
rect 222102 155388 222108 155400
rect 222160 155388 222166 155440
rect 223577 155431 223635 155437
rect 223577 155397 223589 155431
rect 223623 155428 223635 155431
rect 226518 155428 226524 155440
rect 223623 155400 226524 155428
rect 223623 155397 223635 155400
rect 223577 155391 223635 155397
rect 226518 155388 226524 155400
rect 226576 155388 226582 155440
rect 226610 155388 226616 155440
rect 226668 155428 226674 155440
rect 269390 155428 269396 155440
rect 226668 155400 269396 155428
rect 226668 155388 226674 155400
rect 269390 155388 269396 155400
rect 269448 155388 269454 155440
rect 269482 155388 269488 155440
rect 269540 155428 269546 155440
rect 269540 155400 277394 155428
rect 269540 155388 269546 155400
rect 224129 155363 224187 155369
rect 224129 155360 224141 155363
rect 215680 155332 224141 155360
rect 214653 155323 214711 155329
rect 224129 155329 224141 155332
rect 224175 155329 224187 155363
rect 224129 155323 224187 155329
rect 224221 155363 224279 155369
rect 224221 155329 224233 155363
rect 224267 155360 224279 155363
rect 229278 155360 229284 155372
rect 224267 155332 229284 155360
rect 224267 155329 224279 155332
rect 224221 155323 224279 155329
rect 229278 155320 229284 155332
rect 229336 155320 229342 155372
rect 229373 155363 229431 155369
rect 229373 155329 229385 155363
rect 229419 155360 229431 155363
rect 233789 155363 233847 155369
rect 233789 155360 233801 155363
rect 229419 155332 233801 155360
rect 229419 155329 229431 155332
rect 229373 155323 229431 155329
rect 233789 155329 233801 155332
rect 233835 155329 233847 155363
rect 233789 155323 233847 155329
rect 233881 155363 233939 155369
rect 233881 155329 233893 155363
rect 233927 155360 233939 155363
rect 258629 155363 258687 155369
rect 258629 155360 258641 155363
rect 233927 155332 258641 155360
rect 233927 155329 233939 155332
rect 233881 155323 233939 155329
rect 258629 155329 258641 155332
rect 258675 155329 258687 155363
rect 258629 155323 258687 155329
rect 258718 155320 258724 155372
rect 258776 155360 258782 155372
rect 260558 155360 260564 155372
rect 258776 155332 260564 155360
rect 258776 155320 258782 155332
rect 260558 155320 260564 155332
rect 260616 155320 260622 155372
rect 260650 155320 260656 155372
rect 260708 155360 260714 155372
rect 264149 155363 264207 155369
rect 264149 155360 264161 155363
rect 260708 155332 264161 155360
rect 260708 155320 260714 155332
rect 264149 155329 264161 155332
rect 264195 155329 264207 155363
rect 264149 155323 264207 155329
rect 265526 155320 265532 155372
rect 265584 155360 265590 155372
rect 272705 155363 272763 155369
rect 272705 155360 272717 155363
rect 265584 155332 272717 155360
rect 265584 155320 265590 155332
rect 272705 155329 272717 155332
rect 272751 155329 272763 155363
rect 272705 155323 272763 155329
rect 272794 155320 272800 155372
rect 272852 155360 272858 155372
rect 277118 155360 277124 155372
rect 272852 155332 277124 155360
rect 272852 155320 272858 155332
rect 277118 155320 277124 155332
rect 277176 155320 277182 155372
rect 277366 155360 277394 155400
rect 277486 155388 277492 155440
rect 277544 155428 277550 155440
rect 279142 155428 279148 155440
rect 277544 155400 279148 155428
rect 277544 155388 277550 155400
rect 279142 155388 279148 155400
rect 279200 155388 279206 155440
rect 279234 155388 279240 155440
rect 279292 155428 279298 155440
rect 296717 155431 296775 155437
rect 296717 155428 296729 155431
rect 279292 155400 296729 155428
rect 279292 155388 279298 155400
rect 296717 155397 296729 155400
rect 296763 155397 296775 155431
rect 296717 155391 296775 155397
rect 296809 155431 296867 155437
rect 296809 155397 296821 155431
rect 296855 155428 296867 155431
rect 298649 155431 298707 155437
rect 298649 155428 298661 155431
rect 296855 155400 298661 155428
rect 296855 155397 296867 155400
rect 296809 155391 296867 155397
rect 298649 155397 298661 155400
rect 298695 155397 298707 155431
rect 298649 155391 298707 155397
rect 298738 155388 298744 155440
rect 298796 155428 298802 155440
rect 302513 155431 302571 155437
rect 298796 155400 302234 155428
rect 298796 155388 298802 155400
rect 288713 155363 288771 155369
rect 288713 155360 288725 155363
rect 277366 155332 288725 155360
rect 288713 155329 288725 155332
rect 288759 155329 288771 155363
rect 288713 155323 288771 155329
rect 288897 155363 288955 155369
rect 288897 155329 288909 155363
rect 288943 155360 288955 155363
rect 289998 155360 290004 155372
rect 288943 155332 290004 155360
rect 288943 155329 288955 155332
rect 288897 155323 288955 155329
rect 289998 155320 290004 155332
rect 290056 155320 290062 155372
rect 290918 155320 290924 155372
rect 290976 155360 290982 155372
rect 301317 155363 301375 155369
rect 301317 155360 301329 155363
rect 290976 155332 301329 155360
rect 290976 155320 290982 155332
rect 301317 155329 301329 155332
rect 301363 155329 301375 155363
rect 302206 155360 302234 155400
rect 302513 155397 302525 155431
rect 302559 155428 302571 155431
rect 308582 155428 308588 155440
rect 302559 155400 308588 155428
rect 302559 155397 302571 155400
rect 302513 155391 302571 155397
rect 308582 155388 308588 155400
rect 308640 155388 308646 155440
rect 310348 155428 310376 155468
rect 310422 155456 310428 155508
rect 310480 155496 310486 155508
rect 313200 155496 313228 155604
rect 321646 155592 321652 155604
rect 321704 155592 321710 155644
rect 322106 155592 322112 155644
rect 322164 155632 322170 155644
rect 334618 155632 334624 155644
rect 322164 155604 334624 155632
rect 322164 155592 322170 155604
rect 334618 155592 334624 155604
rect 334676 155592 334682 155644
rect 337654 155592 337660 155644
rect 337712 155632 337718 155644
rect 342714 155632 342720 155644
rect 337712 155604 342720 155632
rect 337712 155592 337718 155604
rect 342714 155592 342720 155604
rect 342772 155592 342778 155644
rect 344554 155592 344560 155644
rect 344612 155632 344618 155644
rect 349522 155632 349528 155644
rect 344612 155604 349528 155632
rect 344612 155592 344618 155604
rect 349522 155592 349528 155604
rect 349580 155592 349586 155644
rect 385862 155592 385868 155644
rect 385920 155632 385926 155644
rect 389358 155632 389364 155644
rect 385920 155604 389364 155632
rect 385920 155592 385926 155604
rect 389358 155592 389364 155604
rect 389416 155592 389422 155644
rect 406102 155592 406108 155644
rect 406160 155632 406166 155644
rect 412453 155635 412511 155641
rect 412453 155632 412465 155635
rect 406160 155604 412465 155632
rect 406160 155592 406166 155604
rect 412453 155601 412465 155604
rect 412499 155601 412511 155635
rect 437106 155632 437112 155644
rect 412453 155595 412511 155601
rect 412606 155604 437112 155632
rect 313369 155567 313427 155573
rect 313369 155533 313381 155567
rect 313415 155564 313427 155567
rect 319073 155567 319131 155573
rect 319073 155564 319085 155567
rect 313415 155536 319085 155564
rect 313415 155533 313427 155536
rect 313369 155527 313427 155533
rect 319073 155533 319085 155536
rect 319119 155533 319131 155567
rect 319073 155527 319131 155533
rect 319162 155524 319168 155576
rect 319220 155564 319226 155576
rect 332594 155564 332600 155576
rect 319220 155536 332600 155564
rect 319220 155524 319226 155536
rect 332594 155524 332600 155536
rect 332652 155524 332658 155576
rect 335722 155524 335728 155576
rect 335780 155564 335786 155576
rect 340966 155564 340972 155576
rect 335780 155536 340972 155564
rect 335780 155524 335786 155536
rect 340966 155524 340972 155536
rect 341024 155524 341030 155576
rect 358170 155524 358176 155576
rect 358228 155564 358234 155576
rect 358814 155564 358820 155576
rect 358228 155536 358820 155564
rect 358228 155524 358234 155536
rect 358814 155524 358820 155536
rect 358872 155524 358878 155576
rect 379606 155524 379612 155576
rect 379664 155564 379670 155576
rect 382550 155564 382556 155576
rect 379664 155536 382556 155564
rect 379664 155524 379670 155536
rect 382550 155524 382556 155536
rect 382608 155524 382614 155576
rect 385954 155524 385960 155576
rect 386012 155564 386018 155576
rect 390278 155564 390284 155576
rect 386012 155536 390284 155564
rect 386012 155524 386018 155536
rect 390278 155524 390284 155536
rect 390336 155524 390342 155576
rect 411990 155524 411996 155576
rect 412048 155564 412054 155576
rect 412606 155564 412634 155604
rect 437106 155592 437112 155604
rect 437164 155592 437170 155644
rect 438670 155592 438676 155644
rect 438728 155632 438734 155644
rect 477034 155632 477040 155644
rect 438728 155604 477040 155632
rect 438728 155592 438734 155604
rect 477034 155592 477040 155604
rect 477092 155592 477098 155644
rect 479610 155592 479616 155644
rect 479668 155632 479674 155644
rect 538490 155632 538496 155644
rect 479668 155604 538496 155632
rect 479668 155592 479674 155604
rect 538490 155592 538496 155604
rect 538548 155592 538554 155644
rect 412048 155536 412634 155564
rect 412048 155524 412054 155536
rect 413830 155524 413836 155576
rect 413888 155564 413894 155576
rect 416682 155564 416688 155576
rect 413888 155536 416688 155564
rect 413888 155524 413894 155536
rect 416682 155524 416688 155536
rect 416740 155524 416746 155576
rect 417421 155567 417479 155573
rect 417421 155533 417433 155567
rect 417467 155564 417479 155567
rect 430298 155564 430304 155576
rect 417467 155536 430304 155564
rect 417467 155533 417479 155536
rect 417421 155527 417479 155533
rect 430298 155524 430304 155536
rect 430356 155524 430362 155576
rect 433058 155524 433064 155576
rect 433116 155564 433122 155576
rect 469306 155564 469312 155576
rect 433116 155536 469312 155564
rect 433116 155524 433122 155536
rect 469306 155524 469312 155536
rect 469364 155524 469370 155576
rect 482186 155524 482192 155576
rect 482244 155564 482250 155576
rect 542354 155564 542360 155576
rect 482244 155536 542360 155564
rect 482244 155524 482250 155536
rect 542354 155524 542360 155536
rect 542412 155524 542418 155576
rect 575474 155524 575480 155576
rect 575532 155564 575538 155576
rect 576486 155564 576492 155576
rect 575532 155536 576492 155564
rect 575532 155524 575538 155536
rect 576486 155524 576492 155536
rect 576544 155524 576550 155576
rect 578237 155567 578295 155573
rect 578237 155533 578249 155567
rect 578283 155564 578295 155567
rect 578418 155564 578424 155576
rect 578283 155536 578424 155564
rect 578283 155533 578295 155536
rect 578237 155527 578295 155533
rect 578418 155524 578424 155536
rect 578476 155524 578482 155576
rect 310480 155468 313228 155496
rect 310480 155456 310486 155468
rect 313274 155456 313280 155508
rect 313332 155496 313338 155508
rect 328362 155496 328368 155508
rect 313332 155468 328368 155496
rect 313332 155456 313338 155468
rect 328362 155456 328368 155468
rect 328420 155456 328426 155508
rect 330846 155456 330852 155508
rect 330904 155496 330910 155508
rect 336550 155496 336556 155508
rect 330904 155468 336556 155496
rect 330904 155456 330910 155468
rect 336550 155456 336556 155468
rect 336608 155456 336614 155508
rect 378134 155456 378140 155508
rect 378192 155496 378198 155508
rect 380618 155496 380624 155508
rect 378192 155468 380624 155496
rect 378192 155456 378198 155468
rect 380618 155456 380624 155468
rect 380676 155456 380682 155508
rect 382366 155456 382372 155508
rect 382424 155496 382430 155508
rect 385494 155496 385500 155508
rect 382424 155468 385500 155496
rect 382424 155456 382430 155468
rect 385494 155456 385500 155468
rect 385552 155456 385558 155508
rect 386782 155456 386788 155508
rect 386840 155496 386846 155508
rect 391290 155496 391296 155508
rect 386840 155468 391296 155496
rect 386840 155456 386846 155468
rect 391290 155456 391296 155468
rect 391348 155456 391354 155508
rect 404262 155456 404268 155508
rect 404320 155496 404326 155508
rect 405918 155496 405924 155508
rect 404320 155468 405924 155496
rect 404320 155456 404326 155468
rect 405918 155456 405924 155468
rect 405976 155456 405982 155508
rect 407758 155456 407764 155508
rect 407816 155496 407822 155508
rect 412361 155499 412419 155505
rect 412361 155496 412373 155499
rect 407816 155468 412373 155496
rect 407816 155456 407822 155468
rect 412361 155465 412373 155468
rect 412407 155465 412419 155499
rect 412361 155459 412419 155465
rect 412450 155456 412456 155508
rect 412508 155496 412514 155508
rect 438118 155496 438124 155508
rect 412508 155468 438124 155496
rect 412508 155456 412514 155468
rect 438118 155456 438124 155468
rect 438176 155456 438182 155508
rect 476114 155496 476120 155508
rect 438228 155468 476120 155496
rect 311158 155428 311164 155440
rect 310348 155400 311164 155428
rect 311158 155388 311164 155400
rect 311216 155388 311222 155440
rect 311342 155388 311348 155440
rect 311400 155428 311406 155440
rect 326706 155428 326712 155440
rect 311400 155400 326712 155428
rect 311400 155388 311406 155400
rect 326706 155388 326712 155400
rect 326764 155388 326770 155440
rect 327902 155388 327908 155440
rect 327960 155428 327966 155440
rect 338482 155428 338488 155440
rect 327960 155400 338488 155428
rect 327960 155388 327966 155400
rect 338482 155388 338488 155400
rect 338540 155388 338546 155440
rect 398558 155388 398564 155440
rect 398616 155428 398622 155440
rect 398616 155400 407436 155428
rect 398616 155388 398622 155400
rect 318978 155360 318984 155372
rect 302206 155332 318984 155360
rect 301317 155323 301375 155329
rect 318978 155320 318984 155332
rect 319036 155320 319042 155372
rect 321094 155320 321100 155372
rect 321152 155360 321158 155372
rect 334158 155360 334164 155372
rect 321152 155332 334164 155360
rect 321152 155320 321158 155332
rect 334158 155320 334164 155332
rect 334216 155320 334222 155372
rect 382274 155320 382280 155372
rect 382332 155360 382338 155372
rect 386414 155360 386420 155372
rect 382332 155332 386420 155360
rect 382332 155320 382338 155332
rect 386414 155320 386420 155332
rect 386472 155320 386478 155372
rect 401594 155320 401600 155372
rect 401652 155360 401658 155372
rect 404906 155360 404912 155372
rect 401652 155332 404912 155360
rect 401652 155320 401658 155332
rect 404906 155320 404912 155332
rect 404964 155320 404970 155372
rect 407408 155360 407436 155400
rect 411162 155388 411168 155440
rect 411220 155428 411226 155440
rect 436094 155428 436100 155440
rect 411220 155400 436100 155428
rect 411220 155388 411226 155400
rect 436094 155388 436100 155400
rect 436152 155388 436158 155440
rect 438026 155388 438032 155440
rect 438084 155428 438090 155440
rect 438228 155428 438256 155468
rect 476114 155456 476120 155468
rect 476172 155456 476178 155508
rect 484762 155456 484768 155508
rect 484820 155496 484826 155508
rect 546310 155496 546316 155508
rect 484820 155468 546316 155496
rect 484820 155456 484826 155468
rect 546310 155456 546316 155468
rect 546368 155456 546374 155508
rect 438084 155400 438256 155428
rect 438084 155388 438090 155400
rect 441246 155388 441252 155440
rect 441304 155428 441310 155440
rect 480990 155428 480996 155440
rect 441304 155400 480996 155428
rect 441304 155388 441310 155400
rect 480990 155388 480996 155400
rect 481048 155388 481054 155440
rect 483566 155388 483572 155440
rect 483624 155428 483630 155440
rect 544286 155428 544292 155440
rect 483624 155400 544292 155428
rect 483624 155388 483630 155400
rect 544286 155388 544292 155400
rect 544344 155388 544350 155440
rect 417602 155360 417608 155372
rect 407408 155332 417608 155360
rect 417602 155320 417608 155332
rect 417660 155320 417666 155372
rect 417970 155320 417976 155372
rect 418028 155360 418034 155372
rect 444926 155360 444932 155372
rect 418028 155332 444932 155360
rect 418028 155320 418034 155332
rect 444926 155320 444932 155332
rect 444984 155320 444990 155372
rect 445662 155320 445668 155372
rect 445720 155360 445726 155372
rect 484854 155360 484860 155372
rect 445720 155332 484860 155360
rect 445720 155320 445726 155332
rect 484854 155320 484860 155332
rect 484912 155320 484918 155372
rect 488350 155320 488356 155372
rect 488408 155360 488414 155372
rect 552106 155360 552112 155372
rect 488408 155332 552112 155360
rect 488408 155320 488414 155332
rect 552106 155320 552112 155332
rect 552164 155320 552170 155372
rect 137373 155295 137431 155301
rect 137373 155261 137385 155295
rect 137419 155261 137431 155295
rect 137373 155255 137431 155261
rect 138017 155295 138075 155301
rect 138017 155261 138029 155295
rect 138063 155292 138075 155295
rect 203061 155295 203119 155301
rect 203061 155292 203073 155295
rect 138063 155264 203073 155292
rect 138063 155261 138075 155264
rect 138017 155255 138075 155261
rect 203061 155261 203073 155264
rect 203107 155261 203119 155295
rect 203061 155255 203119 155261
rect 137388 155224 137416 155255
rect 203150 155252 203156 155304
rect 203208 155292 203214 155304
rect 213181 155295 213239 155301
rect 213181 155292 213193 155295
rect 203208 155264 213193 155292
rect 203208 155252 203214 155264
rect 213181 155261 213193 155264
rect 213227 155261 213239 155295
rect 213181 155255 213239 155261
rect 214469 155295 214527 155301
rect 214469 155261 214481 155295
rect 214515 155292 214527 155295
rect 219345 155295 219403 155301
rect 219345 155292 219357 155295
rect 214515 155264 219357 155292
rect 214515 155261 214527 155264
rect 214469 155255 214527 155261
rect 219345 155261 219357 155264
rect 219391 155261 219403 155295
rect 219345 155255 219403 155261
rect 219437 155295 219495 155301
rect 219437 155261 219449 155295
rect 219483 155292 219495 155295
rect 220630 155292 220636 155304
rect 219483 155264 220636 155292
rect 219483 155261 219495 155264
rect 219437 155255 219495 155261
rect 220630 155252 220636 155264
rect 220688 155252 220694 155304
rect 221553 155295 221611 155301
rect 221553 155261 221565 155295
rect 221599 155292 221611 155295
rect 223577 155295 223635 155301
rect 223577 155292 223589 155295
rect 221599 155264 223589 155292
rect 221599 155261 221611 155264
rect 221553 155255 221611 155261
rect 223577 155261 223589 155264
rect 223623 155261 223635 155295
rect 223577 155255 223635 155261
rect 223666 155252 223672 155304
rect 223724 155292 223730 155304
rect 269022 155292 269028 155304
rect 223724 155264 269028 155292
rect 223724 155252 223730 155264
rect 269022 155252 269028 155264
rect 269080 155252 269086 155304
rect 270402 155252 270408 155304
rect 270460 155292 270466 155304
rect 270460 155264 273944 155292
rect 270460 155252 270466 155264
rect 202141 155227 202199 155233
rect 202141 155224 202153 155227
rect 137388 155196 202153 155224
rect 202141 155193 202153 155196
rect 202187 155193 202199 155227
rect 202141 155187 202199 155193
rect 202230 155184 202236 155236
rect 202288 155224 202294 155236
rect 206005 155227 206063 155233
rect 206005 155224 206017 155227
rect 202288 155196 206017 155224
rect 202288 155184 202294 155196
rect 206005 155193 206017 155196
rect 206051 155193 206063 155227
rect 206005 155187 206063 155193
rect 206097 155227 206155 155233
rect 206097 155193 206109 155227
rect 206143 155224 206155 155227
rect 209038 155224 209044 155236
rect 206143 155196 209044 155224
rect 206143 155193 206155 155196
rect 206097 155187 206155 155193
rect 209038 155184 209044 155196
rect 209096 155184 209102 155236
rect 210970 155184 210976 155236
rect 211028 155224 211034 155236
rect 249245 155227 249303 155233
rect 211028 155196 249196 155224
rect 211028 155184 211034 155196
rect 52144 155128 137324 155156
rect 137373 155159 137431 155165
rect 52144 155116 52150 155128
rect 137373 155125 137385 155159
rect 137419 155156 137431 155159
rect 143629 155159 143687 155165
rect 143629 155156 143641 155159
rect 137419 155128 143641 155156
rect 137419 155125 137431 155128
rect 137373 155119 137431 155125
rect 143629 155125 143641 155128
rect 143675 155125 143687 155159
rect 143629 155119 143687 155125
rect 143721 155159 143779 155165
rect 143721 155125 143733 155159
rect 143767 155156 143779 155159
rect 146849 155159 146907 155165
rect 146849 155156 146861 155159
rect 143767 155128 146861 155156
rect 143767 155125 143779 155128
rect 143721 155119 143779 155125
rect 146849 155125 146861 155128
rect 146895 155125 146907 155159
rect 146849 155119 146907 155125
rect 146941 155159 146999 155165
rect 146941 155125 146953 155159
rect 146987 155156 146999 155159
rect 185578 155156 185584 155168
rect 146987 155128 185584 155156
rect 146987 155125 146999 155128
rect 146941 155119 146999 155125
rect 185578 155116 185584 155128
rect 185636 155116 185642 155168
rect 185673 155159 185731 155165
rect 185673 155125 185685 155159
rect 185719 155156 185731 155159
rect 240226 155156 240232 155168
rect 185719 155128 240232 155156
rect 185719 155125 185731 155128
rect 185673 155119 185731 155125
rect 240226 155116 240232 155128
rect 240284 155116 240290 155168
rect 241977 155159 242035 155165
rect 241977 155125 241989 155159
rect 242023 155156 242035 155159
rect 242023 155128 243584 155156
rect 242023 155125 242035 155128
rect 241977 155119 242035 155125
rect 39390 155048 39396 155100
rect 39448 155088 39454 155100
rect 124122 155088 124128 155100
rect 39448 155060 124128 155088
rect 39448 155048 39454 155060
rect 124122 155048 124128 155060
rect 124180 155048 124186 155100
rect 124769 155091 124827 155097
rect 124769 155057 124781 155091
rect 124815 155088 124827 155091
rect 127437 155091 127495 155097
rect 127437 155088 127449 155091
rect 124815 155060 127449 155088
rect 124815 155057 124827 155060
rect 124769 155051 124827 155057
rect 127437 155057 127449 155060
rect 127483 155057 127495 155091
rect 127437 155051 127495 155057
rect 127529 155091 127587 155097
rect 127529 155057 127541 155091
rect 127575 155088 127587 155091
rect 127713 155091 127771 155097
rect 127713 155088 127725 155091
rect 127575 155060 127725 155088
rect 127575 155057 127587 155060
rect 127529 155051 127587 155057
rect 127713 155057 127725 155060
rect 127759 155057 127771 155091
rect 127713 155051 127771 155057
rect 128817 155091 128875 155097
rect 128817 155057 128829 155091
rect 128863 155088 128875 155091
rect 202874 155088 202880 155100
rect 128863 155060 202880 155088
rect 128863 155057 128875 155060
rect 128817 155051 128875 155057
rect 202874 155048 202880 155060
rect 202932 155048 202938 155100
rect 202969 155091 203027 155097
rect 202969 155057 202981 155091
rect 203015 155088 203027 155091
rect 209869 155091 209927 155097
rect 209869 155088 209881 155091
rect 203015 155060 209881 155088
rect 203015 155057 203027 155060
rect 202969 155051 203027 155057
rect 209869 155057 209881 155060
rect 209915 155057 209927 155091
rect 209869 155051 209927 155057
rect 209958 155048 209964 155100
rect 210016 155088 210022 155100
rect 214469 155091 214527 155097
rect 214469 155088 214481 155091
rect 210016 155060 214481 155088
rect 210016 155048 210022 155060
rect 214469 155057 214481 155060
rect 214515 155057 214527 155091
rect 214469 155051 214527 155057
rect 214561 155091 214619 155097
rect 214561 155057 214573 155091
rect 214607 155088 214619 155091
rect 243446 155088 243452 155100
rect 214607 155060 243452 155088
rect 214607 155057 214619 155060
rect 214561 155051 214619 155057
rect 243446 155048 243452 155060
rect 243504 155048 243510 155100
rect 243556 155088 243584 155128
rect 244826 155088 244832 155100
rect 243556 155060 244832 155088
rect 244826 155048 244832 155060
rect 244884 155048 244890 155100
rect 244921 155091 244979 155097
rect 244921 155057 244933 155091
rect 244967 155088 244979 155091
rect 249061 155091 249119 155097
rect 249061 155088 249073 155091
rect 244967 155060 249073 155088
rect 244967 155057 244979 155060
rect 244921 155051 244979 155057
rect 249061 155057 249073 155060
rect 249107 155057 249119 155091
rect 249168 155088 249196 155196
rect 249245 155193 249257 155227
rect 249291 155224 249303 155227
rect 252646 155224 252652 155236
rect 249291 155196 252652 155224
rect 249291 155193 249303 155196
rect 249245 155187 249303 155193
rect 252646 155184 252652 155196
rect 252704 155184 252710 155236
rect 253842 155184 253848 155236
rect 253900 155224 253906 155236
rect 262953 155227 263011 155233
rect 262953 155224 262965 155227
rect 253900 155196 262965 155224
rect 253900 155184 253906 155196
rect 262953 155193 262965 155196
rect 262999 155193 263011 155227
rect 262953 155187 263011 155193
rect 264149 155227 264207 155233
rect 264149 155193 264161 155227
rect 264195 155224 264207 155227
rect 272613 155227 272671 155233
rect 272613 155224 272625 155227
rect 264195 155196 272625 155224
rect 264195 155193 264207 155196
rect 264149 155187 264207 155193
rect 272613 155193 272625 155196
rect 272659 155193 272671 155227
rect 273916 155224 273944 155264
rect 275278 155252 275284 155304
rect 275336 155292 275342 155304
rect 296717 155295 296775 155301
rect 296717 155292 296729 155295
rect 275336 155264 296729 155292
rect 275336 155252 275342 155264
rect 296717 155261 296729 155264
rect 296763 155261 296775 155295
rect 300118 155292 300124 155304
rect 296717 155255 296775 155261
rect 296824 155264 300124 155292
rect 296824 155224 296852 155264
rect 300118 155252 300124 155264
rect 300176 155252 300182 155304
rect 301590 155252 301596 155304
rect 301648 155292 301654 155304
rect 307113 155295 307171 155301
rect 307113 155292 307125 155295
rect 301648 155264 307125 155292
rect 301648 155252 301654 155264
rect 307113 155261 307125 155264
rect 307159 155261 307171 155295
rect 307113 155255 307171 155261
rect 308490 155252 308496 155304
rect 308548 155292 308554 155304
rect 324406 155292 324412 155304
rect 308548 155264 324412 155292
rect 308548 155252 308554 155264
rect 324406 155252 324412 155264
rect 324464 155252 324470 155304
rect 331858 155252 331864 155304
rect 331916 155292 331922 155304
rect 337930 155292 337936 155304
rect 331916 155264 337936 155292
rect 331916 155252 331922 155264
rect 337930 155252 337936 155264
rect 337988 155252 337994 155304
rect 402238 155252 402244 155304
rect 402296 155292 402302 155304
rect 422478 155292 422484 155304
rect 402296 155264 422484 155292
rect 402296 155252 402302 155264
rect 422478 155252 422484 155264
rect 422536 155252 422542 155304
rect 424962 155252 424968 155304
rect 425020 155292 425026 155304
rect 456610 155292 456616 155304
rect 425020 155264 456616 155292
rect 425020 155252 425026 155264
rect 456610 155252 456616 155264
rect 456668 155252 456674 155304
rect 456702 155252 456708 155304
rect 456760 155292 456766 155304
rect 502426 155292 502432 155304
rect 456760 155264 502432 155292
rect 456760 155252 456766 155264
rect 502426 155252 502432 155264
rect 502484 155252 502490 155304
rect 502978 155252 502984 155304
rect 503036 155292 503042 155304
rect 569678 155292 569684 155304
rect 503036 155264 569684 155292
rect 503036 155252 503042 155264
rect 569678 155252 569684 155264
rect 569736 155252 569742 155304
rect 273916 155196 296852 155224
rect 272613 155187 272671 155193
rect 296898 155184 296904 155236
rect 296956 155224 296962 155236
rect 304902 155224 304908 155236
rect 296956 155196 304908 155224
rect 296956 155184 296962 155196
rect 304902 155184 304908 155196
rect 304960 155184 304966 155236
rect 305546 155184 305552 155236
rect 305604 155224 305610 155236
rect 322842 155224 322848 155236
rect 305604 155196 322848 155224
rect 305604 155184 305610 155196
rect 322842 155184 322848 155196
rect 322900 155184 322906 155236
rect 323026 155184 323032 155236
rect 323084 155224 323090 155236
rect 334066 155224 334072 155236
rect 323084 155196 334072 155224
rect 323084 155184 323090 155196
rect 334066 155184 334072 155196
rect 334124 155184 334130 155236
rect 343542 155184 343548 155236
rect 343600 155224 343606 155236
rect 349062 155224 349068 155236
rect 343600 155196 349068 155224
rect 343600 155184 343606 155196
rect 349062 155184 349068 155196
rect 349120 155184 349126 155236
rect 384850 155184 384856 155236
rect 384908 155224 384914 155236
rect 388346 155224 388352 155236
rect 384908 155196 388352 155224
rect 384908 155184 384914 155196
rect 388346 155184 388352 155196
rect 388404 155184 388410 155236
rect 401502 155184 401508 155236
rect 401560 155224 401566 155236
rect 421558 155224 421564 155236
rect 401560 155196 421564 155224
rect 401560 155184 401566 155196
rect 421558 155184 421564 155196
rect 421616 155184 421622 155236
rect 422018 155184 422024 155236
rect 422076 155224 422082 155236
rect 452746 155224 452752 155236
rect 422076 155196 452752 155224
rect 422076 155184 422082 155196
rect 452746 155184 452752 155196
rect 452804 155184 452810 155236
rect 454862 155184 454868 155236
rect 454920 155224 454926 155236
rect 501414 155224 501420 155236
rect 454920 155196 501420 155224
rect 454920 155184 454926 155196
rect 501414 155184 501420 155196
rect 501472 155184 501478 155236
rect 502242 155184 502248 155236
rect 502300 155224 502306 155236
rect 572622 155224 572628 155236
rect 502300 155196 572628 155224
rect 502300 155184 502306 155196
rect 572622 155184 572628 155196
rect 572680 155184 572686 155236
rect 249978 155116 249984 155168
rect 250036 155156 250042 155168
rect 277397 155159 277455 155165
rect 277397 155156 277409 155159
rect 250036 155128 277409 155156
rect 250036 155116 250042 155128
rect 277397 155125 277409 155128
rect 277443 155125 277455 155159
rect 277397 155119 277455 155125
rect 277489 155159 277547 155165
rect 277489 155125 277501 155159
rect 277535 155156 277547 155159
rect 281442 155156 281448 155168
rect 277535 155128 281448 155156
rect 277535 155125 277547 155128
rect 277489 155119 277547 155125
rect 281442 155116 281448 155128
rect 281500 155116 281506 155168
rect 282181 155159 282239 155165
rect 282181 155125 282193 155159
rect 282227 155156 282239 155159
rect 288621 155159 288679 155165
rect 288621 155156 288633 155159
rect 282227 155128 288633 155156
rect 282227 155125 282239 155128
rect 282181 155119 282239 155125
rect 288621 155125 288633 155128
rect 288667 155125 288679 155159
rect 288621 155119 288679 155125
rect 288713 155159 288771 155165
rect 288713 155125 288725 155159
rect 288759 155156 288771 155159
rect 297910 155156 297916 155168
rect 288759 155128 297916 155156
rect 288759 155125 288771 155128
rect 288713 155119 288771 155125
rect 297910 155116 297916 155128
rect 297968 155116 297974 155168
rect 298649 155159 298707 155165
rect 298649 155125 298661 155159
rect 298695 155156 298707 155159
rect 301409 155159 301467 155165
rect 301409 155156 301421 155159
rect 298695 155128 301421 155156
rect 298695 155125 298707 155128
rect 298649 155119 298707 155125
rect 301409 155125 301421 155128
rect 301455 155125 301467 155159
rect 301409 155119 301467 155125
rect 301501 155159 301559 155165
rect 301501 155125 301513 155159
rect 301547 155156 301559 155159
rect 306929 155159 306987 155165
rect 306929 155156 306941 155159
rect 301547 155128 306941 155156
rect 301547 155125 301559 155128
rect 301501 155119 301559 155125
rect 306929 155125 306941 155128
rect 306975 155125 306987 155159
rect 306929 155119 306987 155125
rect 307205 155159 307263 155165
rect 307205 155125 307217 155159
rect 307251 155156 307263 155159
rect 316402 155156 316408 155168
rect 307251 155128 316408 155156
rect 307251 155125 307263 155128
rect 307205 155119 307263 155125
rect 316402 155116 316408 155128
rect 316460 155116 316466 155168
rect 320082 155156 320088 155168
rect 317156 155128 320088 155156
rect 259362 155088 259368 155100
rect 249168 155060 259368 155088
rect 249061 155051 249119 155057
rect 259362 155048 259368 155060
rect 259420 155048 259426 155100
rect 259457 155091 259515 155097
rect 259457 155057 259469 155091
rect 259503 155088 259515 155091
rect 262677 155091 262735 155097
rect 262677 155088 262689 155091
rect 259503 155060 262689 155088
rect 259503 155057 259515 155060
rect 259457 155051 259515 155057
rect 262677 155057 262689 155060
rect 262723 155057 262735 155091
rect 262677 155051 262735 155057
rect 262769 155091 262827 155097
rect 262769 155057 262781 155091
rect 262815 155088 262827 155091
rect 282089 155091 282147 155097
rect 282089 155088 282101 155091
rect 262815 155060 282101 155088
rect 262815 155057 262827 155060
rect 262769 155051 262827 155057
rect 282089 155057 282101 155060
rect 282135 155057 282147 155091
rect 282089 155051 282147 155057
rect 285030 155048 285036 155100
rect 285088 155088 285094 155100
rect 291841 155091 291899 155097
rect 291841 155088 291853 155091
rect 285088 155060 291853 155088
rect 285088 155048 285094 155060
rect 291841 155057 291853 155060
rect 291887 155057 291899 155091
rect 291841 155051 291899 155057
rect 292853 155091 292911 155097
rect 292853 155057 292865 155091
rect 292899 155088 292911 155091
rect 302234 155088 302240 155100
rect 292899 155060 302240 155088
rect 292899 155057 292911 155060
rect 292853 155051 292911 155057
rect 302234 155048 302240 155060
rect 302292 155048 302298 155100
rect 302329 155091 302387 155097
rect 302329 155057 302341 155091
rect 302375 155088 302387 155091
rect 314654 155088 314660 155100
rect 302375 155060 314660 155088
rect 302375 155057 302387 155060
rect 302329 155051 302387 155057
rect 314654 155048 314660 155060
rect 314712 155048 314718 155100
rect 317156 155088 317184 155128
rect 320082 155116 320088 155128
rect 320140 155116 320146 155168
rect 324038 155116 324044 155168
rect 324096 155156 324102 155168
rect 333974 155156 333980 155168
rect 324096 155128 333980 155156
rect 324096 155116 324102 155128
rect 333974 155116 333980 155128
rect 334032 155116 334038 155168
rect 355226 155116 355232 155168
rect 355284 155156 355290 155168
rect 356698 155156 356704 155168
rect 355284 155128 356704 155156
rect 355284 155116 355290 155128
rect 356698 155116 356704 155128
rect 356756 155116 356762 155168
rect 405918 155116 405924 155168
rect 405976 155156 405982 155168
rect 409782 155156 409788 155168
rect 405976 155128 409788 155156
rect 405976 155116 405982 155128
rect 409782 155116 409788 155128
rect 409840 155116 409846 155168
rect 409877 155159 409935 155165
rect 409877 155125 409889 155159
rect 409923 155156 409935 155159
rect 426342 155156 426348 155168
rect 409923 155128 426348 155156
rect 409923 155125 409935 155128
rect 409877 155119 409935 155125
rect 426342 155116 426348 155128
rect 426400 155116 426406 155168
rect 428274 155116 428280 155168
rect 428332 155156 428338 155168
rect 428332 155128 460934 155156
rect 428332 155116 428338 155128
rect 316006 155060 317184 155088
rect 86218 154980 86224 155032
rect 86276 155020 86282 155032
rect 156141 155023 156199 155029
rect 156141 155020 156153 155023
rect 86276 154992 156153 155020
rect 86276 154980 86282 154992
rect 156141 154989 156153 154992
rect 156187 154989 156199 155023
rect 166994 155020 167000 155032
rect 156141 154983 156199 154989
rect 156248 154992 167000 155020
rect 74534 154912 74540 154964
rect 74592 154952 74598 154964
rect 143537 154955 143595 154961
rect 143537 154952 143549 154955
rect 74592 154924 143549 154952
rect 74592 154912 74598 154924
rect 143537 154921 143549 154924
rect 143583 154921 143595 154955
rect 143537 154915 143595 154921
rect 143629 154955 143687 154961
rect 143629 154921 143641 154955
rect 143675 154952 143687 154955
rect 156248 154952 156276 154992
rect 166994 154980 167000 154992
rect 167052 154980 167058 155032
rect 167086 154980 167092 155032
rect 167144 155020 167150 155032
rect 171137 155023 171195 155029
rect 171137 155020 171149 155023
rect 167144 154992 171149 155020
rect 167144 154980 167150 154992
rect 171137 154989 171149 154992
rect 171183 154989 171195 155023
rect 171137 154983 171195 154989
rect 171226 154980 171232 155032
rect 171284 155020 171290 155032
rect 182082 155020 182088 155032
rect 171284 154992 182088 155020
rect 171284 154980 171290 154992
rect 182082 154980 182088 154992
rect 182140 154980 182146 155032
rect 187602 154980 187608 155032
rect 187660 155020 187666 155032
rect 195241 155023 195299 155029
rect 187660 154992 194916 155020
rect 187660 154980 187666 154992
rect 143675 154924 156276 154952
rect 156417 154955 156475 154961
rect 143675 154921 143687 154924
rect 143629 154915 143687 154921
rect 156417 154921 156429 154955
rect 156463 154952 156475 154955
rect 194888 154952 194916 154992
rect 195241 154989 195253 155023
rect 195287 155020 195299 155023
rect 242250 155020 242256 155032
rect 195287 154992 242256 155020
rect 195287 154989 195299 154992
rect 195241 154983 195299 154989
rect 242250 154980 242256 154992
rect 242308 154980 242314 155032
rect 243541 155023 243599 155029
rect 243541 154989 243553 155023
rect 243587 155020 243599 155023
rect 268289 155023 268347 155029
rect 268289 155020 268301 155023
rect 243587 154992 268301 155020
rect 243587 154989 243599 154992
rect 243541 154983 243599 154989
rect 268289 154989 268301 154992
rect 268335 154989 268347 155023
rect 272429 155023 272487 155029
rect 272429 155020 272441 155023
rect 268289 154983 268347 154989
rect 268396 154992 272441 155020
rect 241977 154955 242035 154961
rect 241977 154952 241989 154955
rect 156463 154924 194364 154952
rect 194888 154924 241989 154952
rect 156463 154921 156475 154924
rect 156417 154915 156475 154921
rect 474 154844 480 154896
rect 532 154884 538 154896
rect 1302 154884 1308 154896
rect 532 154856 1308 154884
rect 532 154844 538 154856
rect 1302 154844 1308 154856
rect 1360 154844 1366 154896
rect 97902 154844 97908 154896
rect 97960 154884 97966 154896
rect 169754 154884 169760 154896
rect 97960 154856 169760 154884
rect 97960 154844 97966 154856
rect 169754 154844 169760 154856
rect 169812 154844 169818 154896
rect 171137 154887 171195 154893
rect 171137 154853 171149 154887
rect 171183 154884 171195 154887
rect 175826 154884 175832 154896
rect 171183 154856 175832 154884
rect 171183 154853 171195 154856
rect 171137 154847 171195 154853
rect 175826 154844 175832 154856
rect 175884 154844 175890 154896
rect 176838 154844 176844 154896
rect 176896 154884 176902 154896
rect 177942 154884 177948 154896
rect 176896 154856 177948 154884
rect 176896 154844 176902 154856
rect 177942 154844 177948 154856
rect 178000 154844 178006 154896
rect 190457 154887 190515 154893
rect 190457 154853 190469 154887
rect 190503 154884 190515 154887
rect 194226 154884 194232 154896
rect 190503 154856 194232 154884
rect 190503 154853 190515 154856
rect 190457 154847 190515 154853
rect 194226 154844 194232 154856
rect 194284 154844 194290 154896
rect 94958 154776 94964 154828
rect 95016 154816 95022 154828
rect 137373 154819 137431 154825
rect 137373 154816 137385 154819
rect 95016 154788 137385 154816
rect 95016 154776 95022 154788
rect 137373 154785 137385 154788
rect 137419 154785 137431 154819
rect 137373 154779 137431 154785
rect 137465 154819 137523 154825
rect 137465 154785 137477 154819
rect 137511 154816 137523 154819
rect 193122 154816 193128 154828
rect 137511 154788 193128 154816
rect 137511 154785 137523 154788
rect 137465 154779 137523 154785
rect 193122 154776 193128 154788
rect 193180 154776 193186 154828
rect 194336 154816 194364 154924
rect 241977 154921 241989 154924
rect 242023 154921 242035 154955
rect 241977 154915 242035 154921
rect 242069 154955 242127 154961
rect 242069 154921 242081 154955
rect 242115 154952 242127 154955
rect 242115 154924 245056 154952
rect 242115 154921 242127 154924
rect 242069 154915 242127 154921
rect 194410 154844 194416 154896
rect 194468 154884 194474 154896
rect 197449 154887 197507 154893
rect 197449 154884 197461 154887
rect 194468 154856 197461 154884
rect 194468 154844 194474 154856
rect 197449 154853 197461 154856
rect 197495 154853 197507 154887
rect 197449 154847 197507 154853
rect 197541 154887 197599 154893
rect 197541 154853 197553 154887
rect 197587 154884 197599 154887
rect 241057 154887 241115 154893
rect 241057 154884 241069 154887
rect 197587 154856 241069 154884
rect 197587 154853 197599 154856
rect 197541 154847 197599 154853
rect 241057 154853 241069 154856
rect 241103 154853 241115 154887
rect 241057 154847 241115 154853
rect 241146 154844 241152 154896
rect 241204 154884 241210 154896
rect 244277 154887 244335 154893
rect 244277 154884 244289 154887
rect 241204 154856 244289 154884
rect 241204 154844 241210 154856
rect 244277 154853 244289 154856
rect 244323 154853 244335 154887
rect 244921 154887 244979 154893
rect 244921 154884 244933 154887
rect 244277 154847 244335 154853
rect 244384 154856 244933 154884
rect 195514 154816 195520 154828
rect 194336 154788 195520 154816
rect 195514 154776 195520 154788
rect 195572 154776 195578 154828
rect 204809 154819 204867 154825
rect 204809 154816 204821 154819
rect 197740 154788 204821 154816
rect 78398 154708 78404 154760
rect 78456 154748 78462 154760
rect 110414 154748 110420 154760
rect 78456 154720 110420 154748
rect 78456 154708 78462 154720
rect 110414 154708 110420 154720
rect 110472 154708 110478 154760
rect 113542 154708 113548 154760
rect 113600 154748 113606 154760
rect 117869 154751 117927 154757
rect 113600 154720 117820 154748
rect 113600 154708 113606 154720
rect 56962 154640 56968 154692
rect 57020 154680 57026 154692
rect 116762 154680 116768 154692
rect 57020 154652 116768 154680
rect 57020 154640 57026 154652
rect 116762 154640 116768 154652
rect 116820 154640 116826 154692
rect 117792 154680 117820 154720
rect 117869 154717 117881 154751
rect 117915 154748 117927 154751
rect 120718 154748 120724 154760
rect 117915 154720 120724 154748
rect 117915 154717 117927 154720
rect 117869 154711 117927 154717
rect 120718 154708 120724 154720
rect 120776 154708 120782 154760
rect 178034 154748 178040 154760
rect 120828 154720 178040 154748
rect 120828 154680 120856 154720
rect 178034 154708 178040 154720
rect 178092 154708 178098 154760
rect 178770 154708 178776 154760
rect 178828 154748 178834 154760
rect 186314 154748 186320 154760
rect 178828 154720 186320 154748
rect 178828 154708 178834 154720
rect 186314 154708 186320 154720
rect 186372 154708 186378 154760
rect 194962 154748 194968 154760
rect 190426 154720 194968 154748
rect 117792 154652 120856 154680
rect 121270 154640 121276 154692
rect 121328 154680 121334 154692
rect 127621 154683 127679 154689
rect 127621 154680 127633 154683
rect 121328 154652 127633 154680
rect 121328 154640 121334 154652
rect 127621 154649 127633 154652
rect 127667 154649 127679 154683
rect 127621 154643 127679 154649
rect 127713 154683 127771 154689
rect 127713 154649 127725 154683
rect 127759 154680 127771 154683
rect 182082 154680 182088 154692
rect 127759 154652 182088 154680
rect 127759 154649 127771 154652
rect 127713 154643 127771 154649
rect 182082 154640 182088 154652
rect 182140 154640 182146 154692
rect 182726 154640 182732 154692
rect 182784 154680 182790 154692
rect 190426 154680 190454 154720
rect 194962 154708 194968 154720
rect 195020 154708 195026 154760
rect 195330 154708 195336 154760
rect 195388 154748 195394 154760
rect 197740 154748 197768 154788
rect 204809 154785 204821 154788
rect 204855 154785 204867 154819
rect 244384 154816 244412 154856
rect 244921 154853 244933 154856
rect 244967 154853 244979 154887
rect 245028 154884 245056 154924
rect 245102 154912 245108 154964
rect 245160 154952 245166 154964
rect 268396 154952 268424 154992
rect 272429 154989 272441 154992
rect 272475 154989 272487 155023
rect 272429 154983 272487 154989
rect 272521 155023 272579 155029
rect 272521 154989 272533 155023
rect 272567 155020 272579 155023
rect 277397 155023 277455 155029
rect 277397 155020 277409 155023
rect 272567 154992 277409 155020
rect 272567 154989 272579 154992
rect 272521 154983 272579 154989
rect 277397 154989 277409 154992
rect 277443 154989 277455 155023
rect 277397 154983 277455 154989
rect 277486 154980 277492 155032
rect 277544 155020 277550 155032
rect 285674 155020 285680 155032
rect 277544 154992 285680 155020
rect 277544 154980 277550 154992
rect 285674 154980 285680 154992
rect 285732 154980 285738 155032
rect 285769 155023 285827 155029
rect 285769 154989 285781 155023
rect 285815 155020 285827 155023
rect 285815 154992 297680 155020
rect 285815 154989 285827 154992
rect 285769 154983 285827 154989
rect 245160 154924 268424 154952
rect 245160 154912 245166 154924
rect 268470 154912 268476 154964
rect 268528 154952 268534 154964
rect 276201 154955 276259 154961
rect 276201 154952 276213 154955
rect 268528 154924 276213 154952
rect 268528 154912 268534 154924
rect 276201 154921 276213 154924
rect 276247 154921 276259 154955
rect 276201 154915 276259 154921
rect 276290 154912 276296 154964
rect 276348 154952 276354 154964
rect 282181 154955 282239 154961
rect 282181 154952 282193 154955
rect 276348 154924 282193 154952
rect 276348 154912 276354 154924
rect 282181 154921 282193 154924
rect 282227 154921 282239 154955
rect 282181 154915 282239 154921
rect 282273 154955 282331 154961
rect 282273 154921 282285 154955
rect 282319 154952 282331 154955
rect 296901 154955 296959 154961
rect 296901 154952 296913 154955
rect 282319 154924 296913 154952
rect 282319 154921 282331 154924
rect 282273 154915 282331 154921
rect 296901 154921 296913 154924
rect 296947 154921 296959 154955
rect 297652 154952 297680 154992
rect 297726 154980 297732 155032
rect 297784 155020 297790 155032
rect 306929 155023 306987 155029
rect 306929 155020 306941 155023
rect 297784 154992 306941 155020
rect 297784 154980 297790 154992
rect 306929 154989 306941 154992
rect 306975 154989 306987 155023
rect 306929 154983 306987 154989
rect 307036 154992 307248 155020
rect 302513 154955 302571 154961
rect 302513 154952 302525 154955
rect 297652 154924 302525 154952
rect 296901 154915 296959 154921
rect 302513 154921 302525 154924
rect 302559 154921 302571 154955
rect 302513 154915 302571 154921
rect 302602 154912 302608 154964
rect 302660 154952 302666 154964
rect 307036 154952 307064 154992
rect 302660 154924 307064 154952
rect 307220 154952 307248 154992
rect 307478 154980 307484 155032
rect 307536 155020 307542 155032
rect 316006 155020 316034 155060
rect 317230 155048 317236 155100
rect 317288 155088 317294 155100
rect 326890 155088 326896 155100
rect 317288 155060 326896 155088
rect 317288 155048 317294 155060
rect 326890 155048 326896 155060
rect 326948 155048 326954 155100
rect 326982 155048 326988 155100
rect 327040 155088 327046 155100
rect 338022 155088 338028 155100
rect 327040 155060 338028 155088
rect 327040 155048 327046 155060
rect 338022 155048 338028 155060
rect 338080 155048 338086 155100
rect 356238 155048 356244 155100
rect 356296 155088 356302 155100
rect 357434 155088 357440 155100
rect 356296 155060 357440 155088
rect 356296 155048 356302 155060
rect 357434 155048 357440 155060
rect 357492 155048 357498 155100
rect 400306 155048 400312 155100
rect 400364 155088 400370 155100
rect 402054 155088 402060 155100
rect 400364 155060 402060 155088
rect 400364 155048 400370 155060
rect 402054 155048 402060 155060
rect 402112 155048 402118 155100
rect 418614 155088 418620 155100
rect 402164 155060 418620 155088
rect 321554 155020 321560 155032
rect 307536 154992 316034 155020
rect 316098 154992 321560 155020
rect 307536 154980 307542 154992
rect 316098 154952 316126 154992
rect 321554 154980 321560 154992
rect 321612 154980 321618 155032
rect 325050 154980 325056 155032
rect 325108 155020 325114 155032
rect 336642 155020 336648 155032
rect 325108 154992 336648 155020
rect 325108 154980 325114 154992
rect 336642 154980 336648 154992
rect 336700 154980 336706 155032
rect 399570 154980 399576 155032
rect 399628 155020 399634 155032
rect 402164 155020 402192 155060
rect 418614 155048 418620 155060
rect 418672 155048 418678 155100
rect 424410 155088 424416 155100
rect 418724 155060 424416 155088
rect 399628 154992 402192 155020
rect 402241 155023 402299 155029
rect 399628 154980 399634 154992
rect 402241 154989 402253 155023
rect 402287 155020 402299 155023
rect 413738 155020 413744 155032
rect 402287 154992 413744 155020
rect 402287 154989 402299 154992
rect 402241 154983 402299 154989
rect 413738 154980 413744 154992
rect 413796 154980 413802 155032
rect 418724 155020 418752 155060
rect 424410 155048 424416 155060
rect 424468 155048 424474 155100
rect 425606 155048 425612 155100
rect 425664 155088 425670 155100
rect 457622 155088 457628 155100
rect 425664 155060 457628 155088
rect 425664 155048 425670 155060
rect 457622 155048 457628 155060
rect 457680 155048 457686 155100
rect 413848 154992 418752 155020
rect 319622 154952 319628 154964
rect 307220 154924 316126 154952
rect 316236 154924 319628 154952
rect 302660 154912 302666 154924
rect 248785 154887 248843 154893
rect 248785 154884 248797 154887
rect 245028 154856 248797 154884
rect 244921 154847 244979 154853
rect 248785 154853 248797 154856
rect 248831 154853 248843 154887
rect 248785 154847 248843 154853
rect 248877 154887 248935 154893
rect 248877 154853 248889 154887
rect 248923 154884 248935 154887
rect 255314 154884 255320 154896
rect 248923 154856 255320 154884
rect 248923 154853 248935 154856
rect 248877 154847 248935 154853
rect 255314 154844 255320 154856
rect 255372 154844 255378 154896
rect 262769 154887 262827 154893
rect 262769 154884 262781 154887
rect 256436 154856 262781 154884
rect 204809 154779 204867 154785
rect 204916 154788 244412 154816
rect 244461 154819 244519 154825
rect 195388 154720 197768 154748
rect 195388 154708 195394 154720
rect 199286 154708 199292 154760
rect 199344 154748 199350 154760
rect 204916 154748 204944 154788
rect 244461 154785 244473 154819
rect 244507 154816 244519 154819
rect 246942 154816 246948 154828
rect 244507 154788 246948 154816
rect 244507 154785 244519 154788
rect 244461 154779 244519 154785
rect 246942 154776 246948 154788
rect 247000 154776 247006 154828
rect 247034 154776 247040 154828
rect 247092 154816 247098 154828
rect 247402 154816 247408 154828
rect 247092 154788 247408 154816
rect 247092 154776 247098 154788
rect 247402 154776 247408 154788
rect 247460 154776 247466 154828
rect 248966 154776 248972 154828
rect 249024 154816 249030 154828
rect 254765 154819 254823 154825
rect 254765 154816 254777 154819
rect 249024 154788 254777 154816
rect 249024 154776 249030 154788
rect 254765 154785 254777 154788
rect 254811 154785 254823 154819
rect 254765 154779 254823 154785
rect 254854 154776 254860 154828
rect 254912 154816 254918 154828
rect 256436 154816 256464 154856
rect 262769 154853 262781 154856
rect 262815 154853 262827 154887
rect 262769 154847 262827 154853
rect 262858 154844 262864 154896
rect 262916 154884 262922 154896
rect 270402 154884 270408 154896
rect 262916 154856 270408 154884
rect 262916 154844 262922 154856
rect 270402 154844 270408 154856
rect 270460 154844 270466 154896
rect 272705 154887 272763 154893
rect 272705 154853 272717 154887
rect 272751 154884 272763 154887
rect 288529 154887 288587 154893
rect 288529 154884 288541 154887
rect 272751 154856 288541 154884
rect 272751 154853 272763 154856
rect 272705 154847 272763 154853
rect 288529 154853 288541 154856
rect 288575 154853 288587 154887
rect 288529 154847 288587 154853
rect 288621 154887 288679 154893
rect 288621 154853 288633 154887
rect 288667 154884 288679 154887
rect 291102 154884 291108 154896
rect 288667 154856 291108 154884
rect 288667 154853 288679 154856
rect 288621 154847 288679 154853
rect 291102 154844 291108 154856
rect 291160 154844 291166 154896
rect 292850 154844 292856 154896
rect 292908 154884 292914 154896
rect 296625 154887 296683 154893
rect 296625 154884 296637 154887
rect 292908 154856 296637 154884
rect 292908 154844 292914 154856
rect 296625 154853 296637 154856
rect 296671 154853 296683 154887
rect 296625 154847 296683 154853
rect 296717 154887 296775 154893
rect 296717 154853 296729 154887
rect 296763 154884 296775 154887
rect 306282 154884 306288 154896
rect 296763 154856 306288 154884
rect 296763 154853 296775 154856
rect 296717 154847 296775 154853
rect 306282 154844 306288 154856
rect 306340 154844 306346 154896
rect 307021 154887 307079 154893
rect 307021 154853 307033 154887
rect 307067 154884 307079 154887
rect 316236 154884 316264 154924
rect 319622 154912 319628 154924
rect 319680 154912 319686 154964
rect 325970 154912 325976 154964
rect 326028 154952 326034 154964
rect 337194 154952 337200 154964
rect 326028 154924 337200 154952
rect 326028 154912 326034 154924
rect 337194 154912 337200 154924
rect 337252 154912 337258 154964
rect 345474 154912 345480 154964
rect 345532 154952 345538 154964
rect 347590 154952 347596 154964
rect 345532 154924 347596 154952
rect 345532 154912 345538 154924
rect 347590 154912 347596 154924
rect 347648 154912 347654 154964
rect 357158 154912 357164 154964
rect 357216 154952 357222 154964
rect 357986 154952 357992 154964
rect 357216 154924 357992 154952
rect 357216 154912 357222 154924
rect 357986 154912 357992 154924
rect 358044 154912 358050 154964
rect 384206 154912 384212 154964
rect 384264 154952 384270 154964
rect 387426 154952 387432 154964
rect 384264 154924 387432 154952
rect 384264 154912 384270 154924
rect 387426 154912 387432 154924
rect 387484 154912 387490 154964
rect 400214 154912 400220 154964
rect 400272 154952 400278 154964
rect 402974 154952 402980 154964
rect 400272 154924 402980 154952
rect 400272 154912 400278 154924
rect 402974 154912 402980 154924
rect 403032 154912 403038 154964
rect 404722 154912 404728 154964
rect 404780 154952 404786 154964
rect 409877 154955 409935 154961
rect 409877 154952 409889 154955
rect 404780 154924 409889 154952
rect 404780 154912 404786 154924
rect 409877 154921 409889 154924
rect 409923 154921 409935 154955
rect 409877 154915 409935 154921
rect 413646 154912 413652 154964
rect 413704 154952 413710 154964
rect 413848 154952 413876 154992
rect 419442 154980 419448 155032
rect 419500 155020 419506 155032
rect 448790 155020 448796 155032
rect 419500 154992 448796 155020
rect 419500 154980 419506 154992
rect 448790 154980 448796 154992
rect 448848 154980 448854 155032
rect 460906 155020 460934 155128
rect 464614 155116 464620 155168
rect 464672 155156 464678 155168
rect 516042 155156 516048 155168
rect 464672 155128 516048 155156
rect 464672 155116 464678 155128
rect 516042 155116 516048 155128
rect 516100 155116 516106 155168
rect 463326 155048 463332 155100
rect 463384 155088 463390 155100
rect 514110 155088 514116 155100
rect 463384 155060 514116 155088
rect 463384 155048 463390 155060
rect 514110 155048 514116 155060
rect 514168 155048 514174 155100
rect 461486 155020 461492 155032
rect 460906 154992 461492 155020
rect 461486 154980 461492 154992
rect 461544 154980 461550 155032
rect 462038 154980 462044 155032
rect 462096 155020 462102 155032
rect 512178 155020 512184 155032
rect 462096 154992 512184 155020
rect 462096 154980 462102 154992
rect 512178 154980 512184 154992
rect 512236 154980 512242 155032
rect 413704 154924 413876 154952
rect 413704 154912 413710 154924
rect 415210 154912 415216 154964
rect 415268 154952 415274 154964
rect 420825 154955 420883 154961
rect 420825 154952 420837 154955
rect 415268 154924 420837 154952
rect 415268 154912 415274 154924
rect 420825 154921 420837 154924
rect 420871 154921 420883 154955
rect 420825 154915 420883 154921
rect 423030 154912 423036 154964
rect 423088 154952 423094 154964
rect 453666 154952 453672 154964
rect 423088 154924 453672 154952
rect 423088 154912 423094 154924
rect 453666 154912 453672 154924
rect 453724 154912 453730 154964
rect 460106 154912 460112 154964
rect 460164 154952 460170 154964
rect 509234 154952 509240 154964
rect 460164 154924 509240 154952
rect 460164 154912 460170 154924
rect 509234 154912 509240 154924
rect 509292 154912 509298 154964
rect 561674 154912 561680 154964
rect 561732 154952 561738 154964
rect 563790 154952 563796 154964
rect 561732 154924 563796 154952
rect 561732 154912 561738 154924
rect 563790 154912 563796 154924
rect 563848 154912 563854 154964
rect 307067 154856 316264 154884
rect 307067 154853 307079 154856
rect 307021 154847 307079 154853
rect 316586 154844 316592 154896
rect 316644 154884 316650 154896
rect 316644 154856 325694 154884
rect 316644 154844 316650 154856
rect 273254 154816 273260 154828
rect 254912 154788 256464 154816
rect 256620 154788 273260 154816
rect 254912 154776 254918 154788
rect 244277 154751 244335 154757
rect 244277 154748 244289 154751
rect 199344 154720 204944 154748
rect 205008 154720 244289 154748
rect 199344 154708 199350 154720
rect 182784 154652 190454 154680
rect 182784 154640 182790 154652
rect 191466 154640 191472 154692
rect 191524 154680 191530 154692
rect 197541 154683 197599 154689
rect 197541 154680 197553 154683
rect 191524 154652 197553 154680
rect 191524 154640 191530 154652
rect 197541 154649 197553 154652
rect 197587 154649 197599 154683
rect 197541 154643 197599 154649
rect 198274 154640 198280 154692
rect 198332 154680 198338 154692
rect 202969 154683 203027 154689
rect 202969 154680 202981 154683
rect 198332 154652 202981 154680
rect 198332 154640 198338 154652
rect 202969 154649 202981 154652
rect 203015 154649 203027 154683
rect 202969 154643 203027 154649
rect 203061 154683 203119 154689
rect 203061 154649 203073 154683
rect 203107 154680 203119 154683
rect 204901 154683 204959 154689
rect 204901 154680 204913 154683
rect 203107 154652 204913 154680
rect 203107 154649 203119 154652
rect 203061 154643 203119 154649
rect 204901 154649 204913 154652
rect 204947 154649 204959 154683
rect 204901 154643 204959 154649
rect 89162 154572 89168 154624
rect 89220 154612 89226 154624
rect 120166 154612 120172 154624
rect 89220 154584 120172 154612
rect 89220 154572 89226 154584
rect 120166 154572 120172 154584
rect 120224 154572 120230 154624
rect 122282 154572 122288 154624
rect 122340 154612 122346 154624
rect 122340 154584 183508 154612
rect 122340 154572 122346 154584
rect 75454 154504 75460 154556
rect 75512 154544 75518 154556
rect 166905 154547 166963 154553
rect 166905 154544 166917 154547
rect 75512 154516 166917 154544
rect 75512 154504 75518 154516
rect 166905 154513 166917 154516
rect 166951 154513 166963 154547
rect 166905 154507 166963 154513
rect 166994 154504 167000 154556
rect 167052 154544 167058 154556
rect 183002 154544 183008 154556
rect 167052 154516 183008 154544
rect 167052 154504 167058 154516
rect 183002 154504 183008 154516
rect 183060 154504 183066 154556
rect 183480 154544 183508 154584
rect 183646 154572 183652 154624
rect 183704 154612 183710 154624
rect 195241 154615 195299 154621
rect 195241 154612 195253 154615
rect 183704 154584 195253 154612
rect 183704 154572 183710 154584
rect 195241 154581 195253 154584
rect 195287 154581 195299 154615
rect 195241 154575 195299 154581
rect 196342 154572 196348 154624
rect 196400 154612 196406 154624
rect 205008 154612 205036 154720
rect 244277 154717 244289 154720
rect 244323 154717 244335 154751
rect 244277 154711 244335 154717
rect 244553 154751 244611 154757
rect 244553 154717 244565 154751
rect 244599 154748 244611 154751
rect 252649 154751 252707 154757
rect 252649 154748 252661 154751
rect 244599 154720 252661 154748
rect 244599 154717 244611 154720
rect 244553 154711 244611 154717
rect 252649 154717 252661 154720
rect 252695 154717 252707 154751
rect 252649 154711 252707 154717
rect 252833 154751 252891 154757
rect 252833 154717 252845 154751
rect 252879 154748 252891 154751
rect 256513 154751 256571 154757
rect 256513 154748 256525 154751
rect 252879 154720 256525 154748
rect 252879 154717 252891 154720
rect 252833 154711 252891 154717
rect 256513 154717 256525 154720
rect 256559 154717 256571 154751
rect 256513 154711 256571 154717
rect 205177 154683 205235 154689
rect 205177 154649 205189 154683
rect 205223 154680 205235 154683
rect 205913 154683 205971 154689
rect 205913 154680 205925 154683
rect 205223 154652 205925 154680
rect 205223 154649 205235 154652
rect 205177 154643 205235 154649
rect 205913 154649 205925 154652
rect 205959 154649 205971 154683
rect 205913 154643 205971 154649
rect 206094 154640 206100 154692
rect 206152 154680 206158 154692
rect 214561 154683 214619 154689
rect 214561 154680 214573 154683
rect 206152 154652 214573 154680
rect 206152 154640 206158 154652
rect 214561 154649 214573 154652
rect 214607 154649 214619 154683
rect 214561 154643 214619 154649
rect 214653 154683 214711 154689
rect 214653 154649 214665 154683
rect 214699 154680 214711 154683
rect 214699 154652 219572 154680
rect 214699 154649 214711 154652
rect 214653 154643 214711 154649
rect 196400 154584 205036 154612
rect 206005 154615 206063 154621
rect 196400 154572 196406 154584
rect 206005 154581 206017 154615
rect 206051 154612 206063 154615
rect 213825 154615 213883 154621
rect 213825 154612 213837 154615
rect 206051 154584 213837 154612
rect 206051 154581 206063 154584
rect 206005 154575 206063 154581
rect 213825 154581 213837 154584
rect 213871 154581 213883 154615
rect 213825 154575 213883 154581
rect 213914 154572 213920 154624
rect 213972 154612 213978 154624
rect 219250 154612 219256 154624
rect 213972 154584 219256 154612
rect 213972 154572 213978 154584
rect 219250 154572 219256 154584
rect 219308 154572 219314 154624
rect 219345 154615 219403 154621
rect 219345 154581 219357 154615
rect 219391 154612 219403 154615
rect 219437 154615 219495 154621
rect 219437 154612 219449 154615
rect 219391 154584 219449 154612
rect 219391 154581 219403 154584
rect 219345 154575 219403 154581
rect 219437 154581 219449 154584
rect 219483 154581 219495 154615
rect 219544 154612 219572 154652
rect 219618 154640 219624 154692
rect 219676 154680 219682 154692
rect 252554 154680 252560 154692
rect 219676 154652 252560 154680
rect 219676 154640 219682 154652
rect 252554 154640 252560 154652
rect 252612 154640 252618 154692
rect 254765 154683 254823 154689
rect 254765 154649 254777 154683
rect 254811 154680 254823 154683
rect 256620 154680 256648 154788
rect 273254 154776 273260 154788
rect 273312 154776 273318 154828
rect 273346 154776 273352 154828
rect 273404 154816 273410 154828
rect 276109 154819 276167 154825
rect 276109 154816 276121 154819
rect 273404 154788 276121 154816
rect 273404 154776 273410 154788
rect 276109 154785 276121 154788
rect 276155 154785 276167 154819
rect 276109 154779 276167 154785
rect 276201 154819 276259 154825
rect 276201 154785 276213 154819
rect 276247 154816 276259 154819
rect 281997 154819 282055 154825
rect 281997 154816 282009 154819
rect 276247 154788 282009 154816
rect 276247 154785 276259 154788
rect 276201 154779 276259 154785
rect 281997 154785 282009 154788
rect 282043 154785 282055 154819
rect 282273 154819 282331 154825
rect 282273 154816 282285 154819
rect 281997 154779 282055 154785
rect 282104 154788 282285 154816
rect 256697 154751 256755 154757
rect 256697 154717 256709 154751
rect 256743 154748 256755 154751
rect 262858 154748 262864 154760
rect 256743 154720 262864 154748
rect 256743 154717 256755 154720
rect 256697 154711 256755 154717
rect 262858 154708 262864 154720
rect 262916 154708 262922 154760
rect 262953 154751 263011 154757
rect 262953 154717 262965 154751
rect 262999 154748 263011 154751
rect 262999 154720 263732 154748
rect 262999 154717 263011 154720
rect 262953 154711 263011 154717
rect 254811 154652 256648 154680
rect 254811 154649 254823 154652
rect 254765 154643 254823 154649
rect 256786 154640 256792 154692
rect 256844 154680 256850 154692
rect 261297 154683 261355 154689
rect 261297 154680 261309 154683
rect 256844 154652 261309 154680
rect 256844 154640 256850 154652
rect 261297 154649 261309 154652
rect 261343 154649 261355 154683
rect 263594 154680 263600 154692
rect 261297 154643 261355 154649
rect 261404 154652 263600 154680
rect 222102 154612 222108 154624
rect 219544 154584 222108 154612
rect 219437 154575 219495 154581
rect 222102 154572 222108 154584
rect 222160 154572 222166 154624
rect 222654 154572 222660 154624
rect 222712 154612 222718 154624
rect 233881 154615 233939 154621
rect 233881 154612 233893 154615
rect 222712 154584 233893 154612
rect 222712 154572 222718 154584
rect 233881 154581 233893 154584
rect 233927 154581 233939 154615
rect 233881 154575 233939 154581
rect 233973 154615 234031 154621
rect 233973 154581 233985 154615
rect 234019 154612 234031 154615
rect 261404 154612 261432 154652
rect 263594 154640 263600 154652
rect 263652 154640 263658 154692
rect 263704 154680 263732 154720
rect 264606 154708 264612 154760
rect 264664 154748 264670 154760
rect 272521 154751 272579 154757
rect 272521 154748 272533 154751
rect 264664 154720 272533 154748
rect 264664 154708 264670 154720
rect 272521 154717 272533 154720
rect 272567 154717 272579 154751
rect 272521 154711 272579 154717
rect 272613 154751 272671 154757
rect 272613 154717 272625 154751
rect 272659 154748 272671 154751
rect 279326 154748 279332 154760
rect 272659 154720 279332 154748
rect 272659 154717 272671 154720
rect 272613 154711 272671 154717
rect 279326 154708 279332 154720
rect 279384 154708 279390 154760
rect 280065 154751 280123 154757
rect 280065 154717 280077 154751
rect 280111 154748 280123 154751
rect 281813 154751 281871 154757
rect 281813 154748 281825 154751
rect 280111 154720 281825 154748
rect 280111 154717 280123 154720
rect 280065 154711 280123 154717
rect 281813 154717 281825 154720
rect 281859 154717 281871 154751
rect 281813 154711 281871 154717
rect 263704 154652 276060 154680
rect 234019 154584 261432 154612
rect 261481 154615 261539 154621
rect 234019 154581 234031 154584
rect 233973 154575 234031 154581
rect 261481 154581 261493 154615
rect 261527 154612 261539 154615
rect 275922 154612 275928 154624
rect 261527 154584 275928 154612
rect 261527 154581 261539 154584
rect 261481 154575 261539 154581
rect 275922 154572 275928 154584
rect 275980 154572 275986 154624
rect 201494 154544 201500 154556
rect 183480 154516 201500 154544
rect 201494 154504 201500 154516
rect 201552 154504 201558 154556
rect 202782 154504 202788 154556
rect 202840 154544 202846 154556
rect 202840 154516 252508 154544
rect 202840 154504 202846 154516
rect 71590 154436 71596 154488
rect 71648 154476 71654 154488
rect 71648 154448 164004 154476
rect 71648 154436 71654 154448
rect 59906 154368 59912 154420
rect 59964 154408 59970 154420
rect 159634 154408 159640 154420
rect 59964 154380 159640 154408
rect 59964 154368 59970 154380
rect 159634 154368 159640 154380
rect 159692 154368 159698 154420
rect 159729 154411 159787 154417
rect 159729 154377 159741 154411
rect 159775 154408 159787 154411
rect 163777 154411 163835 154417
rect 163777 154408 163789 154411
rect 159775 154380 163789 154408
rect 159775 154377 159787 154380
rect 159729 154371 159787 154377
rect 163777 154377 163789 154380
rect 163823 154377 163835 154411
rect 163777 154371 163835 154377
rect 64782 154300 64788 154352
rect 64840 154340 64846 154352
rect 162854 154340 162860 154352
rect 64840 154312 162860 154340
rect 64840 154300 64846 154312
rect 162854 154300 162860 154312
rect 162912 154300 162918 154352
rect 163976 154340 164004 154448
rect 164050 154436 164056 154488
rect 164108 154476 164114 154488
rect 172606 154476 172612 154488
rect 164108 154448 172612 154476
rect 164108 154436 164114 154448
rect 172606 154436 172612 154448
rect 172664 154436 172670 154488
rect 175918 154436 175924 154488
rect 175976 154476 175982 154488
rect 192754 154476 192760 154488
rect 175976 154448 192760 154476
rect 175976 154436 175982 154448
rect 192754 154436 192760 154448
rect 192812 154436 192818 154488
rect 192846 154436 192852 154488
rect 192904 154476 192910 154488
rect 248046 154476 248052 154488
rect 192904 154448 248052 154476
rect 192904 154436 192910 154448
rect 248046 154436 248052 154448
rect 248104 154436 248110 154488
rect 248785 154479 248843 154485
rect 248785 154445 248797 154479
rect 248831 154476 248843 154479
rect 249978 154476 249984 154488
rect 248831 154448 249984 154476
rect 248831 154445 248843 154448
rect 248785 154439 248843 154445
rect 249978 154436 249984 154448
rect 250036 154436 250042 154488
rect 252480 154476 252508 154516
rect 252554 154504 252560 154556
rect 252612 154544 252618 154556
rect 262398 154544 262404 154556
rect 252612 154516 262404 154544
rect 252612 154504 252618 154516
rect 262398 154504 262404 154516
rect 262456 154504 262462 154556
rect 264974 154504 264980 154556
rect 265032 154544 265038 154556
rect 272794 154544 272800 154556
rect 265032 154516 272800 154544
rect 265032 154504 265038 154516
rect 272794 154504 272800 154516
rect 272852 154504 272858 154556
rect 276032 154544 276060 154652
rect 277210 154640 277216 154692
rect 277268 154680 277274 154692
rect 282104 154680 282132 154788
rect 282273 154785 282285 154788
rect 282319 154785 282331 154819
rect 282273 154779 282331 154785
rect 283098 154776 283104 154828
rect 283156 154816 283162 154828
rect 285769 154819 285827 154825
rect 285769 154816 285781 154819
rect 283156 154788 285781 154816
rect 283156 154776 283162 154788
rect 285769 154785 285781 154788
rect 285815 154785 285827 154819
rect 285769 154779 285827 154785
rect 286042 154776 286048 154828
rect 286100 154816 286106 154828
rect 303433 154819 303491 154825
rect 303433 154816 303445 154819
rect 286100 154788 303445 154816
rect 286100 154776 286106 154788
rect 303433 154785 303445 154788
rect 303479 154785 303491 154819
rect 306558 154816 306564 154828
rect 303433 154779 303491 154785
rect 303540 154788 306564 154816
rect 298002 154748 298008 154760
rect 277268 154652 282132 154680
rect 282196 154720 298008 154748
rect 277268 154640 277274 154652
rect 276109 154615 276167 154621
rect 276109 154581 276121 154615
rect 276155 154612 276167 154615
rect 282196 154612 282224 154720
rect 298002 154708 298008 154720
rect 298060 154708 298066 154760
rect 300581 154751 300639 154757
rect 300581 154717 300593 154751
rect 300627 154748 300639 154751
rect 303540 154748 303568 154788
rect 306558 154776 306564 154788
rect 306616 154776 306622 154828
rect 306929 154819 306987 154825
rect 306929 154785 306941 154819
rect 306975 154816 306987 154819
rect 317322 154816 317328 154828
rect 306975 154788 317328 154816
rect 306975 154785 306987 154788
rect 306929 154779 306987 154785
rect 317322 154776 317328 154788
rect 317380 154776 317386 154828
rect 319073 154819 319131 154825
rect 319073 154785 319085 154819
rect 319119 154816 319131 154819
rect 321738 154816 321744 154828
rect 319119 154788 321744 154816
rect 319119 154785 319131 154788
rect 319073 154779 319131 154785
rect 321738 154776 321744 154788
rect 321796 154776 321802 154828
rect 300627 154720 303568 154748
rect 300627 154717 300639 154720
rect 300581 154711 300639 154717
rect 303614 154708 303620 154760
rect 303672 154748 303678 154760
rect 322198 154748 322204 154760
rect 303672 154720 322204 154748
rect 303672 154708 303678 154720
rect 322198 154708 322204 154720
rect 322256 154708 322262 154760
rect 325666 154748 325694 154856
rect 332778 154844 332784 154896
rect 332836 154884 332842 154896
rect 338666 154884 338672 154896
rect 332836 154856 338672 154884
rect 332836 154844 332842 154856
rect 338666 154844 338672 154856
rect 338724 154844 338730 154896
rect 400950 154844 400956 154896
rect 401008 154884 401014 154896
rect 420546 154884 420552 154896
rect 401008 154856 420552 154884
rect 401008 154844 401014 154856
rect 420546 154844 420552 154856
rect 420604 154844 420610 154896
rect 449802 154884 449808 154896
rect 420656 154856 449808 154884
rect 341610 154776 341616 154828
rect 341668 154816 341674 154828
rect 347498 154816 347504 154828
rect 341668 154788 347504 154816
rect 341668 154776 341674 154788
rect 347498 154776 347504 154788
rect 347556 154776 347562 154828
rect 395982 154776 395988 154828
rect 396040 154816 396046 154828
rect 402241 154819 402299 154825
rect 402241 154816 402253 154819
rect 396040 154788 402253 154816
rect 396040 154776 396046 154788
rect 402241 154785 402253 154788
rect 402287 154785 402299 154819
rect 402241 154779 402299 154785
rect 407022 154776 407028 154828
rect 407080 154816 407086 154828
rect 417421 154819 417479 154825
rect 417421 154816 417433 154819
rect 407080 154788 417433 154816
rect 407080 154776 407086 154788
rect 417421 154785 417433 154788
rect 417467 154785 417479 154819
rect 417421 154779 417479 154785
rect 420454 154776 420460 154828
rect 420512 154816 420518 154828
rect 420656 154816 420684 154856
rect 449802 154844 449808 154856
rect 449860 154844 449866 154896
rect 459462 154844 459468 154896
rect 459520 154884 459526 154896
rect 508222 154884 508228 154896
rect 459520 154856 508228 154884
rect 459520 154844 459526 154856
rect 508222 154844 508228 154856
rect 508280 154844 508286 154896
rect 445846 154816 445852 154828
rect 420512 154788 420684 154816
rect 420748 154788 445852 154816
rect 420512 154776 420518 154788
rect 325666 154720 328316 154748
rect 282273 154683 282331 154689
rect 282273 154649 282285 154683
rect 282319 154680 282331 154683
rect 289722 154680 289728 154692
rect 282319 154652 289728 154680
rect 282319 154649 282331 154652
rect 282273 154643 282331 154649
rect 289722 154640 289728 154652
rect 289780 154640 289786 154692
rect 289817 154683 289875 154689
rect 289817 154649 289829 154683
rect 289863 154680 289875 154683
rect 299566 154680 299572 154692
rect 289863 154652 299572 154680
rect 289863 154649 289875 154652
rect 289817 154643 289875 154649
rect 299566 154640 299572 154652
rect 299624 154640 299630 154692
rect 299658 154640 299664 154692
rect 299716 154680 299722 154692
rect 307021 154683 307079 154689
rect 307021 154680 307033 154683
rect 299716 154652 307033 154680
rect 299716 154640 299722 154652
rect 307021 154649 307033 154652
rect 307067 154649 307079 154683
rect 307021 154643 307079 154649
rect 307113 154683 307171 154689
rect 307113 154649 307125 154683
rect 307159 154680 307171 154683
rect 307159 154652 317276 154680
rect 307159 154649 307171 154652
rect 307113 154643 307171 154649
rect 276155 154584 282224 154612
rect 276155 154581 276167 154584
rect 276109 154575 276167 154581
rect 282362 154572 282368 154624
rect 282420 154612 282426 154624
rect 285858 154612 285864 154624
rect 282420 154584 285864 154612
rect 282420 154572 282426 154584
rect 285858 154572 285864 154584
rect 285916 154572 285922 154624
rect 287793 154615 287851 154621
rect 287793 154581 287805 154615
rect 287839 154612 287851 154615
rect 288621 154615 288679 154621
rect 287839 154584 288572 154612
rect 287839 154581 287851 154584
rect 287793 154575 287851 154581
rect 288434 154544 288440 154556
rect 276032 154516 288440 154544
rect 288434 154504 288440 154516
rect 288492 154504 288498 154556
rect 288544 154544 288572 154584
rect 288621 154581 288633 154615
rect 288667 154612 288679 154615
rect 291841 154615 291899 154621
rect 288667 154584 291792 154612
rect 288667 154581 288679 154584
rect 288621 154575 288679 154581
rect 291562 154544 291568 154556
rect 288544 154516 291568 154544
rect 291562 154504 291568 154516
rect 291620 154504 291626 154556
rect 291764 154544 291792 154584
rect 291841 154581 291853 154615
rect 291887 154612 291899 154615
rect 304445 154615 304503 154621
rect 291887 154584 301544 154612
rect 291887 154581 291899 154584
rect 291841 154575 291899 154581
rect 293954 154544 293960 154556
rect 291764 154516 293960 154544
rect 293954 154504 293960 154516
rect 294012 154504 294018 154556
rect 301516 154544 301544 154584
rect 304445 154581 304457 154615
rect 304491 154612 304503 154615
rect 305914 154612 305920 154624
rect 304491 154584 305920 154612
rect 304491 154581 304503 154584
rect 304445 154575 304503 154581
rect 305914 154572 305920 154584
rect 305972 154572 305978 154624
rect 306466 154572 306472 154624
rect 306524 154612 306530 154624
rect 317141 154615 317199 154621
rect 317141 154612 317153 154615
rect 306524 154584 317153 154612
rect 306524 154572 306530 154584
rect 317141 154581 317153 154584
rect 317187 154581 317199 154615
rect 317141 154575 317199 154581
rect 309870 154544 309876 154556
rect 301516 154516 309876 154544
rect 309870 154504 309876 154516
rect 309928 154504 309934 154556
rect 253290 154476 253296 154488
rect 252480 154448 253296 154476
rect 253290 154436 253296 154448
rect 253348 154436 253354 154488
rect 255314 154436 255320 154488
rect 255372 154476 255378 154488
rect 267826 154476 267832 154488
rect 255372 154448 267832 154476
rect 255372 154436 255378 154448
rect 267826 154436 267832 154448
rect 267884 154436 267890 154488
rect 268289 154479 268347 154485
rect 268289 154445 268301 154479
rect 268335 154476 268347 154479
rect 271782 154476 271788 154488
rect 268335 154448 271788 154476
rect 268335 154445 268347 154448
rect 268289 154439 268347 154445
rect 271782 154436 271788 154448
rect 271840 154436 271846 154488
rect 272429 154479 272487 154485
rect 272429 154445 272441 154479
rect 272475 154476 272487 154479
rect 273346 154476 273352 154488
rect 272475 154448 273352 154476
rect 272475 154445 272487 154448
rect 272429 154439 272487 154445
rect 273346 154436 273352 154448
rect 273404 154436 273410 154488
rect 279326 154436 279332 154488
rect 279384 154476 279390 154488
rect 293586 154476 293592 154488
rect 279384 154448 293592 154476
rect 279384 154436 279390 154448
rect 293586 154436 293592 154448
rect 293644 154436 293650 154488
rect 296901 154479 296959 154485
rect 296901 154445 296913 154479
rect 296947 154476 296959 154479
rect 304626 154476 304632 154488
rect 296947 154448 304632 154476
rect 296947 154445 296959 154448
rect 296901 154439 296959 154445
rect 304626 154436 304632 154448
rect 304684 154436 304690 154488
rect 317248 154476 317276 154652
rect 318150 154640 318156 154692
rect 318208 154680 318214 154692
rect 318208 154652 328224 154680
rect 318208 154640 318214 154652
rect 317417 154615 317475 154621
rect 317417 154581 317429 154615
rect 317463 154612 317475 154615
rect 317463 154584 320128 154612
rect 317463 154581 317475 154584
rect 317417 154575 317475 154581
rect 320100 154544 320128 154584
rect 324314 154544 324320 154556
rect 320100 154516 324320 154544
rect 324314 154504 324320 154516
rect 324372 154504 324378 154556
rect 320910 154476 320916 154488
rect 317248 154448 320916 154476
rect 320910 154436 320916 154448
rect 320968 154436 320974 154488
rect 328196 154476 328224 154652
rect 328288 154544 328316 154720
rect 340598 154708 340604 154760
rect 340656 154748 340662 154760
rect 340656 154720 346440 154748
rect 340656 154708 340662 154720
rect 339678 154640 339684 154692
rect 339736 154680 339742 154692
rect 346302 154680 346308 154692
rect 339736 154652 346308 154680
rect 339736 154640 339742 154652
rect 346302 154640 346308 154652
rect 346360 154640 346366 154692
rect 336734 154572 336740 154624
rect 336792 154612 336798 154624
rect 336792 154584 343588 154612
rect 336792 154572 336798 154584
rect 330662 154544 330668 154556
rect 328288 154516 330668 154544
rect 330662 154504 330668 154516
rect 330720 154504 330726 154556
rect 343560 154544 343588 154584
rect 344370 154544 344376 154556
rect 343560 154516 344376 154544
rect 344370 154504 344376 154516
rect 344428 154504 344434 154556
rect 346412 154544 346440 154720
rect 406746 154708 406752 154760
rect 406804 154748 406810 154760
rect 417329 154751 417387 154757
rect 417329 154748 417341 154751
rect 406804 154720 417341 154748
rect 406804 154708 406810 154720
rect 417329 154717 417341 154720
rect 417375 154717 417387 154751
rect 417329 154711 417387 154717
rect 417786 154708 417792 154760
rect 417844 154748 417850 154760
rect 420748 154748 420776 154788
rect 445846 154776 445852 154788
rect 445904 154776 445910 154828
rect 460658 154776 460664 154828
rect 460716 154816 460722 154828
rect 510246 154816 510252 154828
rect 460716 154788 510252 154816
rect 460716 154776 460722 154788
rect 510246 154776 510252 154788
rect 510304 154776 510310 154828
rect 417844 154720 420776 154748
rect 420825 154751 420883 154757
rect 417844 154708 417850 154720
rect 420825 154717 420837 154751
rect 420871 154748 420883 154751
rect 441982 154748 441988 154760
rect 420871 154720 441988 154748
rect 420871 154717 420883 154720
rect 420825 154711 420883 154717
rect 441982 154708 441988 154720
rect 442040 154708 442046 154760
rect 457530 154708 457536 154760
rect 457588 154748 457594 154760
rect 505370 154748 505376 154760
rect 457588 154720 505376 154748
rect 457588 154708 457594 154720
rect 505370 154708 505376 154720
rect 505428 154708 505434 154760
rect 352282 154640 352288 154692
rect 352340 154680 352346 154692
rect 353386 154680 353392 154692
rect 352340 154652 353392 154680
rect 352340 154640 352346 154652
rect 353386 154640 353392 154652
rect 353444 154640 353450 154692
rect 409414 154640 409420 154692
rect 409472 154680 409478 154692
rect 433242 154680 433248 154692
rect 409472 154652 433248 154680
rect 409472 154640 409478 154652
rect 433242 154640 433248 154652
rect 433300 154640 433306 154692
rect 433337 154683 433395 154689
rect 433337 154649 433349 154683
rect 433383 154680 433395 154683
rect 468294 154680 468300 154692
rect 433383 154652 468300 154680
rect 433383 154649 433395 154652
rect 433337 154643 433395 154649
rect 468294 154640 468300 154652
rect 468352 154640 468358 154692
rect 511166 154680 511172 154692
rect 470566 154652 511172 154680
rect 346486 154572 346492 154624
rect 346544 154612 346550 154624
rect 346544 154584 348372 154612
rect 346544 154572 346550 154584
rect 347038 154544 347044 154556
rect 346412 154516 347044 154544
rect 347038 154504 347044 154516
rect 347096 154504 347102 154556
rect 331950 154476 331956 154488
rect 328196 154448 331956 154476
rect 331950 154436 331956 154448
rect 332008 154436 332014 154488
rect 340966 154436 340972 154488
rect 341024 154476 341030 154488
rect 343726 154476 343732 154488
rect 341024 154448 343732 154476
rect 341024 154436 341030 154448
rect 343726 154436 343732 154448
rect 343784 154436 343790 154488
rect 164145 154411 164203 154417
rect 164145 154377 164157 154411
rect 164191 154408 164203 154411
rect 184290 154408 184296 154420
rect 164191 154380 184296 154408
rect 164191 154377 164203 154380
rect 164145 154371 164203 154377
rect 184290 154368 184296 154380
rect 184348 154368 184354 154420
rect 184658 154368 184664 154420
rect 184716 154408 184722 154420
rect 184716 154380 187556 154408
rect 184716 154368 184722 154380
rect 167454 154340 167460 154352
rect 163976 154312 167460 154340
rect 167454 154300 167460 154312
rect 167512 154300 167518 154352
rect 168101 154343 168159 154349
rect 168101 154309 168113 154343
rect 168147 154340 168159 154343
rect 169665 154343 169723 154349
rect 169665 154340 169677 154343
rect 168147 154312 169677 154340
rect 168147 154309 168159 154312
rect 168101 154303 168159 154309
rect 169665 154309 169677 154312
rect 169711 154309 169723 154343
rect 169665 154303 169723 154309
rect 169754 154300 169760 154352
rect 169812 154340 169818 154352
rect 184934 154340 184940 154352
rect 169812 154312 184940 154340
rect 169812 154300 169818 154312
rect 184934 154300 184940 154312
rect 184992 154300 184998 154352
rect 187528 154340 187556 154380
rect 188522 154368 188528 154420
rect 188580 154408 188586 154420
rect 245654 154408 245660 154420
rect 188580 154380 245660 154408
rect 188580 154368 188586 154380
rect 245654 154368 245660 154380
rect 245712 154368 245718 154420
rect 249058 154368 249064 154420
rect 249116 154408 249122 154420
rect 261110 154408 261116 154420
rect 249116 154380 261116 154408
rect 249116 154368 249122 154380
rect 261110 154368 261116 154380
rect 261168 154368 261174 154420
rect 262674 154368 262680 154420
rect 262732 154408 262738 154420
rect 294874 154408 294880 154420
rect 262732 154380 294880 154408
rect 262732 154368 262738 154380
rect 294874 154368 294880 154380
rect 294932 154368 294938 154420
rect 301409 154411 301467 154417
rect 301409 154377 301421 154411
rect 301455 154408 301467 154411
rect 303614 154408 303620 154420
rect 301455 154380 303620 154408
rect 301455 154377 301467 154380
rect 301409 154371 301467 154377
rect 303614 154368 303620 154380
rect 303672 154368 303678 154420
rect 242894 154340 242900 154352
rect 187528 154312 242900 154340
rect 242894 154300 242900 154312
rect 242952 154300 242958 154352
rect 243170 154300 243176 154352
rect 243228 154340 243234 154352
rect 281902 154340 281908 154352
rect 243228 154312 281908 154340
rect 243228 154300 243234 154312
rect 281902 154300 281908 154312
rect 281960 154300 281966 154352
rect 291102 154300 291108 154352
rect 291160 154340 291166 154352
rect 303982 154340 303988 154352
rect 291160 154312 303988 154340
rect 291160 154300 291166 154312
rect 303982 154300 303988 154312
rect 304040 154300 304046 154352
rect 53098 154232 53104 154284
rect 53156 154272 53162 154284
rect 155034 154272 155040 154284
rect 53156 154244 155040 154272
rect 53156 154232 53162 154244
rect 155034 154232 155040 154244
rect 155092 154232 155098 154284
rect 155862 154232 155868 154284
rect 155920 154272 155926 154284
rect 159729 154275 159787 154281
rect 159729 154272 159741 154275
rect 155920 154244 159741 154272
rect 155920 154232 155926 154244
rect 159729 154241 159741 154244
rect 159775 154241 159787 154275
rect 159729 154235 159787 154241
rect 162762 154232 162768 154284
rect 162820 154272 162826 154284
rect 177206 154272 177212 154284
rect 162820 154244 177212 154272
rect 162820 154232 162826 154244
rect 177206 154232 177212 154244
rect 177264 154232 177270 154284
rect 177942 154232 177948 154284
rect 178000 154272 178006 154284
rect 237650 154272 237656 154284
rect 178000 154244 237656 154272
rect 178000 154232 178006 154244
rect 237650 154232 237656 154244
rect 237708 154232 237714 154284
rect 239214 154232 239220 154284
rect 239272 154272 239278 154284
rect 279326 154272 279332 154284
rect 239272 154244 279332 154272
rect 239272 154232 239278 154244
rect 279326 154232 279332 154244
rect 279384 154232 279390 154284
rect 281813 154275 281871 154281
rect 281813 154241 281825 154275
rect 281859 154272 281871 154275
rect 284478 154272 284484 154284
rect 281859 154244 284484 154272
rect 281859 154241 281871 154244
rect 281813 154235 281871 154241
rect 284478 154232 284484 154244
rect 284536 154232 284542 154284
rect 285674 154232 285680 154284
rect 285732 154272 285738 154284
rect 301406 154272 301412 154284
rect 285732 154244 301412 154272
rect 285732 154232 285738 154244
rect 301406 154232 301412 154244
rect 301464 154232 301470 154284
rect 306282 154232 306288 154284
rect 306340 154272 306346 154284
rect 315022 154272 315028 154284
rect 306340 154244 315028 154272
rect 306340 154232 306346 154244
rect 315022 154232 315028 154244
rect 315080 154232 315086 154284
rect 348344 154272 348372 154584
rect 348418 154572 348424 154624
rect 348476 154612 348482 154624
rect 348476 154584 349292 154612
rect 348476 154572 348482 154584
rect 349264 154340 349292 154584
rect 349338 154572 349344 154624
rect 349396 154612 349402 154624
rect 349396 154584 350304 154612
rect 349396 154572 349402 154584
rect 350276 154544 350304 154584
rect 350350 154572 350356 154624
rect 350408 154612 350414 154624
rect 350408 154584 351316 154612
rect 350408 154572 350414 154584
rect 350276 154516 351224 154544
rect 351196 154408 351224 154516
rect 351288 154476 351316 154584
rect 351362 154572 351368 154624
rect 351420 154612 351426 154624
rect 367922 154612 367928 154624
rect 351420 154584 353248 154612
rect 351420 154572 351426 154584
rect 353220 154544 353248 154584
rect 365732 154584 367928 154612
rect 354122 154544 354128 154556
rect 353220 154516 354128 154544
rect 354122 154504 354128 154516
rect 354180 154504 354186 154556
rect 361482 154504 361488 154556
rect 361540 154544 361546 154556
rect 362034 154544 362040 154556
rect 361540 154516 362040 154544
rect 361540 154504 361546 154516
rect 362034 154504 362040 154516
rect 362092 154504 362098 154556
rect 362586 154504 362592 154556
rect 362644 154544 362650 154556
rect 363046 154544 363052 154556
rect 362644 154516 363052 154544
rect 362644 154504 362650 154516
rect 363046 154504 363052 154516
rect 363104 154504 363110 154556
rect 365622 154504 365628 154556
rect 365680 154544 365686 154556
rect 365732 154544 365760 154584
rect 367922 154572 367928 154584
rect 367980 154572 367986 154624
rect 368842 154612 368848 154624
rect 368032 154584 368848 154612
rect 365680 154516 365760 154544
rect 365680 154504 365686 154516
rect 366450 154504 366456 154556
rect 366508 154544 366514 154556
rect 368032 154544 368060 154584
rect 368842 154572 368848 154584
rect 368900 154572 368906 154624
rect 370866 154612 370872 154624
rect 369964 154584 370872 154612
rect 366508 154516 368060 154544
rect 366508 154504 366514 154516
rect 353478 154476 353484 154488
rect 351288 154448 353484 154476
rect 353478 154436 353484 154448
rect 353536 154436 353542 154488
rect 362862 154436 362868 154488
rect 362920 154476 362926 154488
rect 363966 154476 363972 154488
rect 362920 154448 363972 154476
rect 362920 154436 362926 154448
rect 363966 154436 363972 154448
rect 364024 154436 364030 154488
rect 367002 154436 367008 154488
rect 367060 154476 367066 154488
rect 369854 154476 369860 154488
rect 367060 154448 369860 154476
rect 367060 154436 367066 154448
rect 369854 154436 369860 154448
rect 369912 154436 369918 154488
rect 352834 154408 352840 154420
rect 351196 154380 352840 154408
rect 352834 154368 352840 154380
rect 352892 154368 352898 154420
rect 367738 154368 367744 154420
rect 367796 154408 367802 154420
rect 369964 154408 369992 154584
rect 370866 154572 370872 154584
rect 370924 154572 370930 154624
rect 381538 154612 381544 154624
rect 379532 154584 381544 154612
rect 374914 154504 374920 154556
rect 374972 154544 374978 154556
rect 379532 154544 379560 154584
rect 381538 154572 381544 154584
rect 381596 154572 381602 154624
rect 383470 154612 383476 154624
rect 381648 154584 383476 154612
rect 374972 154516 379560 154544
rect 374972 154504 374978 154516
rect 375190 154436 375196 154488
rect 375248 154476 375254 154488
rect 379606 154476 379612 154488
rect 375248 154448 379612 154476
rect 375248 154436 375254 154448
rect 379606 154436 379612 154448
rect 379664 154436 379670 154488
rect 367796 154380 369992 154408
rect 367796 154368 367802 154380
rect 376202 154368 376208 154420
rect 376260 154408 376266 154420
rect 381648 154408 381676 154584
rect 383470 154572 383476 154584
rect 383528 154572 383534 154624
rect 401042 154612 401048 154624
rect 398852 154584 401048 154612
rect 387702 154504 387708 154556
rect 387760 154544 387766 154556
rect 398852 154544 398880 154584
rect 401042 154572 401048 154584
rect 401100 154572 401106 154624
rect 414566 154572 414572 154624
rect 414624 154612 414630 154624
rect 440970 154612 440976 154624
rect 414624 154584 440976 154612
rect 414624 154572 414630 154584
rect 440970 154572 440976 154584
rect 441028 154572 441034 154624
rect 470566 154612 470594 154652
rect 511166 154640 511172 154652
rect 511224 154640 511230 154692
rect 467852 154584 470594 154612
rect 387760 154516 398880 154544
rect 387760 154504 387766 154516
rect 410702 154504 410708 154556
rect 410760 154544 410766 154556
rect 435174 154544 435180 154556
rect 410760 154516 435180 154544
rect 410760 154504 410766 154516
rect 435174 154504 435180 154516
rect 435232 154504 435238 154556
rect 461394 154504 461400 154556
rect 461452 154544 461458 154556
rect 467852 154544 467880 154584
rect 500126 154572 500132 154624
rect 500184 154612 500190 154624
rect 503346 154612 503352 154624
rect 500184 154584 503352 154612
rect 500184 154572 500190 154584
rect 503346 154572 503352 154584
rect 503404 154572 503410 154624
rect 461452 154516 467880 154544
rect 461452 154504 461458 154516
rect 471790 154504 471796 154556
rect 471848 154544 471854 154556
rect 526806 154544 526812 154556
rect 471848 154516 526812 154544
rect 471848 154504 471854 154516
rect 526806 154504 526812 154516
rect 526864 154504 526870 154556
rect 390462 154436 390468 154488
rect 390520 154476 390526 154488
rect 401594 154476 401600 154488
rect 390520 154448 401600 154476
rect 390520 154436 390526 154448
rect 401594 154436 401600 154448
rect 401652 154436 401658 154488
rect 408310 154436 408316 154488
rect 408368 154476 408374 154488
rect 432230 154476 432236 154488
rect 408368 154448 432236 154476
rect 408368 154436 408374 154448
rect 432230 154436 432236 154448
rect 432288 154436 432294 154488
rect 432598 154436 432604 154488
rect 432656 154476 432662 154488
rect 433337 154479 433395 154485
rect 433337 154476 433349 154479
rect 432656 154448 433349 154476
rect 432656 154436 432662 154448
rect 433337 154445 433349 154448
rect 433383 154445 433395 154479
rect 433337 154439 433395 154445
rect 480898 154436 480904 154488
rect 480956 154476 480962 154488
rect 484946 154476 484952 154488
rect 480956 154448 484952 154476
rect 480956 154436 480962 154448
rect 484946 154436 484952 154448
rect 485004 154436 485010 154488
rect 487062 154436 487068 154488
rect 487120 154476 487126 154488
rect 550174 154476 550180 154488
rect 487120 154448 550180 154476
rect 487120 154436 487126 154448
rect 550174 154436 550180 154448
rect 550232 154436 550238 154488
rect 376260 154380 381676 154408
rect 376260 154368 376266 154380
rect 383286 154368 383292 154420
rect 383344 154408 383350 154420
rect 394234 154408 394240 154420
rect 383344 154380 394240 154408
rect 383344 154368 383350 154380
rect 394234 154368 394240 154380
rect 394292 154368 394298 154420
rect 395062 154368 395068 154420
rect 395120 154408 395126 154420
rect 395525 154411 395583 154417
rect 395120 154380 395476 154408
rect 395120 154368 395126 154380
rect 352098 154340 352104 154352
rect 349264 154312 352104 154340
rect 352098 154300 352104 154312
rect 352156 154300 352162 154352
rect 368382 154300 368388 154352
rect 368440 154340 368446 154352
rect 371786 154340 371792 154352
rect 368440 154312 371792 154340
rect 368440 154300 368446 154312
rect 371786 154300 371792 154312
rect 371844 154300 371850 154352
rect 384022 154300 384028 154352
rect 384080 154340 384086 154352
rect 395154 154340 395160 154352
rect 384080 154312 395160 154340
rect 384080 154300 384086 154312
rect 395154 154300 395160 154312
rect 395212 154300 395218 154352
rect 395448 154340 395476 154380
rect 395525 154377 395537 154411
rect 395571 154408 395583 154411
rect 410794 154408 410800 154420
rect 395571 154380 410800 154408
rect 395571 154377 395583 154380
rect 395525 154371 395583 154377
rect 410794 154368 410800 154380
rect 410852 154368 410858 154420
rect 413922 154368 413928 154420
rect 413980 154408 413986 154420
rect 440050 154408 440056 154420
rect 413980 154380 440056 154408
rect 413980 154368 413986 154380
rect 440050 154368 440056 154380
rect 440108 154368 440114 154420
rect 491202 154368 491208 154420
rect 491260 154408 491266 154420
rect 556062 154408 556068 154420
rect 491260 154380 556068 154408
rect 491260 154368 491266 154380
rect 556062 154368 556068 154380
rect 556120 154368 556126 154420
rect 411806 154340 411812 154352
rect 395448 154312 411812 154340
rect 411806 154300 411812 154312
rect 411864 154300 411870 154352
rect 413278 154300 413284 154352
rect 413336 154340 413342 154352
rect 439038 154340 439044 154352
rect 413336 154312 439044 154340
rect 413336 154300 413342 154312
rect 439038 154300 439044 154312
rect 439096 154300 439102 154352
rect 493962 154300 493968 154352
rect 494020 154340 494026 154352
rect 559926 154340 559932 154352
rect 494020 154312 559932 154340
rect 494020 154300 494026 154312
rect 559926 154300 559932 154312
rect 559984 154300 559990 154352
rect 350810 154272 350816 154284
rect 348344 154244 350816 154272
rect 350810 154232 350816 154244
rect 350868 154232 350874 154284
rect 369670 154232 369676 154284
rect 369728 154272 369734 154284
rect 373718 154272 373724 154284
rect 369728 154244 373724 154272
rect 369728 154232 369734 154244
rect 373718 154232 373724 154244
rect 373776 154232 373782 154284
rect 381446 154232 381452 154284
rect 381504 154272 381510 154284
rect 386782 154272 386788 154284
rect 381504 154244 386788 154272
rect 381504 154232 381510 154244
rect 386782 154232 386788 154244
rect 386840 154232 386846 154284
rect 393038 154232 393044 154284
rect 393096 154272 393102 154284
rect 408862 154272 408868 154284
rect 393096 154244 408868 154272
rect 393096 154232 393102 154244
rect 408862 154232 408868 154244
rect 408920 154232 408926 154284
rect 494606 154232 494612 154284
rect 494664 154272 494670 154284
rect 560938 154272 560944 154284
rect 494664 154244 560944 154272
rect 494664 154232 494670 154244
rect 560938 154232 560944 154244
rect 560996 154232 561002 154284
rect 48222 154164 48228 154216
rect 48280 154204 48286 154216
rect 48280 154176 151814 154204
rect 48280 154164 48286 154176
rect 36538 154096 36544 154148
rect 36596 154136 36602 154148
rect 36596 154108 137324 154136
rect 36596 154096 36602 154108
rect 24762 154028 24768 154080
rect 24820 154068 24826 154080
rect 136174 154068 136180 154080
rect 24820 154040 136180 154068
rect 24820 154028 24826 154040
rect 136174 154028 136180 154040
rect 136232 154028 136238 154080
rect 137189 154071 137247 154077
rect 137189 154068 137201 154071
rect 136468 154040 137201 154068
rect 20898 153960 20904 154012
rect 20956 154000 20962 154012
rect 133874 154000 133880 154012
rect 20956 153972 133880 154000
rect 20956 153960 20962 153972
rect 133874 153960 133880 153972
rect 133932 153960 133938 154012
rect 135162 153960 135168 154012
rect 135220 154000 135226 154012
rect 136468 154000 136496 154040
rect 137189 154037 137201 154040
rect 137235 154037 137247 154071
rect 137189 154031 137247 154037
rect 135220 153972 136496 154000
rect 135220 153960 135226 153972
rect 136542 153960 136548 154012
rect 136600 154000 136606 154012
rect 137296 154000 137324 154108
rect 137830 154096 137836 154148
rect 137888 154136 137894 154148
rect 140777 154139 140835 154145
rect 140777 154136 140789 154139
rect 137888 154108 140789 154136
rect 137888 154096 137894 154108
rect 140777 154105 140789 154108
rect 140823 154105 140835 154139
rect 140777 154099 140835 154105
rect 140866 154096 140872 154148
rect 140924 154136 140930 154148
rect 144733 154139 144791 154145
rect 144733 154136 144745 154139
rect 140924 154108 144745 154136
rect 140924 154096 140930 154108
rect 144733 154105 144745 154108
rect 144779 154105 144791 154139
rect 144733 154099 144791 154105
rect 144822 154096 144828 154148
rect 144880 154136 144886 154148
rect 147125 154139 147183 154145
rect 144880 154108 147076 154136
rect 144880 154096 144886 154108
rect 137465 154071 137523 154077
rect 137465 154037 137477 154071
rect 137511 154068 137523 154071
rect 140958 154068 140964 154080
rect 137511 154040 140964 154068
rect 137511 154037 137523 154040
rect 137465 154031 137523 154037
rect 140958 154028 140964 154040
rect 141016 154028 141022 154080
rect 141053 154071 141111 154077
rect 141053 154037 141065 154071
rect 141099 154068 141111 154071
rect 146941 154071 146999 154077
rect 146941 154068 146953 154071
rect 141099 154040 146953 154068
rect 141099 154037 141111 154040
rect 141053 154031 141111 154037
rect 146941 154037 146953 154040
rect 146987 154037 146999 154071
rect 147048 154068 147076 154108
rect 147125 154105 147137 154139
rect 147171 154136 147183 154139
rect 149333 154139 149391 154145
rect 149333 154136 149345 154139
rect 147171 154108 149345 154136
rect 147171 154105 147183 154108
rect 147125 154099 147183 154105
rect 149333 154105 149345 154108
rect 149379 154105 149391 154139
rect 151786 154136 151814 154176
rect 156506 154164 156512 154216
rect 156564 154204 156570 154216
rect 166261 154207 166319 154213
rect 166261 154204 166273 154207
rect 156564 154176 166273 154204
rect 156564 154164 156570 154176
rect 166261 154173 166273 154176
rect 166307 154173 166319 154207
rect 166261 154167 166319 154173
rect 166905 154207 166963 154213
rect 166905 154173 166917 154207
rect 166951 154204 166963 154207
rect 170030 154204 170036 154216
rect 166951 154176 170036 154204
rect 166951 154173 166963 154176
rect 166905 154167 166963 154173
rect 170030 154164 170036 154176
rect 170088 154164 170094 154216
rect 232498 154204 232504 154216
rect 170140 154176 232504 154204
rect 151998 154136 152004 154148
rect 151786 154108 152004 154136
rect 149333 154099 149391 154105
rect 151998 154096 152004 154108
rect 152056 154096 152062 154148
rect 160094 154096 160100 154148
rect 160152 154136 160158 154148
rect 164786 154136 164792 154148
rect 160152 154108 164792 154136
rect 160152 154096 160158 154108
rect 164786 154096 164792 154108
rect 164844 154096 164850 154148
rect 165154 154096 165160 154148
rect 165212 154136 165218 154148
rect 168101 154139 168159 154145
rect 168101 154136 168113 154139
rect 165212 154108 168113 154136
rect 165212 154096 165218 154108
rect 168101 154105 168113 154108
rect 168147 154105 168159 154139
rect 168101 154099 168159 154105
rect 169018 154096 169024 154148
rect 169076 154136 169082 154148
rect 170140 154136 170168 154176
rect 232498 154164 232504 154176
rect 232556 154164 232562 154216
rect 235350 154164 235356 154216
rect 235408 154204 235414 154216
rect 276658 154204 276664 154216
rect 235408 154176 276664 154204
rect 235408 154164 235414 154176
rect 276658 154164 276664 154176
rect 276716 154164 276722 154216
rect 281997 154207 282055 154213
rect 281997 154173 282009 154207
rect 282043 154204 282055 154207
rect 298830 154204 298836 154216
rect 282043 154176 298836 154204
rect 282043 154173 282055 154176
rect 281997 154167 282055 154173
rect 298830 154164 298836 154176
rect 298888 154164 298894 154216
rect 302234 154164 302240 154216
rect 302292 154204 302298 154216
rect 312446 154204 312452 154216
rect 302292 154176 312452 154204
rect 302292 154164 302298 154176
rect 312446 154164 312452 154176
rect 312504 154164 312510 154216
rect 347590 154164 347596 154216
rect 347648 154204 347654 154216
rect 350166 154204 350172 154216
rect 347648 154176 350172 154204
rect 347648 154164 347654 154176
rect 350166 154164 350172 154176
rect 350224 154164 350230 154216
rect 372982 154164 372988 154216
rect 373040 154204 373046 154216
rect 378594 154204 378600 154216
rect 373040 154176 378600 154204
rect 373040 154164 373046 154176
rect 378594 154164 378600 154176
rect 378652 154164 378658 154216
rect 382090 154164 382096 154216
rect 382148 154204 382154 154216
rect 392302 154204 392308 154216
rect 382148 154176 392308 154204
rect 382148 154164 382154 154176
rect 392302 154164 392308 154176
rect 392360 154164 392366 154216
rect 394418 154164 394424 154216
rect 394476 154204 394482 154216
rect 395525 154207 395583 154213
rect 395525 154204 395537 154207
rect 394476 154176 395537 154204
rect 394476 154164 394482 154176
rect 395525 154173 395537 154176
rect 395571 154173 395583 154207
rect 395525 154167 395583 154173
rect 395706 154164 395712 154216
rect 395764 154204 395770 154216
rect 412542 154204 412548 154216
rect 395764 154176 412548 154204
rect 395764 154164 395770 154176
rect 412542 154164 412548 154176
rect 412600 154164 412606 154216
rect 419166 154164 419172 154216
rect 419224 154204 419230 154216
rect 447870 154204 447876 154216
rect 419224 154176 447876 154204
rect 419224 154164 419230 154176
rect 447870 154164 447876 154176
rect 447928 154164 447934 154216
rect 496538 154164 496544 154216
rect 496596 154204 496602 154216
rect 561674 154204 561680 154216
rect 496596 154176 561680 154204
rect 496596 154164 496602 154176
rect 561674 154164 561680 154176
rect 561732 154164 561738 154216
rect 169076 154108 170168 154136
rect 170217 154139 170275 154145
rect 169076 154096 169082 154108
rect 170217 154105 170229 154139
rect 170263 154136 170275 154139
rect 229830 154136 229836 154148
rect 170263 154108 229836 154136
rect 170263 154105 170275 154108
rect 170217 154099 170275 154105
rect 229830 154096 229836 154108
rect 229888 154096 229894 154148
rect 231486 154096 231492 154148
rect 231544 154136 231550 154148
rect 231544 154108 273024 154136
rect 231544 154096 231550 154108
rect 154574 154068 154580 154080
rect 147048 154040 154580 154068
rect 146941 154031 146999 154037
rect 154574 154028 154580 154040
rect 154632 154028 154638 154080
rect 155310 154028 155316 154080
rect 155368 154068 155374 154080
rect 156966 154068 156972 154080
rect 155368 154040 156972 154068
rect 155368 154028 155374 154040
rect 156966 154028 156972 154040
rect 157024 154028 157030 154080
rect 157334 154028 157340 154080
rect 157392 154068 157398 154080
rect 224954 154068 224960 154080
rect 157392 154040 224960 154068
rect 157392 154028 157398 154040
rect 224954 154028 224960 154040
rect 225012 154028 225018 154080
rect 227530 154028 227536 154080
rect 227588 154068 227594 154080
rect 271506 154068 271512 154080
rect 227588 154040 271512 154068
rect 227588 154028 227594 154040
rect 271506 154028 271512 154040
rect 271564 154028 271570 154080
rect 272996 154068 273024 154108
rect 273254 154096 273260 154148
rect 273312 154136 273318 154148
rect 285766 154136 285772 154148
rect 273312 154108 285772 154136
rect 273312 154096 273318 154108
rect 285766 154096 285772 154108
rect 285824 154096 285830 154148
rect 291746 154096 291752 154148
rect 291804 154136 291810 154148
rect 306650 154136 306656 154148
rect 291804 154108 306656 154136
rect 291804 154096 291810 154108
rect 306650 154096 306656 154108
rect 306708 154096 306714 154148
rect 372338 154096 372344 154148
rect 372396 154136 372402 154148
rect 377674 154136 377680 154148
rect 372396 154108 377680 154136
rect 372396 154096 372402 154108
rect 377674 154096 377680 154108
rect 377732 154096 377738 154148
rect 384942 154096 384948 154148
rect 385000 154136 385006 154148
rect 397178 154136 397184 154148
rect 385000 154108 397184 154136
rect 385000 154096 385006 154108
rect 397178 154096 397184 154108
rect 397236 154096 397242 154148
rect 397270 154096 397276 154148
rect 397328 154136 397334 154148
rect 415670 154136 415676 154148
rect 397328 154108 415676 154136
rect 397328 154096 397334 154108
rect 415670 154096 415676 154108
rect 415728 154096 415734 154148
rect 421742 154096 421748 154148
rect 421800 154136 421806 154148
rect 451734 154136 451740 154148
rect 421800 154108 451740 154136
rect 421800 154096 421806 154108
rect 451734 154096 451740 154108
rect 451792 154096 451798 154148
rect 497826 154096 497832 154148
rect 497884 154136 497890 154148
rect 565722 154136 565728 154148
rect 497884 154108 565728 154136
rect 497884 154096 497890 154108
rect 565722 154096 565728 154108
rect 565780 154096 565786 154148
rect 274082 154068 274088 154080
rect 272996 154040 274088 154068
rect 274082 154028 274088 154040
rect 274140 154028 274146 154080
rect 281442 154028 281448 154080
rect 281500 154068 281506 154080
rect 296162 154068 296168 154080
rect 281500 154040 296168 154068
rect 281500 154028 281506 154040
rect 296162 154028 296168 154040
rect 296220 154028 296226 154080
rect 304902 154028 304908 154080
rect 304960 154068 304966 154080
rect 317690 154068 317696 154080
rect 304960 154040 317696 154068
rect 304960 154028 304966 154040
rect 317690 154028 317696 154040
rect 317748 154028 317754 154080
rect 386230 154028 386236 154080
rect 386288 154068 386294 154080
rect 398742 154068 398748 154080
rect 386288 154040 398748 154068
rect 386288 154028 386294 154040
rect 398742 154028 398748 154040
rect 398800 154028 398806 154080
rect 400122 154028 400128 154080
rect 400180 154068 400186 154080
rect 419534 154068 419540 154080
rect 400180 154040 419540 154068
rect 400180 154028 400186 154040
rect 419534 154028 419540 154040
rect 419592 154028 419598 154080
rect 426894 154028 426900 154080
rect 426952 154068 426958 154080
rect 459554 154068 459560 154080
rect 426952 154040 459560 154068
rect 426952 154028 426958 154040
rect 459554 154028 459560 154040
rect 459612 154028 459618 154080
rect 499114 154028 499120 154080
rect 499172 154068 499178 154080
rect 567746 154068 567752 154080
rect 499172 154040 567752 154068
rect 499172 154028 499178 154040
rect 567746 154028 567752 154040
rect 567804 154028 567810 154080
rect 143994 154000 144000 154012
rect 136600 153972 137232 154000
rect 137296 153972 144000 154000
rect 136600 153960 136606 153972
rect 17034 153892 17040 153944
rect 17092 153932 17098 153944
rect 131114 153932 131120 153944
rect 17092 153904 131120 153932
rect 17092 153892 17098 153904
rect 131114 153892 131120 153904
rect 131172 153892 131178 153944
rect 131298 153892 131304 153944
rect 131356 153932 131362 153944
rect 137204 153932 137232 153972
rect 143994 153960 144000 153972
rect 144052 153960 144058 154012
rect 144733 154003 144791 154009
rect 144733 153969 144745 154003
rect 144779 154000 144791 154003
rect 149238 154000 149244 154012
rect 144779 153972 149244 154000
rect 144779 153969 144791 153972
rect 144733 153963 144791 153969
rect 149238 153960 149244 153972
rect 149296 153960 149302 154012
rect 149333 154003 149391 154009
rect 149333 153969 149345 154003
rect 149379 154000 149391 154003
rect 216858 154000 216864 154012
rect 149379 153972 216864 154000
rect 149379 153969 149391 153972
rect 149333 153963 149391 153969
rect 216858 153960 216864 153972
rect 216916 153960 216922 154012
rect 219710 153960 219716 154012
rect 219768 154000 219774 154012
rect 266354 154000 266360 154012
rect 219768 153972 266360 154000
rect 219768 153960 219774 153972
rect 266354 153960 266360 153972
rect 266412 153960 266418 154012
rect 276014 153960 276020 154012
rect 276072 154000 276078 154012
rect 291194 154000 291200 154012
rect 276072 153972 291200 154000
rect 276072 153960 276078 153972
rect 291194 153960 291200 153972
rect 291252 153960 291258 154012
rect 293034 153960 293040 154012
rect 293092 154000 293098 154012
rect 311894 154000 311900 154012
rect 293092 153972 311900 154000
rect 293092 153960 293098 153972
rect 311894 153960 311900 153972
rect 311952 153960 311958 154012
rect 311986 153960 311992 154012
rect 312044 154000 312050 154012
rect 322934 154000 322940 154012
rect 312044 153972 322940 154000
rect 312044 153960 312050 153972
rect 322934 153960 322940 153972
rect 322992 153960 322998 154012
rect 347774 153960 347780 154012
rect 347832 154000 347838 154012
rect 351454 154000 351460 154012
rect 347832 153972 351460 154000
rect 347832 153960 347838 153972
rect 351454 153960 351460 153972
rect 351512 153960 351518 154012
rect 373902 153960 373908 154012
rect 373960 154000 373966 154012
rect 378134 154000 378140 154012
rect 373960 153972 378140 154000
rect 373960 153960 373966 153972
rect 378134 153960 378140 153972
rect 378192 153960 378198 154012
rect 389818 153960 389824 154012
rect 389876 154000 389882 154012
rect 401686 154000 401692 154012
rect 389876 153972 401692 154000
rect 389876 153960 389882 153972
rect 401686 153960 401692 153972
rect 401744 153960 401750 154012
rect 405458 153960 405464 154012
rect 405516 154000 405522 154012
rect 427354 154000 427360 154012
rect 405516 153972 427360 154000
rect 405516 153960 405522 153972
rect 427354 153960 427360 153972
rect 427412 153960 427418 154012
rect 429562 153960 429568 154012
rect 429620 154000 429626 154012
rect 463418 154000 463424 154012
rect 429620 153972 463424 154000
rect 429620 153960 429626 153972
rect 463418 153960 463424 153972
rect 463476 153960 463482 154012
rect 500862 153960 500868 154012
rect 500920 154000 500926 154012
rect 570690 154000 570696 154012
rect 500920 153972 570696 154000
rect 500920 153960 500926 153972
rect 570690 153960 570696 153972
rect 570748 153960 570754 154012
rect 138106 153932 138112 153944
rect 131356 153904 136956 153932
rect 137204 153904 138112 153932
rect 131356 153892 131362 153904
rect 1394 153824 1400 153876
rect 1452 153864 1458 153876
rect 120626 153864 120632 153876
rect 1452 153836 120632 153864
rect 1452 153824 1458 153836
rect 120626 153824 120632 153836
rect 120684 153824 120690 153876
rect 120718 153824 120724 153876
rect 120776 153864 120782 153876
rect 125778 153864 125784 153876
rect 120776 153836 125784 153864
rect 120776 153824 120782 153836
rect 125778 153824 125784 153836
rect 125836 153824 125842 153876
rect 127437 153867 127495 153873
rect 127437 153833 127449 153867
rect 127483 153864 127495 153867
rect 130378 153864 130384 153876
rect 127483 153836 130384 153864
rect 127483 153833 127495 153836
rect 127437 153827 127495 153833
rect 130378 153824 130384 153836
rect 130436 153824 130442 153876
rect 131206 153824 131212 153876
rect 131264 153864 131270 153876
rect 132954 153864 132960 153876
rect 131264 153836 132960 153864
rect 131264 153824 131270 153836
rect 132954 153824 132960 153836
rect 133012 153824 133018 153876
rect 133046 153824 133052 153876
rect 133104 153864 133110 153876
rect 135530 153864 135536 153876
rect 133104 153836 135536 153864
rect 133104 153824 133110 153836
rect 135530 153824 135536 153836
rect 135588 153824 135594 153876
rect 136928 153864 136956 153904
rect 138106 153892 138112 153904
rect 138164 153892 138170 153944
rect 138198 153892 138204 153944
rect 138256 153932 138262 153944
rect 140682 153932 140688 153944
rect 138256 153904 140688 153932
rect 138256 153892 138262 153904
rect 140682 153892 140688 153904
rect 140740 153892 140746 153944
rect 140774 153892 140780 153944
rect 140832 153932 140838 153944
rect 143534 153932 143540 153944
rect 140832 153904 143540 153932
rect 140832 153892 140838 153904
rect 143534 153892 143540 153904
rect 143592 153892 143598 153944
rect 143626 153892 143632 153944
rect 143684 153932 143690 153944
rect 146570 153932 146576 153944
rect 143684 153904 146576 153932
rect 143684 153892 143690 153904
rect 146570 153892 146576 153904
rect 146628 153892 146634 153944
rect 146941 153935 146999 153941
rect 146941 153901 146953 153935
rect 146987 153932 146999 153935
rect 211614 153932 211620 153944
rect 146987 153904 211620 153932
rect 146987 153901 146999 153904
rect 146941 153895 146999 153901
rect 211614 153892 211620 153904
rect 211672 153892 211678 153944
rect 215846 153892 215852 153944
rect 215904 153932 215910 153944
rect 215904 153904 258074 153932
rect 215904 153892 215910 153904
rect 203886 153864 203892 153876
rect 136928 153836 203892 153864
rect 203886 153824 203892 153836
rect 203944 153824 203950 153876
rect 204162 153824 204168 153876
rect 204220 153864 204226 153876
rect 255866 153864 255872 153876
rect 204220 153836 255872 153864
rect 204220 153824 204226 153836
rect 255866 153824 255872 153836
rect 255924 153824 255930 153876
rect 258046 153864 258074 153904
rect 263594 153892 263600 153944
rect 263652 153932 263658 153944
rect 270494 153932 270500 153944
rect 263652 153904 270500 153932
rect 263652 153892 263658 153904
rect 270494 153892 270500 153904
rect 270552 153892 270558 153944
rect 278222 153892 278228 153944
rect 278280 153932 278286 153944
rect 305270 153932 305276 153944
rect 278280 153904 305276 153932
rect 278280 153892 278286 153904
rect 305270 153892 305276 153904
rect 305328 153892 305334 153944
rect 309134 153892 309140 153944
rect 309192 153932 309198 153944
rect 320266 153932 320272 153944
rect 309192 153904 320272 153932
rect 309192 153892 309198 153904
rect 320266 153892 320272 153904
rect 320324 153892 320330 153944
rect 334434 153892 334440 153944
rect 334492 153932 334498 153944
rect 339126 153932 339132 153944
rect 334492 153904 339132 153932
rect 334492 153892 334498 153904
rect 339126 153892 339132 153904
rect 339184 153892 339190 153944
rect 376478 153892 376484 153944
rect 376536 153932 376542 153944
rect 380894 153932 380900 153944
rect 376536 153904 380900 153932
rect 376536 153892 376542 153904
rect 380894 153892 380900 153904
rect 380952 153892 380958 153944
rect 382734 153892 382740 153944
rect 382792 153932 382798 153944
rect 388162 153932 388168 153944
rect 382792 153904 388168 153932
rect 382792 153892 382798 153904
rect 388162 153892 388168 153904
rect 388220 153892 388226 153944
rect 391198 153892 391204 153944
rect 391256 153932 391262 153944
rect 404262 153932 404268 153944
rect 391256 153904 404268 153932
rect 391256 153892 391262 153904
rect 404262 153892 404268 153904
rect 404320 153892 404326 153944
rect 408034 153892 408040 153944
rect 408092 153932 408098 153944
rect 431218 153932 431224 153944
rect 408092 153904 431224 153932
rect 408092 153892 408098 153904
rect 431218 153892 431224 153904
rect 431276 153892 431282 153944
rect 431770 153892 431776 153944
rect 431828 153932 431834 153944
rect 467282 153932 467288 153944
rect 431828 153904 467288 153932
rect 431828 153892 431834 153904
rect 467282 153892 467288 153904
rect 467340 153892 467346 153944
rect 503070 153892 503076 153944
rect 503128 153932 503134 153944
rect 573542 153932 573548 153944
rect 503128 153904 573548 153932
rect 503128 153892 503134 153904
rect 573542 153892 573548 153904
rect 573600 153892 573606 153944
rect 263686 153864 263692 153876
rect 258046 153836 263692 153864
rect 263686 153824 263692 153836
rect 263744 153824 263750 153876
rect 292574 153864 292580 153876
rect 267706 153836 292580 153864
rect 83274 153756 83280 153808
rect 83332 153796 83338 153808
rect 175274 153796 175280 153808
rect 83332 153768 175280 153796
rect 83332 153756 83338 153768
rect 175274 153756 175280 153768
rect 175332 153756 175338 153808
rect 179414 153756 179420 153808
rect 179472 153796 179478 153808
rect 211154 153796 211160 153808
rect 179472 153768 211160 153796
rect 179472 153756 179478 153768
rect 211154 153756 211160 153768
rect 211212 153756 211218 153808
rect 260558 153756 260564 153808
rect 260616 153796 260622 153808
rect 267706 153796 267734 153836
rect 292574 153824 292580 153836
rect 292632 153824 292638 153876
rect 295794 153824 295800 153876
rect 295852 153864 295858 153876
rect 317046 153864 317052 153876
rect 295852 153836 317052 153864
rect 295852 153824 295858 153836
rect 317046 153824 317052 153836
rect 317104 153824 317110 153876
rect 336458 153824 336464 153876
rect 336516 153864 336522 153876
rect 339770 153864 339776 153876
rect 336516 153836 339776 153864
rect 336516 153824 336522 153836
rect 339770 153824 339776 153836
rect 339828 153824 339834 153876
rect 340782 153824 340788 153876
rect 340840 153864 340846 153876
rect 342990 153864 342996 153876
rect 340840 153836 342996 153864
rect 340840 153824 340846 153836
rect 342990 153824 342996 153836
rect 343048 153824 343054 153876
rect 373626 153824 373632 153876
rect 373684 153864 373690 153876
rect 379422 153864 379428 153876
rect 373684 153836 379428 153864
rect 373684 153824 373690 153836
rect 379422 153824 379428 153836
rect 379480 153824 379486 153876
rect 389082 153824 389088 153876
rect 389140 153864 389146 153876
rect 400214 153864 400220 153876
rect 389140 153836 400220 153864
rect 389140 153824 389146 153836
rect 400214 153824 400220 153836
rect 400272 153824 400278 153876
rect 402698 153824 402704 153876
rect 402756 153864 402762 153876
rect 423490 153864 423496 153876
rect 402756 153836 423496 153864
rect 402756 153824 402762 153836
rect 423490 153824 423496 153836
rect 423548 153824 423554 153876
rect 456242 153824 456248 153876
rect 456300 153864 456306 153876
rect 500126 153864 500132 153876
rect 456300 153836 500132 153864
rect 456300 153824 456306 153836
rect 500126 153824 500132 153836
rect 500184 153824 500190 153876
rect 501690 153824 501696 153876
rect 501748 153864 501754 153876
rect 571610 153864 571616 153876
rect 501748 153836 571616 153864
rect 501748 153824 501754 153836
rect 571610 153824 571616 153836
rect 571668 153824 571674 153876
rect 260616 153768 267734 153796
rect 260616 153756 260622 153768
rect 270402 153756 270408 153808
rect 270460 153796 270466 153808
rect 280614 153796 280620 153808
rect 270460 153768 280620 153796
rect 270460 153756 270466 153768
rect 280614 153756 280620 153768
rect 280672 153756 280678 153808
rect 287054 153756 287060 153808
rect 287112 153796 287118 153808
rect 289078 153796 289084 153808
rect 287112 153768 289084 153796
rect 287112 153756 287118 153768
rect 289078 153756 289084 153768
rect 289136 153756 289142 153808
rect 289998 153756 290004 153808
rect 290056 153796 290062 153808
rect 291654 153796 291660 153808
rect 290056 153768 291660 153796
rect 290056 153756 290062 153768
rect 291654 153756 291660 153768
rect 291712 153756 291718 153808
rect 326798 153756 326804 153808
rect 326856 153796 326862 153808
rect 328086 153796 328092 153808
rect 326856 153768 328092 153796
rect 326856 153756 326862 153768
rect 328086 153756 328092 153768
rect 328144 153756 328150 153808
rect 328178 153756 328184 153808
rect 328236 153796 328242 153808
rect 329374 153796 329380 153808
rect 328236 153768 329380 153796
rect 328236 153756 328242 153768
rect 329374 153756 329380 153768
rect 329432 153756 329438 153808
rect 339402 153756 339408 153808
rect 339460 153796 339466 153808
rect 342346 153796 342352 153808
rect 339460 153768 342352 153796
rect 339460 153756 339466 153768
rect 342346 153756 342352 153768
rect 342404 153756 342410 153808
rect 377490 153756 377496 153808
rect 377548 153796 377554 153808
rect 382366 153796 382372 153808
rect 377548 153768 382372 153796
rect 377548 153756 377554 153768
rect 382366 153756 382372 153768
rect 382424 153756 382430 153808
rect 385770 153756 385776 153808
rect 385828 153796 385834 153808
rect 398098 153796 398104 153808
rect 385828 153768 398104 153796
rect 385828 153756 385834 153768
rect 398098 153756 398104 153768
rect 398156 153756 398162 153808
rect 398282 153756 398288 153808
rect 398340 153796 398346 153808
rect 413830 153796 413836 153808
rect 398340 153768 413836 153796
rect 398340 153756 398346 153768
rect 413830 153756 413836 153768
rect 413888 153756 413894 153808
rect 416498 153756 416504 153808
rect 416556 153796 416562 153808
rect 443914 153796 443920 153808
rect 416556 153768 443920 153796
rect 416556 153756 416562 153768
rect 443914 153756 443920 153768
rect 443972 153756 443978 153808
rect 470318 153756 470324 153808
rect 470376 153796 470382 153808
rect 524874 153796 524880 153808
rect 470376 153768 524880 153796
rect 470376 153756 470382 153768
rect 524874 153756 524880 153768
rect 524932 153756 524938 153808
rect 93026 153688 93032 153740
rect 93084 153728 93090 153740
rect 175921 153731 175979 153737
rect 175921 153728 175933 153731
rect 93084 153700 175933 153728
rect 93084 153688 93090 153700
rect 175921 153697 175933 153700
rect 175967 153697 175979 153731
rect 180426 153728 180432 153740
rect 175921 153691 175979 153697
rect 177960 153700 180432 153728
rect 91094 153620 91100 153672
rect 91152 153660 91158 153672
rect 177960 153660 177988 153700
rect 180426 153688 180432 153700
rect 180484 153688 180490 153740
rect 185578 153688 185584 153740
rect 185636 153728 185642 153740
rect 213914 153728 213920 153740
rect 185636 153700 213920 153728
rect 185636 153688 185642 153700
rect 213914 153688 213920 153700
rect 213972 153688 213978 153740
rect 262214 153688 262220 153740
rect 262272 153728 262278 153740
rect 265618 153728 265624 153740
rect 262272 153700 265624 153728
rect 262272 153688 262278 153700
rect 265618 153688 265624 153700
rect 265676 153688 265682 153740
rect 273346 153688 273352 153740
rect 273404 153728 273410 153740
rect 283190 153728 283196 153740
rect 273404 153700 283196 153728
rect 273404 153688 273410 153700
rect 283190 153688 283196 153700
rect 283248 153688 283254 153740
rect 327074 153688 327080 153740
rect 327132 153728 327138 153740
rect 331306 153728 331312 153740
rect 327132 153700 331312 153728
rect 327132 153688 327138 153700
rect 331306 153688 331312 153700
rect 331364 153688 331370 153740
rect 378778 153688 378784 153740
rect 378836 153728 378842 153740
rect 384206 153728 384212 153740
rect 378836 153700 384212 153728
rect 378836 153688 378842 153700
rect 384206 153688 384212 153700
rect 384264 153688 384270 153740
rect 391842 153688 391848 153740
rect 391900 153728 391906 153740
rect 403434 153728 403440 153740
rect 391900 153700 403440 153728
rect 391900 153688 391906 153700
rect 403434 153688 403440 153700
rect 403492 153688 403498 153740
rect 424318 153688 424324 153740
rect 424376 153728 424382 153740
rect 455598 153728 455604 153740
rect 424376 153700 455604 153728
rect 424376 153688 424382 153700
rect 455598 153688 455604 153700
rect 455656 153688 455662 153740
rect 469122 153688 469128 153740
rect 469180 153728 469186 153740
rect 522850 153728 522856 153740
rect 469180 153700 522856 153728
rect 469180 153688 469186 153700
rect 522850 153688 522856 153700
rect 522908 153688 522914 153740
rect 91152 153632 177988 153660
rect 91152 153620 91158 153632
rect 178034 153620 178040 153672
rect 178092 153660 178098 153672
rect 195422 153660 195428 153672
rect 178092 153632 195428 153660
rect 178092 153620 178098 153632
rect 195422 153620 195428 153632
rect 195480 153620 195486 153672
rect 195514 153620 195520 153672
rect 195572 153660 195578 153672
rect 219618 153660 219624 153672
rect 195572 153632 219624 153660
rect 195572 153620 195578 153632
rect 219618 153620 219624 153632
rect 219676 153620 219682 153672
rect 260926 153620 260932 153672
rect 260984 153660 260990 153672
rect 263042 153660 263048 153672
rect 260984 153632 263048 153660
rect 260984 153620 260990 153632
rect 263042 153620 263048 153632
rect 263100 153620 263106 153672
rect 269390 153620 269396 153672
rect 269448 153660 269454 153672
rect 270862 153660 270868 153672
rect 269448 153632 270868 153660
rect 269448 153620 269454 153632
rect 270862 153620 270868 153632
rect 270920 153620 270926 153672
rect 321738 153620 321744 153672
rect 321796 153660 321802 153672
rect 324961 153663 325019 153669
rect 324961 153660 324973 153663
rect 321796 153632 324973 153660
rect 321796 153620 321802 153632
rect 324961 153629 324973 153632
rect 325007 153629 325019 153663
rect 324961 153623 325019 153629
rect 326706 153620 326712 153672
rect 326764 153660 326770 153672
rect 327442 153660 327448 153672
rect 326764 153632 327448 153660
rect 326764 153620 326770 153632
rect 327442 153620 327448 153632
rect 327500 153620 327506 153672
rect 336550 153620 336556 153672
rect 336608 153660 336614 153672
rect 340414 153660 340420 153672
rect 336608 153632 340420 153660
rect 336608 153620 336614 153632
rect 340414 153620 340420 153632
rect 340472 153620 340478 153672
rect 370958 153620 370964 153672
rect 371016 153660 371022 153672
rect 375742 153660 375748 153672
rect 371016 153632 375748 153660
rect 371016 153620 371022 153632
rect 375742 153620 375748 153632
rect 375800 153620 375806 153672
rect 380066 153620 380072 153672
rect 380124 153660 380130 153672
rect 385862 153660 385868 153672
rect 380124 153632 385868 153660
rect 380124 153620 380130 153632
rect 385862 153620 385868 153632
rect 385920 153620 385926 153672
rect 388530 153620 388536 153672
rect 388588 153660 388594 153672
rect 400306 153660 400312 153672
rect 388588 153632 400312 153660
rect 388588 153620 388594 153632
rect 400306 153620 400312 153632
rect 400364 153620 400370 153672
rect 403526 153620 403532 153672
rect 403584 153660 403590 153672
rect 413646 153660 413652 153672
rect 403584 153632 413652 153660
rect 403584 153620 403590 153632
rect 413646 153620 413652 153632
rect 413704 153620 413710 153672
rect 466178 153620 466184 153672
rect 466236 153660 466242 153672
rect 518986 153660 518992 153672
rect 466236 153632 518992 153660
rect 466236 153620 466242 153632
rect 518986 153620 518992 153632
rect 519044 153620 519050 153672
rect 98914 153552 98920 153604
rect 98972 153592 98978 153604
rect 185670 153592 185676 153604
rect 98972 153564 185676 153592
rect 98972 153552 98978 153564
rect 185670 153552 185676 153564
rect 185728 153552 185734 153604
rect 193122 153552 193128 153604
rect 193180 153592 193186 153604
rect 208394 153592 208400 153604
rect 193180 153564 208400 153592
rect 193180 153552 193186 153564
rect 208394 153552 208400 153564
rect 208452 153552 208458 153604
rect 208486 153552 208492 153604
rect 208544 153592 208550 153604
rect 214282 153592 214288 153604
rect 208544 153564 214288 153592
rect 208544 153552 208550 153564
rect 214282 153552 214288 153564
rect 214340 153552 214346 153604
rect 321646 153552 321652 153604
rect 321704 153592 321710 153604
rect 327074 153592 327080 153604
rect 321704 153564 327080 153592
rect 321704 153552 321710 153564
rect 327074 153552 327080 153564
rect 327132 153552 327138 153604
rect 337930 153552 337936 153604
rect 337988 153592 337994 153604
rect 341058 153592 341064 153604
rect 337988 153564 341064 153592
rect 337988 153552 337994 153564
rect 341058 153552 341064 153564
rect 341116 153552 341122 153604
rect 369026 153552 369032 153604
rect 369084 153592 369090 153604
rect 372798 153592 372804 153604
rect 369084 153564 372804 153592
rect 369084 153552 369090 153564
rect 372798 153552 372804 153564
rect 372856 153552 372862 153604
rect 378042 153552 378048 153604
rect 378100 153592 378106 153604
rect 382274 153592 382280 153604
rect 378100 153564 382280 153592
rect 378100 153552 378106 153564
rect 382274 153552 382280 153564
rect 382332 153552 382338 153604
rect 393774 153552 393780 153604
rect 393832 153592 393838 153604
rect 405918 153592 405924 153604
rect 393832 153564 405924 153592
rect 393832 153552 393838 153564
rect 405918 153552 405924 153564
rect 405976 153552 405982 153604
rect 417142 153552 417148 153604
rect 417200 153592 417206 153604
rect 417970 153592 417976 153604
rect 417200 153564 417976 153592
rect 417200 153552 417206 153564
rect 417970 153552 417976 153564
rect 418028 153552 418034 153604
rect 443822 153552 443828 153604
rect 443880 153592 443886 153604
rect 445662 153592 445668 153604
rect 443880 153564 445668 153592
rect 443880 153552 443886 153564
rect 445662 153552 445668 153564
rect 445720 153552 445726 153604
rect 455230 153552 455236 153604
rect 455288 153592 455294 153604
rect 456702 153592 456708 153604
rect 455288 153564 456708 153592
rect 455288 153552 455294 153564
rect 456702 153552 456708 153564
rect 456760 153552 456766 153604
rect 463602 153552 463608 153604
rect 463660 153592 463666 153604
rect 515122 153592 515128 153604
rect 463660 153564 515128 153592
rect 463660 153552 463666 153564
rect 515122 153552 515128 153564
rect 515180 153552 515186 153604
rect 1302 153484 1308 153536
rect 1360 153524 1366 153536
rect 120074 153524 120080 153536
rect 1360 153496 120080 153524
rect 1360 153484 1366 153496
rect 120074 153484 120080 153496
rect 120132 153484 120138 153536
rect 120169 153527 120227 153533
rect 120169 153493 120181 153527
rect 120215 153524 120227 153527
rect 193398 153524 193404 153536
rect 120215 153496 193404 153524
rect 120215 153493 120227 153496
rect 120169 153487 120227 153493
rect 193398 153484 193404 153496
rect 193456 153484 193462 153536
rect 200114 153484 200120 153536
rect 200172 153524 200178 153536
rect 200574 153524 200580 153536
rect 200172 153496 200580 153524
rect 200172 153484 200178 153496
rect 200574 153484 200580 153496
rect 200632 153484 200638 153536
rect 249794 153484 249800 153536
rect 249852 153524 249858 153536
rect 257154 153524 257160 153536
rect 249852 153496 257160 153524
rect 249852 153484 249858 153496
rect 257154 153484 257160 153496
rect 257212 153484 257218 153536
rect 259362 153484 259368 153536
rect 259420 153524 259426 153536
rect 260466 153524 260472 153536
rect 259420 153496 260472 153524
rect 259420 153484 259426 153496
rect 260466 153484 260472 153496
rect 260524 153484 260530 153536
rect 284294 153484 284300 153536
rect 284352 153524 284358 153536
rect 286410 153524 286416 153536
rect 284352 153496 286416 153524
rect 284352 153484 284358 153496
rect 286410 153484 286416 153496
rect 286468 153484 286474 153536
rect 291562 153484 291568 153536
rect 291620 153524 291626 153536
rect 297542 153524 297548 153536
rect 291620 153496 297548 153524
rect 291620 153484 291626 153496
rect 297542 153484 297548 153496
rect 297600 153484 297606 153536
rect 297910 153484 297916 153536
rect 297968 153524 297974 153536
rect 299474 153524 299480 153536
rect 297968 153496 299480 153524
rect 297968 153484 297974 153496
rect 299474 153484 299480 153496
rect 299532 153484 299538 153536
rect 322842 153484 322848 153536
rect 322900 153524 322906 153536
rect 323486 153524 323492 153536
rect 322900 153496 323492 153524
rect 322900 153484 322906 153496
rect 323486 153484 323492 153496
rect 323544 153484 323550 153536
rect 344186 153484 344192 153536
rect 344244 153524 344250 153536
rect 345658 153524 345664 153536
rect 344244 153496 345664 153524
rect 344244 153484 344250 153496
rect 345658 153484 345664 153496
rect 345716 153484 345722 153536
rect 370314 153484 370320 153536
rect 370372 153524 370378 153536
rect 374730 153524 374736 153536
rect 370372 153496 374736 153524
rect 370372 153484 370378 153496
rect 374730 153484 374736 153496
rect 374788 153484 374794 153536
rect 380710 153484 380716 153536
rect 380768 153524 380774 153536
rect 385954 153524 385960 153536
rect 380768 153496 385960 153524
rect 380768 153484 380774 153496
rect 385954 153484 385960 153496
rect 386012 153484 386018 153536
rect 392486 153484 392492 153536
rect 392544 153524 392550 153536
rect 404814 153524 404820 153536
rect 392544 153496 404820 153524
rect 392544 153484 392550 153496
rect 404814 153484 404820 153496
rect 404872 153484 404878 153536
rect 458082 153484 458088 153536
rect 458140 153524 458146 153536
rect 458140 153496 489914 153524
rect 458140 153484 458146 153496
rect 108301 153459 108359 153465
rect 108301 153425 108313 153459
rect 108347 153456 108359 153459
rect 113545 153459 113603 153465
rect 113545 153456 113557 153459
rect 108347 153428 113557 153456
rect 108347 153425 108359 153428
rect 108301 153419 108359 153425
rect 113545 153425 113557 153428
rect 113591 153425 113603 153459
rect 113545 153419 113603 153425
rect 113637 153459 113695 153465
rect 113637 153425 113649 153459
rect 113683 153456 113695 153459
rect 171962 153456 171968 153468
rect 113683 153428 171968 153456
rect 113683 153425 113695 153428
rect 113637 153419 113695 153425
rect 171962 153416 171968 153428
rect 172020 153416 172026 153468
rect 175921 153459 175979 153465
rect 175921 153425 175933 153459
rect 175967 153456 175979 153459
rect 181714 153456 181720 153468
rect 175967 153428 181720 153456
rect 175967 153425 175979 153428
rect 175921 153419 175979 153425
rect 181714 153416 181720 153428
rect 181772 153416 181778 153468
rect 182082 153416 182088 153468
rect 182140 153456 182146 153468
rect 198734 153456 198740 153468
rect 182140 153428 198740 153456
rect 182140 153416 182146 153428
rect 198734 153416 198740 153428
rect 198792 153416 198798 153468
rect 271782 153416 271788 153468
rect 271840 153456 271846 153468
rect 277946 153456 277952 153468
rect 271840 153428 277952 153456
rect 271840 153416 271846 153428
rect 277946 153416 277952 153428
rect 278004 153416 278010 153468
rect 299566 153416 299572 153468
rect 299624 153456 299630 153468
rect 307294 153456 307300 153468
rect 299624 153428 307300 153456
rect 299624 153416 299630 153428
rect 307294 153416 307300 153428
rect 307352 153416 307358 153468
rect 320082 153416 320088 153468
rect 320140 153456 320146 153468
rect 324866 153456 324872 153468
rect 320140 153428 324872 153456
rect 320140 153416 320146 153428
rect 324866 153416 324872 153428
rect 324924 153416 324930 153468
rect 324961 153459 325019 153465
rect 324961 153425 324973 153459
rect 325007 153456 325019 153459
rect 326154 153456 326160 153468
rect 325007 153428 326160 153456
rect 325007 153425 325019 153428
rect 324961 153419 325019 153425
rect 326154 153416 326160 153428
rect 326212 153416 326218 153468
rect 333974 153416 333980 153468
rect 334032 153456 334038 153468
rect 335906 153456 335912 153468
rect 334032 153428 335912 153456
rect 334032 153416 334038 153428
rect 335906 153416 335912 153428
rect 335964 153416 335970 153468
rect 342714 153416 342720 153468
rect 342772 153456 342778 153468
rect 345198 153456 345204 153468
rect 342772 153428 345204 153456
rect 342772 153416 342778 153428
rect 345198 153416 345204 153428
rect 345256 153416 345262 153468
rect 364150 153416 364156 153468
rect 364208 153456 364214 153468
rect 365070 153456 365076 153468
rect 364208 153428 365076 153456
rect 364208 153416 364214 153428
rect 365070 153416 365076 153428
rect 365128 153416 365134 153468
rect 365162 153416 365168 153468
rect 365220 153456 365226 153468
rect 366910 153456 366916 153468
rect 365220 153428 366916 153456
rect 365220 153416 365226 153428
rect 366910 153416 366916 153428
rect 366968 153416 366974 153468
rect 371602 153416 371608 153468
rect 371660 153456 371666 153468
rect 376662 153456 376668 153468
rect 371660 153428 376668 153456
rect 371660 153416 371666 153428
rect 376662 153416 376668 153428
rect 376720 153416 376726 153468
rect 384666 153416 384672 153468
rect 384724 153456 384730 153468
rect 396166 153456 396172 153468
rect 384724 153428 396172 153456
rect 384724 153416 384730 153428
rect 396166 153416 396172 153428
rect 396224 153416 396230 153468
rect 396994 153416 397000 153468
rect 397052 153456 397058 153468
rect 407758 153456 407764 153468
rect 397052 153428 407764 153456
rect 397052 153416 397058 153428
rect 407758 153416 407764 153428
rect 407816 153416 407822 153468
rect 489886 153456 489914 153496
rect 500402 153484 500408 153536
rect 500460 153524 500466 153536
rect 502978 153524 502984 153536
rect 500460 153496 502984 153524
rect 500460 153484 500466 153496
rect 502978 153484 502984 153496
rect 503036 153484 503042 153536
rect 506290 153456 506296 153468
rect 489886 153428 506296 153456
rect 506290 153416 506296 153428
rect 506348 153416 506354 153468
rect 511810 153416 511816 153468
rect 511868 153456 511874 153468
rect 523034 153456 523040 153468
rect 511868 153428 523040 153456
rect 511868 153416 511874 153428
rect 523034 153416 523040 153428
rect 523092 153416 523098 153468
rect 74258 153348 74264 153400
rect 74316 153388 74322 153400
rect 99282 153388 99288 153400
rect 74316 153360 99288 153388
rect 74316 153348 74322 153360
rect 99282 153348 99288 153360
rect 99340 153348 99346 153400
rect 102134 153348 102140 153400
rect 102192 153388 102198 153400
rect 114925 153391 114983 153397
rect 114925 153388 114937 153391
rect 102192 153360 114937 153388
rect 102192 153348 102198 153360
rect 114925 153357 114937 153360
rect 114971 153357 114983 153391
rect 120077 153391 120135 153397
rect 120077 153388 120089 153391
rect 114925 153351 114983 153357
rect 115032 153360 120089 153388
rect 36906 153280 36912 153332
rect 36964 153320 36970 153332
rect 108301 153323 108359 153329
rect 108301 153320 108313 153323
rect 36964 153292 108313 153320
rect 36964 153280 36970 153292
rect 108301 153289 108313 153292
rect 108347 153289 108359 153323
rect 108301 153283 108359 153289
rect 110414 153280 110420 153332
rect 110472 153320 110478 153332
rect 113637 153323 113695 153329
rect 113637 153320 113649 153323
rect 110472 153292 113649 153320
rect 110472 153280 110478 153292
rect 113637 153289 113649 153292
rect 113683 153289 113695 153323
rect 113637 153283 113695 153289
rect 113729 153323 113787 153329
rect 113729 153289 113741 153323
rect 113775 153320 113787 153323
rect 113775 153292 114140 153320
rect 113775 153289 113787 153292
rect 113729 153283 113787 153289
rect 23106 153212 23112 153264
rect 23164 153252 23170 153264
rect 75178 153252 75184 153264
rect 23164 153224 75184 153252
rect 23164 153212 23170 153224
rect 75178 153212 75184 153224
rect 75236 153212 75242 153264
rect 108942 153212 108948 153264
rect 109000 153252 109006 153264
rect 113910 153252 113916 153264
rect 109000 153224 113916 153252
rect 109000 153212 109006 153224
rect 113910 153212 113916 153224
rect 113968 153212 113974 153264
rect 114112 153252 114140 153292
rect 114186 153280 114192 153332
rect 114244 153320 114250 153332
rect 115032 153320 115060 153360
rect 120077 153357 120089 153360
rect 120123 153357 120135 153391
rect 120077 153351 120135 153357
rect 120166 153348 120172 153400
rect 120224 153388 120230 153400
rect 179414 153388 179420 153400
rect 120224 153360 179420 153388
rect 120224 153348 120230 153360
rect 179414 153348 179420 153360
rect 179472 153348 179478 153400
rect 179506 153348 179512 153400
rect 179564 153388 179570 153400
rect 188246 153388 188252 153400
rect 179564 153360 188252 153388
rect 179564 153348 179570 153360
rect 188246 153348 188252 153360
rect 188304 153348 188310 153400
rect 246942 153348 246948 153400
rect 247000 153388 247006 153400
rect 250714 153388 250720 153400
rect 247000 153360 250720 153388
rect 247000 153348 247006 153360
rect 250714 153348 250720 153360
rect 250772 153348 250778 153400
rect 262677 153391 262735 153397
rect 262677 153357 262689 153391
rect 262723 153388 262735 153391
rect 268194 153388 268200 153400
rect 262723 153360 268200 153388
rect 262723 153357 262735 153360
rect 262677 153351 262735 153357
rect 268194 153348 268200 153360
rect 268252 153348 268258 153400
rect 280706 153348 280712 153400
rect 280764 153388 280770 153400
rect 283834 153388 283840 153400
rect 280764 153360 283840 153388
rect 280764 153348 280770 153360
rect 283834 153348 283840 153360
rect 283892 153348 283898 153400
rect 285858 153348 285864 153400
rect 285916 153388 285922 153400
rect 287238 153388 287244 153400
rect 285916 153360 287244 153388
rect 285916 153348 285922 153360
rect 287238 153348 287244 153360
rect 287296 153348 287302 153400
rect 293954 153348 293960 153400
rect 294012 153388 294018 153400
rect 296990 153388 296996 153400
rect 294012 153360 296996 153388
rect 294012 153348 294018 153360
rect 296990 153348 296996 153360
rect 297048 153348 297054 153400
rect 298002 153348 298008 153400
rect 298060 153388 298066 153400
rect 302326 153388 302332 153400
rect 298060 153360 302332 153388
rect 298060 153348 298066 153360
rect 302326 153348 302332 153360
rect 302384 153348 302390 153400
rect 306558 153348 306564 153400
rect 306616 153388 306622 153400
rect 307938 153388 307944 153400
rect 306616 153360 307944 153388
rect 306616 153348 306622 153360
rect 307938 153348 307944 153360
rect 307996 153348 308002 153400
rect 308030 153348 308036 153400
rect 308088 153388 308094 153400
rect 310514 153388 310520 153400
rect 308088 153360 310520 153388
rect 308088 153348 308094 153360
rect 310514 153348 310520 153360
rect 310572 153348 310578 153400
rect 317322 153348 317328 153400
rect 317380 153388 317386 153400
rect 318334 153388 318340 153400
rect 317380 153360 318340 153388
rect 317380 153348 317386 153360
rect 318334 153348 318340 153360
rect 318392 153348 318398 153400
rect 324406 153348 324412 153400
rect 324464 153388 324470 153400
rect 325786 153388 325792 153400
rect 324464 153360 325792 153388
rect 324464 153348 324470 153360
rect 325786 153348 325792 153360
rect 325844 153348 325850 153400
rect 334066 153348 334072 153400
rect 334124 153388 334130 153400
rect 335446 153388 335452 153400
rect 334124 153360 335452 153388
rect 334124 153348 334130 153360
rect 335446 153348 335452 153360
rect 335504 153348 335510 153400
rect 338666 153348 338672 153400
rect 338724 153388 338730 153400
rect 341702 153388 341708 153400
rect 338724 153360 341708 153388
rect 338724 153348 338730 153360
rect 341702 153348 341708 153360
rect 341760 153348 341766 153400
rect 353386 153348 353392 153400
rect 353444 153388 353450 153400
rect 354858 153388 354864 153400
rect 353444 153360 354864 153388
rect 353444 153348 353450 153360
rect 354858 153348 354864 153360
rect 354916 153348 354922 153400
rect 363874 153348 363880 153400
rect 363932 153388 363938 153400
rect 364978 153388 364984 153400
rect 363932 153360 364984 153388
rect 363932 153348 363938 153360
rect 364978 153348 364984 153360
rect 365036 153348 365042 153400
rect 379422 153348 379428 153400
rect 379480 153388 379486 153400
rect 384850 153388 384856 153400
rect 379480 153360 384856 153388
rect 379480 153348 379486 153360
rect 384850 153348 384856 153360
rect 384908 153348 384914 153400
rect 387242 153348 387248 153400
rect 387300 153388 387306 153400
rect 400030 153388 400036 153400
rect 387300 153360 400036 153388
rect 387300 153348 387306 153360
rect 400030 153348 400036 153360
rect 400088 153348 400094 153400
rect 512730 153348 512736 153400
rect 512788 153388 512794 153400
rect 512788 153360 518894 153388
rect 512788 153348 512794 153360
rect 114244 153292 115060 153320
rect 115109 153323 115167 153329
rect 114244 153280 114250 153292
rect 115109 153289 115121 153323
rect 115155 153320 115167 153323
rect 123202 153320 123208 153332
rect 115155 153292 123208 153320
rect 115155 153289 115167 153292
rect 115109 153283 115167 153289
rect 123202 153280 123208 153292
rect 123260 153280 123266 153332
rect 124122 153280 124128 153332
rect 124180 153320 124186 153332
rect 125045 153323 125103 153329
rect 124180 153292 124996 153320
rect 124180 153280 124186 153292
rect 115198 153252 115204 153264
rect 114112 153224 115204 153252
rect 115198 153212 115204 153224
rect 115256 153212 115262 153264
rect 116762 153212 116768 153264
rect 116820 153252 116826 153264
rect 124861 153255 124919 153261
rect 124861 153252 124873 153255
rect 116820 153224 124873 153252
rect 116820 153212 116826 153224
rect 124861 153221 124873 153224
rect 124907 153221 124919 153255
rect 124968 153252 124996 153292
rect 125045 153289 125057 153323
rect 125091 153320 125103 153323
rect 157702 153320 157708 153332
rect 125091 153292 157708 153320
rect 125091 153289 125103 153292
rect 125045 153283 125103 153289
rect 157702 153280 157708 153292
rect 157760 153280 157766 153332
rect 158806 153280 158812 153332
rect 158864 153320 158870 153332
rect 162210 153320 162216 153332
rect 158864 153292 162216 153320
rect 158864 153280 158870 153292
rect 162210 153280 162216 153292
rect 162268 153280 162274 153332
rect 166261 153323 166319 153329
rect 166261 153289 166273 153323
rect 166307 153320 166319 153323
rect 194778 153320 194784 153332
rect 166307 153292 194784 153320
rect 166307 153289 166319 153292
rect 166261 153283 166319 153289
rect 194778 153280 194784 153292
rect 194836 153280 194842 153332
rect 197262 153280 197268 153332
rect 197320 153320 197326 153332
rect 512822 153320 512828 153332
rect 197320 153292 512828 153320
rect 197320 153280 197326 153292
rect 512822 153280 512828 153292
rect 512880 153280 512886 153332
rect 518866 153320 518894 153360
rect 520274 153320 520280 153332
rect 518866 153292 520280 153320
rect 520274 153280 520280 153292
rect 520332 153280 520338 153332
rect 145926 153252 145932 153264
rect 124968 153224 145932 153252
rect 124861 153215 124919 153221
rect 145926 153212 145932 153224
rect 145984 153212 145990 153264
rect 149054 153212 149060 153264
rect 149112 153252 149118 153264
rect 169386 153252 169392 153264
rect 149112 153224 169392 153252
rect 149112 153212 149118 153224
rect 169386 153212 169392 153224
rect 169444 153212 169450 153264
rect 171134 153212 171140 153264
rect 171192 153252 171198 153264
rect 514110 153252 514116 153264
rect 171192 153224 514116 153252
rect 171192 153212 171198 153224
rect 514110 153212 514116 153224
rect 514168 153212 514174 153264
rect 515398 153212 515404 153264
rect 515456 153252 515462 153264
rect 520458 153252 520464 153264
rect 515456 153224 520464 153252
rect 515456 153212 515462 153224
rect 520458 153212 520464 153224
rect 520516 153212 520522 153264
rect 60826 153144 60832 153196
rect 60884 153184 60890 153196
rect 160278 153184 160284 153196
rect 60884 153156 160284 153184
rect 60884 153144 60890 153156
rect 160278 153144 160284 153156
rect 160336 153144 160342 153196
rect 170122 153144 170128 153196
rect 170180 153184 170186 153196
rect 233234 153184 233240 153196
rect 170180 153156 233240 153184
rect 170180 153144 170186 153156
rect 233234 153144 233240 153156
rect 233292 153144 233298 153196
rect 471146 153144 471152 153196
rect 471204 153184 471210 153196
rect 525794 153184 525800 153196
rect 471204 153156 525800 153184
rect 471204 153144 471210 153156
rect 525794 153144 525800 153156
rect 525852 153144 525858 153196
rect 49142 153076 49148 153128
rect 49200 153116 49206 153128
rect 152458 153116 152464 153128
rect 49200 153088 152464 153116
rect 49200 153076 49206 153088
rect 152458 153076 152464 153088
rect 152516 153076 152522 153128
rect 158898 153076 158904 153128
rect 158956 153116 158962 153128
rect 223574 153116 223580 153128
rect 158956 153088 223580 153116
rect 158956 153076 158962 153088
rect 223574 153076 223580 153088
rect 223632 153076 223638 153128
rect 423582 153076 423588 153128
rect 423640 153116 423646 153128
rect 454678 153116 454684 153128
rect 423640 153088 454684 153116
rect 423640 153076 423646 153088
rect 454678 153076 454684 153088
rect 454736 153076 454742 153128
rect 475746 153076 475752 153128
rect 475804 153116 475810 153128
rect 532602 153116 532608 153128
rect 475804 153088 532608 153116
rect 475804 153076 475810 153088
rect 532602 153076 532608 153088
rect 532660 153076 532666 153128
rect 45278 153008 45284 153060
rect 45336 153048 45342 153060
rect 149882 153048 149888 153060
rect 45336 153020 149888 153048
rect 45336 153008 45342 153020
rect 149882 153008 149888 153020
rect 149940 153008 149946 153060
rect 153102 153008 153108 153060
rect 153160 153048 153166 153060
rect 158441 153051 158499 153057
rect 158441 153048 158453 153051
rect 153160 153020 158453 153048
rect 153160 153008 153166 153020
rect 158441 153017 158453 153020
rect 158487 153017 158499 153051
rect 158441 153011 158499 153017
rect 162302 153008 162308 153060
rect 162360 153048 162366 153060
rect 227898 153048 227904 153060
rect 162360 153020 227904 153048
rect 162360 153008 162366 153020
rect 227898 153008 227904 153020
rect 227956 153008 227962 153060
rect 255774 153008 255780 153060
rect 255832 153048 255838 153060
rect 290366 153048 290372 153060
rect 255832 153020 290372 153048
rect 255832 153008 255838 153020
rect 290366 153008 290372 153020
rect 290424 153008 290430 153060
rect 431494 153008 431500 153060
rect 431552 153048 431558 153060
rect 466270 153048 466276 153060
rect 431552 153020 466276 153048
rect 431552 153008 431558 153020
rect 466270 153008 466276 153020
rect 466328 153008 466334 153060
rect 475102 153008 475108 153060
rect 475160 153048 475166 153060
rect 531682 153048 531688 153060
rect 475160 153020 531688 153048
rect 475160 153008 475166 153020
rect 531682 153008 531688 153020
rect 531740 153008 531746 153060
rect 42334 152940 42340 152992
rect 42392 152980 42398 152992
rect 147950 152980 147956 152992
rect 42392 152952 147956 152980
rect 42392 152940 42398 152952
rect 147950 152940 147956 152952
rect 148008 152940 148014 152992
rect 152550 152940 152556 152992
rect 152608 152980 152614 152992
rect 221366 152980 221372 152992
rect 152608 152952 221372 152980
rect 152608 152940 152614 152952
rect 221366 152940 221372 152952
rect 221424 152940 221430 152992
rect 248138 152940 248144 152992
rect 248196 152980 248202 152992
rect 285122 152980 285128 152992
rect 248196 152952 285128 152980
rect 248196 152940 248202 152952
rect 285122 152940 285128 152952
rect 285180 152940 285186 152992
rect 434070 152940 434076 152992
rect 434128 152980 434134 152992
rect 470226 152980 470232 152992
rect 434128 152952 470232 152980
rect 434128 152940 434134 152952
rect 470226 152940 470232 152952
rect 470284 152940 470290 152992
rect 478782 152940 478788 152992
rect 478840 152980 478846 152992
rect 537478 152980 537484 152992
rect 478840 152952 537484 152980
rect 478840 152940 478846 152952
rect 537478 152940 537484 152952
rect 537536 152940 537542 152992
rect 41322 152872 41328 152924
rect 41380 152912 41386 152924
rect 147214 152912 147220 152924
rect 41380 152884 147220 152912
rect 41380 152872 41386 152884
rect 147214 152872 147220 152884
rect 147272 152872 147278 152924
rect 150526 152872 150532 152924
rect 150584 152912 150590 152924
rect 220078 152912 220084 152924
rect 150584 152884 220084 152912
rect 150584 152872 150590 152884
rect 220078 152872 220084 152884
rect 220136 152872 220142 152924
rect 238294 152872 238300 152924
rect 238352 152912 238358 152924
rect 278774 152912 278780 152924
rect 238352 152884 278780 152912
rect 238352 152872 238358 152884
rect 278774 152872 278780 152884
rect 278832 152872 278838 152924
rect 439314 152872 439320 152924
rect 439372 152912 439378 152924
rect 478046 152912 478052 152924
rect 439372 152884 478052 152912
rect 439372 152872 439378 152884
rect 478046 152872 478052 152884
rect 478104 152872 478110 152924
rect 482830 152872 482836 152924
rect 482888 152912 482894 152924
rect 543366 152912 543372 152924
rect 482888 152884 543372 152912
rect 482888 152872 482894 152884
rect 543366 152872 543372 152884
rect 543424 152872 543430 152924
rect 31662 152804 31668 152856
rect 31720 152844 31726 152856
rect 139486 152844 139492 152856
rect 31720 152816 139492 152844
rect 31720 152804 31726 152816
rect 139486 152804 139492 152816
rect 139544 152804 139550 152856
rect 140774 152804 140780 152856
rect 140832 152844 140838 152856
rect 141418 152844 141424 152856
rect 140832 152816 141424 152844
rect 140832 152804 140838 152816
rect 141418 152804 141424 152816
rect 141476 152804 141482 152856
rect 142706 152804 142712 152856
rect 142764 152844 142770 152856
rect 214926 152844 214932 152856
rect 142764 152816 214932 152844
rect 142764 152804 142770 152816
rect 214926 152804 214932 152816
rect 214984 152804 214990 152856
rect 232406 152804 232412 152856
rect 232464 152844 232470 152856
rect 274726 152844 274732 152856
rect 232464 152816 274732 152844
rect 232464 152804 232470 152816
rect 274726 152804 274732 152816
rect 274784 152804 274790 152856
rect 440602 152804 440608 152856
rect 440660 152844 440666 152856
rect 479978 152844 479984 152856
rect 440660 152816 479984 152844
rect 440660 152804 440666 152816
rect 479978 152804 479984 152816
rect 480036 152804 480042 152856
rect 485498 152804 485504 152856
rect 485556 152844 485562 152856
rect 547230 152844 547236 152856
rect 485556 152816 547236 152844
rect 485556 152804 485562 152816
rect 547230 152804 547236 152816
rect 547288 152804 547294 152856
rect 22094 152736 22100 152788
rect 22152 152776 22158 152788
rect 22152 152748 127572 152776
rect 22152 152736 22158 152748
rect 11514 152668 11520 152720
rect 11572 152708 11578 152720
rect 122834 152708 122840 152720
rect 11572 152680 122840 152708
rect 11572 152668 11578 152680
rect 122834 152668 122840 152680
rect 122892 152668 122898 152720
rect 124214 152668 124220 152720
rect 124272 152708 124278 152720
rect 127437 152711 127495 152717
rect 127437 152708 127449 152711
rect 124272 152680 127449 152708
rect 124272 152668 124278 152680
rect 127437 152677 127449 152680
rect 127483 152677 127495 152711
rect 127437 152671 127495 152677
rect 10134 152600 10140 152652
rect 10192 152640 10198 152652
rect 126422 152640 126428 152652
rect 10192 152612 126428 152640
rect 10192 152600 10198 152612
rect 126422 152600 126428 152612
rect 126480 152600 126486 152652
rect 127544 152640 127572 152748
rect 138934 152736 138940 152788
rect 138992 152776 138998 152788
rect 212534 152776 212540 152788
rect 138992 152748 212540 152776
rect 138992 152736 138998 152748
rect 212534 152736 212540 152748
rect 212592 152736 212598 152788
rect 224586 152736 224592 152788
rect 224644 152776 224650 152788
rect 269574 152776 269580 152788
rect 224644 152748 269580 152776
rect 224644 152736 224650 152748
rect 269574 152736 269580 152748
rect 269632 152736 269638 152788
rect 486142 152736 486148 152788
rect 486200 152776 486206 152788
rect 548242 152776 548248 152788
rect 486200 152748 548248 152776
rect 486200 152736 486206 152748
rect 548242 152736 548248 152748
rect 548300 152736 548306 152788
rect 127621 152711 127679 152717
rect 127621 152677 127633 152711
rect 127667 152708 127679 152711
rect 195241 152711 195299 152717
rect 195241 152708 195253 152711
rect 127667 152680 195253 152708
rect 127667 152677 127679 152680
rect 127621 152671 127679 152677
rect 195241 152677 195253 152680
rect 195287 152677 195299 152711
rect 195241 152671 195299 152677
rect 209130 152668 209136 152720
rect 209188 152708 209194 152720
rect 259086 152708 259092 152720
rect 209188 152680 259092 152708
rect 209188 152668 209194 152680
rect 259086 152668 259092 152680
rect 259144 152668 259150 152720
rect 445662 152668 445668 152720
rect 445720 152708 445726 152720
rect 487798 152708 487804 152720
rect 445720 152680 487804 152708
rect 445720 152668 445726 152680
rect 487798 152668 487804 152680
rect 487856 152668 487862 152720
rect 488074 152668 488080 152720
rect 488132 152708 488138 152720
rect 551186 152708 551192 152720
rect 488132 152680 551192 152708
rect 488132 152668 488138 152680
rect 551186 152668 551192 152680
rect 551244 152668 551250 152720
rect 134242 152640 134248 152652
rect 127544 152612 134248 152640
rect 134242 152600 134248 152612
rect 134300 152600 134306 152652
rect 135898 152600 135904 152652
rect 135956 152640 135962 152652
rect 210326 152640 210332 152652
rect 135956 152612 210332 152640
rect 135956 152600 135962 152612
rect 210326 152600 210332 152612
rect 210384 152600 210390 152652
rect 211890 152600 211896 152652
rect 211948 152640 211954 152652
rect 212442 152640 212448 152652
rect 211948 152612 212448 152640
rect 211948 152600 211954 152612
rect 212442 152600 212448 152612
rect 212500 152600 212506 152652
rect 216950 152600 216956 152652
rect 217008 152640 217014 152652
rect 264330 152640 264336 152652
rect 217008 152612 264336 152640
rect 217008 152600 217014 152612
rect 264330 152600 264336 152612
rect 264388 152600 264394 152652
rect 271414 152600 271420 152652
rect 271472 152640 271478 152652
rect 300854 152640 300860 152652
rect 271472 152612 300860 152640
rect 271472 152600 271478 152612
rect 300854 152600 300860 152612
rect 300912 152600 300918 152652
rect 446490 152600 446496 152652
rect 446548 152640 446554 152652
rect 488810 152640 488816 152652
rect 446548 152612 488816 152640
rect 446548 152600 446554 152612
rect 488810 152600 488816 152612
rect 488868 152600 488874 152652
rect 489362 152600 489368 152652
rect 489420 152640 489426 152652
rect 553118 152640 553124 152652
rect 489420 152612 553124 152640
rect 489420 152600 489426 152612
rect 553118 152600 553124 152612
rect 553176 152600 553182 152652
rect 7282 152532 7288 152584
rect 7340 152572 7346 152584
rect 124490 152572 124496 152584
rect 7340 152544 124496 152572
rect 7340 152532 7346 152544
rect 124490 152532 124496 152544
rect 124548 152532 124554 152584
rect 127158 152532 127164 152584
rect 127216 152572 127222 152584
rect 204530 152572 204536 152584
rect 127216 152544 204536 152572
rect 127216 152532 127222 152544
rect 204530 152532 204536 152544
rect 204588 152532 204594 152584
rect 214561 152575 214619 152581
rect 214561 152572 214573 152575
rect 204916 152544 214573 152572
rect 2406 152464 2412 152516
rect 2464 152504 2470 152516
rect 121454 152504 121460 152516
rect 2464 152476 121460 152504
rect 2464 152464 2470 152476
rect 121454 152464 121460 152476
rect 121512 152464 121518 152516
rect 123294 152464 123300 152516
rect 123352 152504 123358 152516
rect 201862 152504 201868 152516
rect 123352 152476 201868 152504
rect 123352 152464 123358 152476
rect 201862 152464 201868 152476
rect 201920 152464 201926 152516
rect 203242 152464 203248 152516
rect 203300 152504 203306 152516
rect 204916 152504 204944 152544
rect 214561 152541 214573 152544
rect 214607 152541 214619 152575
rect 214561 152535 214619 152541
rect 220722 152532 220728 152584
rect 220780 152572 220786 152584
rect 266906 152572 266912 152584
rect 220780 152544 266912 152572
rect 220780 152532 220786 152544
rect 266906 152532 266912 152544
rect 266964 152532 266970 152584
rect 267550 152532 267556 152584
rect 267608 152572 267614 152584
rect 298186 152572 298192 152584
rect 267608 152544 298192 152572
rect 267608 152532 267614 152544
rect 298186 152532 298192 152544
rect 298244 152532 298250 152584
rect 449710 152532 449716 152584
rect 449768 152572 449774 152584
rect 449768 152544 491156 152572
rect 449768 152532 449774 152544
rect 203300 152476 204944 152504
rect 203300 152464 203306 152476
rect 208026 152464 208032 152516
rect 208084 152504 208090 152516
rect 258442 152504 258448 152516
rect 208084 152476 258448 152504
rect 208084 152464 208090 152476
rect 258442 152464 258448 152476
rect 258500 152464 258506 152516
rect 259730 152464 259736 152516
rect 259788 152504 259794 152516
rect 292942 152504 292948 152516
rect 259788 152476 292948 152504
rect 259788 152464 259794 152476
rect 292942 152464 292948 152476
rect 293000 152464 293006 152516
rect 418522 152464 418528 152516
rect 418580 152504 418586 152516
rect 446858 152504 446864 152516
rect 418580 152476 446864 152504
rect 418580 152464 418586 152476
rect 446858 152464 446864 152476
rect 446916 152464 446922 152516
rect 452286 152464 452292 152516
rect 452344 152504 452350 152516
rect 491021 152507 491079 152513
rect 491021 152504 491033 152507
rect 452344 152476 491033 152504
rect 452344 152464 452350 152476
rect 491021 152473 491033 152476
rect 491067 152473 491079 152507
rect 491128 152504 491156 152544
rect 493318 152532 493324 152584
rect 493376 152572 493382 152584
rect 558822 152572 558828 152584
rect 493376 152544 558828 152572
rect 493376 152532 493382 152544
rect 558822 152532 558828 152544
rect 558880 152532 558886 152584
rect 493686 152504 493692 152516
rect 491128 152476 493692 152504
rect 491021 152467 491079 152473
rect 493686 152464 493692 152476
rect 493744 152464 493750 152516
rect 498102 152464 498108 152516
rect 498160 152504 498166 152516
rect 566734 152504 566740 152516
rect 498160 152476 566740 152504
rect 498160 152464 498166 152476
rect 566734 152464 566740 152476
rect 566792 152464 566798 152516
rect 57974 152396 57980 152448
rect 58032 152436 58038 152448
rect 158346 152436 158352 152448
rect 58032 152408 158352 152436
rect 58032 152396 58038 152408
rect 158346 152396 158352 152408
rect 158404 152396 158410 152448
rect 158441 152439 158499 152445
rect 158441 152405 158453 152439
rect 158487 152436 158499 152439
rect 215570 152436 215576 152448
rect 158487 152408 215576 152436
rect 158487 152405 158499 152408
rect 158441 152399 158499 152405
rect 215570 152396 215576 152408
rect 215628 152396 215634 152448
rect 468570 152396 468576 152448
rect 468628 152436 468634 152448
rect 521930 152436 521936 152448
rect 468628 152408 521936 152436
rect 468628 152396 468634 152408
rect 521930 152396 521936 152408
rect 521988 152396 521994 152448
rect 72602 152328 72608 152380
rect 72660 152368 72666 152380
rect 168374 152368 168380 152380
rect 72660 152340 168380 152368
rect 72660 152328 72666 152340
rect 168374 152328 168380 152340
rect 168432 152328 168438 152380
rect 179782 152328 179788 152380
rect 179840 152368 179846 152380
rect 239582 152368 239588 152380
rect 179840 152340 239588 152368
rect 179840 152328 179846 152340
rect 239582 152328 239588 152340
rect 239640 152328 239646 152380
rect 465994 152328 466000 152380
rect 466052 152368 466058 152380
rect 517974 152368 517980 152380
rect 466052 152340 517980 152368
rect 466052 152328 466058 152340
rect 517974 152328 517980 152340
rect 518032 152328 518038 152380
rect 80330 152260 80336 152312
rect 80388 152300 80394 152312
rect 173250 152300 173256 152312
rect 80388 152272 173256 152300
rect 80388 152260 80394 152272
rect 173250 152260 173256 152272
rect 173308 152260 173314 152312
rect 181806 152260 181812 152312
rect 181864 152300 181870 152312
rect 240962 152300 240968 152312
rect 181864 152272 240968 152300
rect 181864 152260 181870 152272
rect 240962 152260 240968 152272
rect 241020 152260 241026 152312
rect 458818 152260 458824 152312
rect 458876 152300 458882 152312
rect 507302 152300 507308 152312
rect 458876 152272 507308 152300
rect 458876 152260 458882 152272
rect 507302 152260 507308 152272
rect 507360 152260 507366 152312
rect 73522 152192 73528 152244
rect 73580 152232 73586 152244
rect 169064 152232 169070 152244
rect 73580 152204 169070 152232
rect 73580 152192 73586 152204
rect 169064 152192 169070 152204
rect 169122 152192 169128 152244
rect 175826 152192 175832 152244
rect 175884 152232 175890 152244
rect 175884 152204 177068 152232
rect 175884 152192 175890 152204
rect 85206 152124 85212 152176
rect 85264 152164 85270 152176
rect 176884 152164 176890 152176
rect 85264 152136 176890 152164
rect 85264 152124 85270 152136
rect 176884 152124 176890 152136
rect 176942 152124 176948 152176
rect 177040 152164 177068 152204
rect 178218 152192 178224 152244
rect 178276 152232 178282 152244
rect 236684 152232 236690 152244
rect 178276 152204 236690 152232
rect 178276 152192 178282 152204
rect 236684 152192 236690 152204
rect 236742 152192 236748 152244
rect 453896 152192 453902 152244
rect 453954 152232 453960 152244
rect 500494 152232 500500 152244
rect 453954 152204 500500 152232
rect 453954 152192 453960 152204
rect 500494 152192 500500 152204
rect 500552 152192 500558 152244
rect 177040 152136 180794 152164
rect 88150 152056 88156 152108
rect 88208 152096 88214 152108
rect 178816 152096 178822 152108
rect 88208 152068 178822 152096
rect 88208 152056 88214 152068
rect 178816 152056 178822 152068
rect 178874 152056 178880 152108
rect 180766 152096 180794 152136
rect 185762 152124 185768 152176
rect 185820 152164 185826 152176
rect 243860 152164 243866 152176
rect 185820 152136 243866 152164
rect 185820 152124 185826 152136
rect 243860 152124 243866 152136
rect 243918 152124 243924 152176
rect 450676 152124 450682 152176
rect 450734 152164 450740 152176
rect 491021 152167 491079 152173
rect 450734 152136 490972 152164
rect 450734 152124 450740 152136
rect 231440 152096 231446 152108
rect 180766 152068 231446 152096
rect 231440 152056 231446 152068
rect 231498 152056 231504 152108
rect 451320 152056 451326 152108
rect 451378 152096 451384 152108
rect 490944 152096 490972 152136
rect 491021 152133 491033 152167
rect 491067 152164 491079 152167
rect 497550 152164 497556 152176
rect 491067 152136 497556 152164
rect 491067 152133 491079 152136
rect 491021 152127 491079 152133
rect 497550 152124 497556 152136
rect 497608 152124 497614 152176
rect 495618 152096 495624 152108
rect 451378 152068 490880 152096
rect 490944 152068 495624 152096
rect 451378 152056 451384 152068
rect 95970 151988 95976 152040
rect 96028 152028 96034 152040
rect 183646 152028 183652 152040
rect 96028 152000 183652 152028
rect 96028 151988 96034 152000
rect 183646 151988 183652 152000
rect 183704 151988 183710 152040
rect 197446 151988 197452 152040
rect 197504 152028 197510 152040
rect 251358 152028 251364 152040
rect 197504 152000 251364 152028
rect 197504 151988 197510 152000
rect 251358 151988 251364 152000
rect 251416 151988 251422 152040
rect 447778 151988 447784 152040
rect 447836 152028 447842 152040
rect 490742 152028 490748 152040
rect 447836 152000 490748 152028
rect 447836 151988 447842 152000
rect 490742 151988 490748 152000
rect 490800 151988 490806 152040
rect 490852 152028 490880 152068
rect 495618 152056 495624 152068
rect 495676 152056 495682 152108
rect 496446 152056 496452 152108
rect 496504 152056 496510 152108
rect 496464 152028 496492 152056
rect 490852 152000 496492 152028
rect 111518 151920 111524 151972
rect 111576 151960 111582 151972
rect 194042 151960 194048 151972
rect 111576 151932 194048 151960
rect 111576 151920 111582 151932
rect 194042 151920 194048 151932
rect 194100 151920 194106 151972
rect 195241 151963 195299 151969
rect 195241 151929 195253 151963
rect 195287 151960 195299 151963
rect 202506 151960 202512 151972
rect 195287 151932 202512 151960
rect 195287 151929 195299 151932
rect 195241 151923 195299 151929
rect 202506 151920 202512 151932
rect 202564 151920 202570 151972
rect 214561 151963 214619 151969
rect 214561 151929 214573 151963
rect 214607 151960 214619 151963
rect 249334 151960 249340 151972
rect 214607 151932 249340 151960
rect 214607 151929 214619 151932
rect 214561 151923 214619 151929
rect 249334 151920 249340 151932
rect 249392 151920 249398 151972
rect 444282 151920 444288 151972
rect 444340 151960 444346 151972
rect 485682 151960 485688 151972
rect 444340 151932 485688 151960
rect 444340 151920 444346 151932
rect 485682 151920 485688 151932
rect 485740 151920 485746 151972
rect 75178 151892 75184 151904
rect 75139 151864 75184 151892
rect 75178 151852 75184 151864
rect 75236 151852 75242 151904
rect 78122 151892 78128 151904
rect 78083 151864 78128 151892
rect 78122 151852 78128 151864
rect 78180 151852 78186 151904
rect 88334 151892 88340 151904
rect 88295 151864 88340 151892
rect 88334 151852 88340 151864
rect 88392 151852 88398 151904
rect 91922 151892 91928 151904
rect 91883 151864 91928 151892
rect 91922 151852 91928 151864
rect 91980 151852 91986 151904
rect 95142 151892 95148 151904
rect 95103 151864 95148 151892
rect 95142 151852 95148 151864
rect 95200 151852 95206 151904
rect 99282 151892 99288 151904
rect 99243 151864 99288 151892
rect 99282 151852 99288 151864
rect 99340 151852 99346 151904
rect 112438 151892 112444 151904
rect 103486 151864 112444 151892
rect 41325 151827 41383 151833
rect 41325 151793 41337 151827
rect 41371 151824 41383 151827
rect 103486 151824 103514 151864
rect 112438 151852 112444 151864
rect 112496 151852 112502 151904
rect 116394 151852 116400 151904
rect 116452 151892 116458 151904
rect 197354 151892 197360 151904
rect 116452 151864 197360 151892
rect 116452 151852 116458 151864
rect 197354 151852 197360 151864
rect 197412 151852 197418 151904
rect 199102 151852 199108 151904
rect 199160 151892 199166 151904
rect 244366 151892 244372 151904
rect 199160 151864 244372 151892
rect 199160 151852 199166 151864
rect 244366 151852 244372 151864
rect 244424 151852 244430 151904
rect 105630 151824 105636 151836
rect 41371 151796 103514 151824
rect 105591 151796 105636 151824
rect 41371 151793 41383 151796
rect 41325 151787 41383 151793
rect 105630 151784 105636 151796
rect 105688 151784 105694 151836
rect 146478 151784 146484 151836
rect 146536 151824 146542 151836
rect 146536 151796 212304 151824
rect 146536 151784 146542 151796
rect 25498 151716 25504 151768
rect 25556 151756 25562 151768
rect 127710 151756 127716 151768
rect 25556 151728 127716 151756
rect 25556 151716 25562 151728
rect 127710 151716 127716 151728
rect 127768 151716 127774 151768
rect 212276 151756 212304 151796
rect 212442 151784 212448 151836
rect 212500 151824 212506 151836
rect 252002 151824 252008 151836
rect 212500 151796 252008 151824
rect 212500 151784 212506 151796
rect 252002 151784 252008 151796
rect 252060 151784 252066 151836
rect 503622 151784 503628 151836
rect 503680 151824 503686 151836
rect 520550 151824 520556 151836
rect 503680 151796 520556 151824
rect 503680 151784 503686 151796
rect 520550 151784 520556 151796
rect 520608 151784 520614 151836
rect 212902 151756 212908 151768
rect 212276 151728 212908 151756
rect 212902 151716 212908 151728
rect 212960 151716 212966 151768
rect 64414 151648 64420 151700
rect 64472 151688 64478 151700
rect 171134 151688 171140 151700
rect 64472 151660 171140 151688
rect 64472 151648 64478 151660
rect 171134 151648 171140 151660
rect 171192 151648 171198 151700
rect 505002 151648 505008 151700
rect 505060 151688 505066 151700
rect 528554 151688 528560 151700
rect 505060 151660 528560 151688
rect 505060 151648 505066 151660
rect 528554 151648 528560 151660
rect 528612 151648 528618 151700
rect 50614 151580 50620 151632
rect 50672 151620 50678 151632
rect 197262 151620 197268 151632
rect 50672 151592 197268 151620
rect 50672 151580 50678 151592
rect 197262 151580 197268 151592
rect 197320 151580 197326 151632
rect 506934 151620 506940 151632
rect 506895 151592 506940 151620
rect 506934 151580 506940 151592
rect 506992 151580 506998 151632
rect 3050 151512 3056 151564
rect 3108 151552 3114 151564
rect 117038 151552 117044 151564
rect 3108 151524 117044 151552
rect 3108 151512 3114 151524
rect 117038 151512 117044 151524
rect 117096 151512 117102 151564
rect 118326 151512 118332 151564
rect 118384 151552 118390 151564
rect 127713 151555 127771 151561
rect 118384 151524 127664 151552
rect 118384 151512 118390 151524
rect 3234 151444 3240 151496
rect 3292 151484 3298 151496
rect 3292 151456 115888 151484
rect 3292 151444 3298 151456
rect 40126 151416 40132 151428
rect 40087 151388 40132 151416
rect 40126 151376 40132 151388
rect 40184 151376 40190 151428
rect 43806 151376 43812 151428
rect 43864 151416 43870 151428
rect 115382 151416 115388 151428
rect 43864 151388 115388 151416
rect 43864 151376 43870 151388
rect 115382 151376 115388 151388
rect 115440 151376 115446 151428
rect 115860 151416 115888 151456
rect 117130 151444 117136 151496
rect 117188 151484 117194 151496
rect 127529 151487 127587 151493
rect 127529 151484 127541 151487
rect 117188 151456 127541 151484
rect 117188 151444 117194 151456
rect 127529 151453 127541 151456
rect 127575 151453 127587 151487
rect 127636 151484 127664 151524
rect 127713 151521 127725 151555
rect 127759 151552 127771 151555
rect 503714 151552 503720 151564
rect 127759 151524 503720 151552
rect 127759 151521 127771 151524
rect 127713 151515 127771 151521
rect 503714 151512 503720 151524
rect 503772 151512 503778 151564
rect 505646 151512 505652 151564
rect 505704 151552 505710 151564
rect 545114 151552 545120 151564
rect 505704 151524 545120 151552
rect 505704 151512 505710 151524
rect 545114 151512 545120 151524
rect 545172 151512 545178 151564
rect 575474 151484 575480 151496
rect 127636 151456 575480 151484
rect 127529 151447 127587 151453
rect 575474 151444 575480 151456
rect 575532 151444 575538 151496
rect 117314 151416 117320 151428
rect 115860 151388 117320 151416
rect 117314 151376 117320 151388
rect 117372 151376 117378 151428
rect 118418 151376 118424 151428
rect 118476 151416 118482 151428
rect 575566 151416 575572 151428
rect 118476 151388 575572 151416
rect 118476 151376 118482 151388
rect 575566 151376 575572 151388
rect 575624 151376 575630 151428
rect 3418 151308 3424 151360
rect 3476 151348 3482 151360
rect 115014 151348 115020 151360
rect 3476 151320 115020 151348
rect 3476 151308 3482 151320
rect 115014 151308 115020 151320
rect 115072 151308 115078 151360
rect 116946 151308 116952 151360
rect 117004 151348 117010 151360
rect 507762 151348 507768 151360
rect 117004 151320 507768 151348
rect 117004 151308 117010 151320
rect 507762 151308 507768 151320
rect 507820 151308 507826 151360
rect 508866 151348 508872 151360
rect 508827 151320 508872 151348
rect 508866 151308 508872 151320
rect 508924 151308 508930 151360
rect 515398 151348 515404 151360
rect 509206 151320 515404 151348
rect 4798 151240 4804 151292
rect 4856 151280 4862 151292
rect 112622 151280 112628 151292
rect 4856 151252 112628 151280
rect 4856 151240 4862 151252
rect 112622 151240 112628 151252
rect 112680 151240 112686 151292
rect 114002 151240 114008 151292
rect 114060 151280 114066 151292
rect 506937 151283 506995 151289
rect 506937 151280 506949 151283
rect 114060 151252 506949 151280
rect 114060 151240 114066 151252
rect 506937 151249 506949 151252
rect 506983 151249 506995 151283
rect 506937 151243 506995 151249
rect 99285 151215 99343 151221
rect 99285 151181 99297 151215
rect 99331 151212 99343 151215
rect 509206 151212 509234 151320
rect 515398 151308 515404 151320
rect 515456 151308 515462 151360
rect 518618 151308 518624 151360
rect 518676 151348 518682 151360
rect 518676 151320 518894 151348
rect 518676 151308 518682 151320
rect 518866 151280 518894 151320
rect 519262 151308 519268 151360
rect 519320 151348 519326 151360
rect 520366 151348 520372 151360
rect 519320 151320 520372 151348
rect 519320 151308 519326 151320
rect 520366 151308 520372 151320
rect 520424 151308 520430 151360
rect 520642 151280 520648 151292
rect 518866 151252 520648 151280
rect 520642 151240 520648 151252
rect 520700 151240 520706 151292
rect 99331 151184 509234 151212
rect 99331 151181 99343 151184
rect 99285 151175 99343 151181
rect 95145 151147 95203 151153
rect 95145 151113 95157 151147
rect 95191 151144 95203 151147
rect 521746 151144 521752 151156
rect 95191 151116 521752 151144
rect 95191 151113 95203 151116
rect 95145 151107 95203 151113
rect 521746 151104 521752 151116
rect 521804 151104 521810 151156
rect 5166 151036 5172 151088
rect 5224 151076 5230 151088
rect 41325 151079 41383 151085
rect 41325 151076 41337 151079
rect 5224 151048 41337 151076
rect 5224 151036 5230 151048
rect 41325 151045 41337 151048
rect 41371 151045 41383 151079
rect 41325 151039 41383 151045
rect 75181 151079 75239 151085
rect 75181 151045 75193 151079
rect 75227 151076 75239 151079
rect 508869 151079 508927 151085
rect 508869 151076 508881 151079
rect 75227 151048 508881 151076
rect 75227 151045 75239 151048
rect 75181 151039 75239 151045
rect 508869 151045 508881 151048
rect 508915 151045 508927 151079
rect 508869 151039 508927 151045
rect 78125 151011 78183 151017
rect 78125 150977 78137 151011
rect 78171 151008 78183 151011
rect 521838 151008 521844 151020
rect 78171 150980 521844 151008
rect 78171 150977 78183 150980
rect 78125 150971 78183 150977
rect 521838 150968 521844 150980
rect 521896 150968 521902 151020
rect 40129 150943 40187 150949
rect 40129 150909 40141 150943
rect 40175 150940 40187 150943
rect 522298 150940 522304 150952
rect 40175 150912 522304 150940
rect 40175 150909 40187 150912
rect 40129 150903 40187 150909
rect 522298 150900 522304 150912
rect 522356 150900 522362 150952
rect 3878 150832 3884 150884
rect 3936 150872 3942 150884
rect 112714 150872 112720 150884
rect 3936 150844 112720 150872
rect 3936 150832 3942 150844
rect 112714 150832 112720 150844
rect 112772 150832 112778 150884
rect 4154 150764 4160 150816
rect 4212 150804 4218 150816
rect 114278 150804 114284 150816
rect 4212 150776 114284 150804
rect 4212 150764 4218 150776
rect 114278 150764 114284 150776
rect 114336 150764 114342 150816
rect 3694 150696 3700 150748
rect 3752 150736 3758 150748
rect 114370 150736 114376 150748
rect 3752 150708 114376 150736
rect 3752 150696 3758 150708
rect 114370 150696 114376 150708
rect 114428 150696 114434 150748
rect 117314 150696 117320 150748
rect 117372 150736 117378 150748
rect 118602 150736 118608 150748
rect 117372 150708 118608 150736
rect 117372 150696 117378 150708
rect 118602 150696 118608 150708
rect 118660 150696 118666 150748
rect 3418 150628 3424 150680
rect 3476 150668 3482 150680
rect 115106 150668 115112 150680
rect 3476 150640 115112 150668
rect 3476 150628 3482 150640
rect 115106 150628 115112 150640
rect 115164 150628 115170 150680
rect 105633 150603 105691 150609
rect 105633 150569 105645 150603
rect 105679 150600 105691 150603
rect 119522 150600 119528 150612
rect 105679 150572 119528 150600
rect 105679 150569 105691 150572
rect 105633 150563 105691 150569
rect 119522 150560 119528 150572
rect 119580 150560 119586 150612
rect 91925 150535 91983 150541
rect 91925 150501 91937 150535
rect 91971 150532 91983 150535
rect 113358 150532 113364 150544
rect 91971 150504 113364 150532
rect 91971 150501 91983 150504
rect 91925 150495 91983 150501
rect 113358 150492 113364 150504
rect 113416 150492 113422 150544
rect 88337 150467 88395 150473
rect 88337 150433 88349 150467
rect 88383 150464 88395 150467
rect 117222 150464 117228 150476
rect 88383 150436 117228 150464
rect 88383 150433 88395 150436
rect 88337 150427 88395 150433
rect 117222 150424 117228 150436
rect 117280 150424 117286 150476
rect 3786 150356 3792 150408
rect 3844 150396 3850 150408
rect 112530 150396 112536 150408
rect 3844 150368 112536 150396
rect 3844 150356 3850 150368
rect 112530 150356 112536 150368
rect 112588 150356 112594 150408
rect 4062 150288 4068 150340
rect 4120 150328 4126 150340
rect 115842 150328 115848 150340
rect 4120 150300 115848 150328
rect 4120 150288 4126 150300
rect 115842 150288 115848 150300
rect 115900 150288 115906 150340
rect 3970 150220 3976 150272
rect 4028 150260 4034 150272
rect 115750 150260 115756 150272
rect 4028 150232 115756 150260
rect 4028 150220 4034 150232
rect 115750 150220 115756 150232
rect 115808 150220 115814 150272
rect 3510 147636 3516 147688
rect 3568 147676 3574 147688
rect 5166 147676 5172 147688
rect 3568 147648 5172 147676
rect 3568 147636 3574 147648
rect 5166 147636 5172 147648
rect 5224 147636 5230 147688
rect 113358 147568 113364 147620
rect 113416 147608 113422 147620
rect 117314 147608 117320 147620
rect 113416 147580 117320 147608
rect 113416 147568 113422 147580
rect 117314 147568 117320 147580
rect 117372 147568 117378 147620
rect 3602 145936 3608 145988
rect 3660 145976 3666 145988
rect 4154 145976 4160 145988
rect 3660 145948 4160 145976
rect 3660 145936 3666 145948
rect 4154 145936 4160 145948
rect 4212 145936 4218 145988
rect 3510 140768 3516 140820
rect 3568 140808 3574 140820
rect 4798 140808 4804 140820
rect 3568 140780 4804 140808
rect 3568 140768 3574 140780
rect 4798 140768 4804 140780
rect 4856 140768 4862 140820
rect 115382 136552 115388 136604
rect 115440 136592 115446 136604
rect 117682 136592 117688 136604
rect 115440 136564 117688 136592
rect 115440 136552 115446 136564
rect 117682 136552 117688 136564
rect 117740 136552 117746 136604
rect 115382 129752 115388 129804
rect 115440 129792 115446 129804
rect 117314 129792 117320 129804
rect 115440 129764 117320 129792
rect 115440 129752 115446 129764
rect 117314 129752 117320 129764
rect 117372 129752 117378 129804
rect 114922 127984 114928 128036
rect 114980 128024 114986 128036
rect 117774 128024 117780 128036
rect 114980 127996 117780 128024
rect 114980 127984 114986 127996
rect 117774 127984 117780 127996
rect 117832 127984 117838 128036
rect 115566 124176 115572 124228
rect 115624 124216 115630 124228
rect 117314 124216 117320 124228
rect 115624 124188 117320 124216
rect 115624 124176 115630 124188
rect 117314 124176 117320 124188
rect 117372 124176 117378 124228
rect 114186 111800 114192 111852
rect 114244 111840 114250 111852
rect 117866 111840 117872 111852
rect 114244 111812 117872 111840
rect 114244 111800 114250 111812
rect 117866 111800 117872 111812
rect 117924 111800 117930 111852
rect 115014 104796 115020 104848
rect 115072 104836 115078 104848
rect 117498 104836 117504 104848
rect 115072 104808 117504 104836
rect 115072 104796 115078 104808
rect 117498 104796 117504 104808
rect 117556 104796 117562 104848
rect 112714 102756 112720 102808
rect 112772 102796 112778 102808
rect 117682 102796 117688 102808
rect 112772 102768 117688 102796
rect 112772 102756 112778 102768
rect 117682 102756 117688 102768
rect 117740 102756 117746 102808
rect 116302 99424 116308 99476
rect 116360 99464 116366 99476
rect 119706 99464 119712 99476
rect 116360 99436 119712 99464
rect 116360 99424 116366 99436
rect 119706 99424 119712 99436
rect 119764 99424 119770 99476
rect 112622 99288 112628 99340
rect 112680 99328 112686 99340
rect 115106 99328 115112 99340
rect 112680 99300 115112 99328
rect 112680 99288 112686 99300
rect 115106 99288 115112 99300
rect 115164 99288 115170 99340
rect 115014 96568 115020 96620
rect 115072 96608 115078 96620
rect 117498 96608 117504 96620
rect 115072 96580 117504 96608
rect 115072 96568 115078 96580
rect 117498 96568 117504 96580
rect 117556 96568 117562 96620
rect 115106 95140 115112 95192
rect 115164 95180 115170 95192
rect 117866 95180 117872 95192
rect 115164 95152 117872 95180
rect 115164 95140 115170 95152
rect 117866 95140 117872 95152
rect 117924 95140 117930 95192
rect 114370 88816 114376 88868
rect 114428 88856 114434 88868
rect 118602 88856 118608 88868
rect 114428 88828 118608 88856
rect 114428 88816 114434 88828
rect 118602 88816 118608 88828
rect 118660 88816 118666 88868
rect 115842 86912 115848 86964
rect 115900 86952 115906 86964
rect 117314 86952 117320 86964
rect 115900 86924 117320 86952
rect 115900 86912 115906 86924
rect 117314 86912 117320 86924
rect 117372 86912 117378 86964
rect 112530 85008 112536 85060
rect 112588 85048 112594 85060
rect 117774 85048 117780 85060
rect 112588 85020 117780 85048
rect 112588 85008 112594 85020
rect 117774 85008 117780 85020
rect 117832 85008 117838 85060
rect 115750 84124 115756 84176
rect 115808 84164 115814 84176
rect 117314 84164 117320 84176
rect 115808 84136 117320 84164
rect 115808 84124 115814 84136
rect 117314 84124 117320 84136
rect 117372 84124 117378 84176
rect 114278 73108 114284 73160
rect 114336 73148 114342 73160
rect 117314 73148 117320 73160
rect 114336 73120 117320 73148
rect 114336 73108 114342 73120
rect 117314 73108 117320 73120
rect 117372 73108 117378 73160
rect 112438 67532 112444 67584
rect 112496 67572 112502 67584
rect 117314 67572 117320 67584
rect 112496 67544 117320 67572
rect 112496 67532 112502 67544
rect 117314 67532 117320 67544
rect 117372 67532 117378 67584
rect 116302 67396 116308 67448
rect 116360 67436 116366 67448
rect 119890 67436 119896 67448
rect 116360 67408 119896 67436
rect 116360 67396 116366 67408
rect 119890 67396 119896 67408
rect 119948 67396 119954 67448
rect 115750 58828 115756 58880
rect 115808 58868 115814 58880
rect 117866 58868 117872 58880
rect 115808 58840 117872 58868
rect 115808 58828 115814 58840
rect 117866 58828 117872 58840
rect 117924 58828 117930 58880
rect 115842 56176 115848 56228
rect 115900 56216 115906 56228
rect 117314 56216 117320 56228
rect 115900 56188 117320 56216
rect 115900 56176 115906 56188
rect 117314 56176 117320 56188
rect 117372 56176 117378 56228
rect 115106 53796 115112 53848
rect 115164 53836 115170 53848
rect 118602 53836 118608 53848
rect 115164 53808 118608 53836
rect 115164 53796 115170 53808
rect 118602 53796 118608 53808
rect 118660 53796 118666 53848
rect 522574 52368 522580 52420
rect 522632 52408 522638 52420
rect 578237 52411 578295 52417
rect 578237 52408 578249 52411
rect 522632 52380 578249 52408
rect 522632 52368 522638 52380
rect 578237 52377 578249 52380
rect 578283 52377 578295 52411
rect 578237 52371 578295 52377
rect 117406 48328 117412 48340
rect 114572 48300 117412 48328
rect 114278 48220 114284 48272
rect 114336 48260 114342 48272
rect 114572 48260 114600 48300
rect 117406 48288 117412 48300
rect 117464 48288 117470 48340
rect 114336 48232 114600 48260
rect 114336 48220 114342 48232
rect 117314 46968 117320 46980
rect 114572 46940 117320 46968
rect 114462 46860 114468 46912
rect 114520 46900 114526 46912
rect 114572 46900 114600 46940
rect 117314 46928 117320 46940
rect 117372 46928 117378 46980
rect 114520 46872 114600 46900
rect 114520 46860 114526 46872
rect 114370 45704 114376 45756
rect 114428 45744 114434 45756
rect 117314 45744 117320 45756
rect 114428 45716 117320 45744
rect 114428 45704 114434 45716
rect 117314 45704 117320 45716
rect 117372 45704 117378 45756
rect 115014 39448 115020 39500
rect 115072 39488 115078 39500
rect 118510 39488 118516 39500
rect 115072 39460 118516 39488
rect 115072 39448 115078 39460
rect 118510 39448 118516 39460
rect 118568 39448 118574 39500
rect 117314 37312 117320 37324
rect 114572 37284 117320 37312
rect 113726 37204 113732 37256
rect 113784 37244 113790 37256
rect 114572 37244 114600 37284
rect 117314 37272 117320 37284
rect 117372 37272 117378 37324
rect 113784 37216 114600 37244
rect 113784 37204 113790 37216
rect 114830 34552 114836 34604
rect 114888 34592 114894 34604
rect 117866 34592 117872 34604
rect 114888 34564 117872 34592
rect 114888 34552 114894 34564
rect 117866 34552 117872 34564
rect 117924 34552 117930 34604
rect 114922 34484 114928 34536
rect 114980 34524 114986 34536
rect 117222 34524 117228 34536
rect 114980 34496 117228 34524
rect 114980 34484 114986 34496
rect 117222 34484 117228 34496
rect 117280 34484 117286 34536
rect 3694 33804 3700 33856
rect 3752 33844 3758 33856
rect 4798 33844 4804 33856
rect 3752 33816 4804 33844
rect 3752 33804 3758 33816
rect 4798 33804 4804 33816
rect 4856 33804 4862 33856
rect 3786 31016 3792 31068
rect 3844 31056 3850 31068
rect 4890 31056 4896 31068
rect 3844 31028 4896 31056
rect 3844 31016 3850 31028
rect 4890 31016 4896 31028
rect 4948 31016 4954 31068
rect 114738 30336 114744 30388
rect 114796 30376 114802 30388
rect 117314 30376 117320 30388
rect 114796 30348 117320 30376
rect 114796 30336 114802 30348
rect 117314 30336 117320 30348
rect 117372 30336 117378 30388
rect 112530 29520 112536 29572
rect 112588 29560 112594 29572
rect 114830 29560 114836 29572
rect 112588 29532 114836 29560
rect 112588 29520 112594 29532
rect 114830 29520 114836 29532
rect 114888 29520 114894 29572
rect 112438 29452 112444 29504
rect 112496 29492 112502 29504
rect 114922 29492 114928 29504
rect 112496 29464 114928 29492
rect 112496 29452 112502 29464
rect 114922 29452 114928 29464
rect 114980 29452 114986 29504
rect 4062 28908 4068 28960
rect 4120 28948 4126 28960
rect 4982 28948 4988 28960
rect 4120 28920 4988 28948
rect 4120 28908 4126 28920
rect 4982 28908 4988 28920
rect 5040 28908 5046 28960
rect 116486 20816 116492 20868
rect 116544 20856 116550 20868
rect 119890 20856 119896 20868
rect 116544 20828 119896 20856
rect 116544 20816 116550 20828
rect 119890 20816 119896 20828
rect 119948 20816 119954 20868
rect 3970 20612 3976 20664
rect 4028 20652 4034 20664
rect 5074 20652 5080 20664
rect 4028 20624 5080 20652
rect 4028 20612 4034 20624
rect 5074 20612 5080 20624
rect 5132 20612 5138 20664
rect 3418 19252 3424 19304
rect 3476 19292 3482 19304
rect 5166 19292 5172 19304
rect 3476 19264 5172 19292
rect 3476 19252 3482 19264
rect 5166 19252 5172 19264
rect 5224 19252 5230 19304
rect 114830 16600 114836 16652
rect 114888 16640 114894 16652
rect 117498 16640 117504 16652
rect 114888 16612 117504 16640
rect 114888 16600 114894 16612
rect 117498 16600 117504 16612
rect 117556 16600 117562 16652
rect 114738 13812 114744 13864
rect 114796 13852 114802 13864
rect 117314 13852 117320 13864
rect 114796 13824 117320 13852
rect 114796 13812 114802 13824
rect 117314 13812 117320 13824
rect 117372 13812 117378 13864
rect 3510 11840 3516 11892
rect 3568 11880 3574 11892
rect 5258 11880 5264 11892
rect 3568 11852 5264 11880
rect 3568 11840 3574 11852
rect 5258 11840 5264 11852
rect 5316 11840 5322 11892
rect 117958 11704 117964 11756
rect 118016 11744 118022 11756
rect 118326 11744 118332 11756
rect 118016 11716 118332 11744
rect 118016 11704 118022 11716
rect 118326 11704 118332 11716
rect 118384 11704 118390 11756
rect 3602 11636 3608 11688
rect 3660 11676 3666 11688
rect 3878 11676 3884 11688
rect 3660 11648 3884 11676
rect 3660 11636 3666 11648
rect 3878 11636 3884 11648
rect 3936 11636 3942 11688
rect 114646 11024 114652 11076
rect 114704 11064 114710 11076
rect 117314 11064 117320 11076
rect 114704 11036 117320 11064
rect 114704 11024 114710 11036
rect 117314 11024 117320 11036
rect 117372 11024 117378 11076
rect 3326 9596 3332 9648
rect 3384 9636 3390 9648
rect 5442 9636 5448 9648
rect 3384 9608 5448 9636
rect 3384 9596 3390 9608
rect 5442 9596 5448 9608
rect 5500 9596 5506 9648
rect 114554 7216 114560 7268
rect 114612 7256 114618 7268
rect 117314 7256 117320 7268
rect 114612 7228 117320 7256
rect 114612 7216 114618 7228
rect 117314 7216 117320 7228
rect 117372 7216 117378 7268
rect 3510 6468 3516 6520
rect 3568 6508 3574 6520
rect 4338 6508 4344 6520
rect 3568 6480 4344 6508
rect 3568 6468 3574 6480
rect 4338 6468 4344 6480
rect 4396 6468 4402 6520
rect 2866 5856 2872 5908
rect 2924 5896 2930 5908
rect 118602 5896 118608 5908
rect 2924 5868 118608 5896
rect 2924 5856 2930 5868
rect 118602 5856 118608 5868
rect 118660 5856 118666 5908
rect 2958 5788 2964 5840
rect 3016 5828 3022 5840
rect 118510 5828 118516 5840
rect 3016 5800 118516 5828
rect 3016 5788 3022 5800
rect 118510 5788 118516 5800
rect 118568 5788 118574 5840
rect 3694 5720 3700 5772
rect 3752 5760 3758 5772
rect 117866 5760 117872 5772
rect 3752 5732 117872 5760
rect 3752 5720 3758 5732
rect 117866 5720 117872 5732
rect 117924 5720 117930 5772
rect 3142 5652 3148 5704
rect 3200 5692 3206 5704
rect 117130 5692 117136 5704
rect 3200 5664 117136 5692
rect 3200 5652 3206 5664
rect 117130 5652 117136 5664
rect 117188 5652 117194 5704
rect 3878 5584 3884 5636
rect 3936 5624 3942 5636
rect 117774 5624 117780 5636
rect 3936 5596 117780 5624
rect 3936 5584 3942 5596
rect 117774 5584 117780 5596
rect 117832 5584 117838 5636
rect 3050 5516 3056 5568
rect 3108 5556 3114 5568
rect 114922 5556 114928 5568
rect 3108 5528 114928 5556
rect 3108 5516 3114 5528
rect 114922 5516 114928 5528
rect 114980 5516 114986 5568
rect 3418 5448 3424 5500
rect 3476 5488 3482 5500
rect 114738 5488 114744 5500
rect 3476 5460 114744 5488
rect 3476 5448 3482 5460
rect 114738 5448 114744 5460
rect 114796 5448 114802 5500
rect 3234 5380 3240 5432
rect 3292 5420 3298 5432
rect 114554 5420 114560 5432
rect 3292 5392 114560 5420
rect 3292 5380 3298 5392
rect 114554 5380 114560 5392
rect 114612 5380 114618 5432
rect 4798 5312 4804 5364
rect 4856 5352 4862 5364
rect 115750 5352 115756 5364
rect 4856 5324 115756 5352
rect 4856 5312 4862 5324
rect 115750 5312 115756 5324
rect 115808 5312 115814 5364
rect 4062 5244 4068 5296
rect 4120 5284 4126 5296
rect 114830 5284 114836 5296
rect 4120 5256 114836 5284
rect 4120 5244 4126 5256
rect 114830 5244 114836 5256
rect 114888 5244 114894 5296
rect 117038 5244 117044 5296
rect 117096 5284 117102 5296
rect 520918 5284 520924 5296
rect 117096 5256 520924 5284
rect 117096 5244 117102 5256
rect 520918 5244 520924 5256
rect 520976 5244 520982 5296
rect 3970 5176 3976 5228
rect 4028 5216 4034 5228
rect 114646 5216 114652 5228
rect 4028 5188 114652 5216
rect 4028 5176 4034 5188
rect 114646 5176 114652 5188
rect 114704 5176 114710 5228
rect 5166 5108 5172 5160
rect 5224 5148 5230 5160
rect 115842 5148 115848 5160
rect 5224 5120 115848 5148
rect 5224 5108 5230 5120
rect 115842 5108 115848 5120
rect 115900 5108 115906 5160
rect 119890 5108 119896 5160
rect 119948 5148 119954 5160
rect 444377 5151 444435 5157
rect 444377 5148 444389 5151
rect 119948 5120 444389 5148
rect 119948 5108 119954 5120
rect 444377 5117 444389 5120
rect 444423 5117 444435 5151
rect 444377 5111 444435 5117
rect 463329 5151 463387 5157
rect 463329 5117 463341 5151
rect 463375 5148 463387 5151
rect 576854 5148 576860 5160
rect 463375 5120 576860 5148
rect 463375 5117 463387 5120
rect 463329 5111 463387 5117
rect 576854 5108 576860 5120
rect 576912 5108 576918 5160
rect 95973 5083 96031 5089
rect 95973 5049 95985 5083
rect 96019 5080 96031 5083
rect 520734 5080 520740 5092
rect 96019 5052 520740 5080
rect 96019 5049 96031 5052
rect 95973 5043 96031 5049
rect 520734 5040 520740 5052
rect 520792 5040 520798 5092
rect 79321 5015 79379 5021
rect 79321 4981 79333 5015
rect 79367 5012 79379 5015
rect 521838 5012 521844 5024
rect 79367 4984 521844 5012
rect 79367 4981 79379 4984
rect 79321 4975 79379 4981
rect 521838 4972 521844 4984
rect 521896 4972 521902 5024
rect 4890 4904 4896 4956
rect 4948 4944 4954 4956
rect 115106 4944 115112 4956
rect 4948 4916 115112 4944
rect 4948 4904 4954 4916
rect 115106 4904 115112 4916
rect 115164 4904 115170 4956
rect 118694 4904 118700 4956
rect 118752 4944 118758 4956
rect 577222 4944 577228 4956
rect 118752 4916 577228 4944
rect 118752 4904 118758 4916
rect 577222 4904 577228 4916
rect 577280 4904 577286 4956
rect 62669 4879 62727 4885
rect 62669 4845 62681 4879
rect 62715 4876 62727 4879
rect 522022 4876 522028 4888
rect 62715 4848 522028 4876
rect 62715 4845 62727 4848
rect 62669 4839 62727 4845
rect 522022 4836 522028 4848
rect 522080 4836 522086 4888
rect 12161 4811 12219 4817
rect 12161 4777 12173 4811
rect 12207 4808 12219 4811
rect 522390 4808 522396 4820
rect 12207 4780 522396 4808
rect 12207 4777 12219 4780
rect 12161 4771 12219 4777
rect 522390 4768 522396 4780
rect 522448 4768 522454 4820
rect 3602 4700 3608 4752
rect 3660 4740 3666 4752
rect 113726 4740 113732 4752
rect 3660 4712 113732 4740
rect 3660 4700 3666 4712
rect 113726 4700 113732 4712
rect 113784 4700 113790 4752
rect 5074 4632 5080 4684
rect 5132 4672 5138 4684
rect 114462 4672 114468 4684
rect 5132 4644 114468 4672
rect 5132 4632 5138 4644
rect 114462 4632 114468 4644
rect 114520 4632 114526 4684
rect 444374 4672 444380 4684
rect 444335 4644 444380 4672
rect 444374 4632 444380 4644
rect 444432 4632 444438 4684
rect 463326 4672 463332 4684
rect 463287 4644 463332 4672
rect 463326 4632 463332 4644
rect 463384 4632 463390 4684
rect 5258 4564 5264 4616
rect 5316 4604 5322 4616
rect 114278 4604 114284 4616
rect 5316 4576 114284 4604
rect 5316 4564 5322 4576
rect 114278 4564 114284 4576
rect 114336 4564 114342 4616
rect 4338 4496 4344 4548
rect 4396 4536 4402 4548
rect 114370 4536 114376 4548
rect 4396 4508 114376 4536
rect 4396 4496 4402 4508
rect 114370 4496 114376 4508
rect 114428 4496 114434 4548
rect 12158 4468 12164 4480
rect 12119 4440 12164 4468
rect 12158 4428 12164 4440
rect 12216 4428 12222 4480
rect 48222 4428 48228 4480
rect 48280 4468 48286 4480
rect 118418 4468 118424 4480
rect 48280 4440 118424 4468
rect 48280 4428 48286 4440
rect 118418 4428 118424 4440
rect 118476 4428 118482 4480
rect 62666 4400 62672 4412
rect 62627 4372 62672 4400
rect 62666 4360 62672 4372
rect 62724 4360 62730 4412
rect 71958 4360 71964 4412
rect 72016 4400 72022 4412
rect 74902 4400 74908 4412
rect 72016 4372 74908 4400
rect 72016 4360 72022 4372
rect 74902 4360 74908 4372
rect 74960 4360 74966 4412
rect 79318 4400 79324 4412
rect 79279 4372 79324 4400
rect 79318 4360 79324 4372
rect 79376 4360 79382 4412
rect 82170 4360 82176 4412
rect 82228 4400 82234 4412
rect 82814 4400 82820 4412
rect 82228 4372 82820 4400
rect 82228 4360 82234 4372
rect 82814 4360 82820 4372
rect 82872 4360 82878 4412
rect 85942 4360 85948 4412
rect 86000 4400 86006 4412
rect 116670 4400 116676 4412
rect 86000 4372 116676 4400
rect 86000 4360 86006 4372
rect 116670 4360 116676 4372
rect 116728 4360 116734 4412
rect 81986 4292 81992 4344
rect 82044 4332 82050 4344
rect 86402 4332 86408 4344
rect 82044 4304 86408 4332
rect 82044 4292 82050 4304
rect 86402 4292 86408 4304
rect 86460 4292 86466 4344
rect 95970 4332 95976 4344
rect 95931 4304 95976 4332
rect 95970 4292 95976 4304
rect 96028 4292 96034 4344
rect 106182 4292 106188 4344
rect 106240 4332 106246 4344
rect 118234 4332 118240 4344
rect 106240 4304 118240 4332
rect 106240 4292 106246 4304
rect 118234 4292 118240 4304
rect 118292 4292 118298 4344
rect 3326 4224 3332 4276
rect 3384 4264 3390 4276
rect 112438 4264 112444 4276
rect 3384 4236 112444 4264
rect 3384 4224 3390 4236
rect 112438 4224 112444 4236
rect 112496 4224 112502 4276
rect 2958 4156 2964 4208
rect 3016 4196 3022 4208
rect 117314 4196 117320 4208
rect 3016 4168 117320 4196
rect 3016 4156 3022 4168
rect 117314 4156 117320 4168
rect 117372 4156 117378 4208
rect 45922 4088 45928 4140
rect 45980 4128 45986 4140
rect 522206 4128 522212 4140
rect 45980 4100 522212 4128
rect 45980 4088 45986 4100
rect 522206 4088 522212 4100
rect 522264 4088 522270 4140
rect 61102 4020 61108 4072
rect 61160 4060 61166 4072
rect 111794 4060 111800 4072
rect 61160 4032 111800 4060
rect 61160 4020 61166 4032
rect 111794 4020 111800 4032
rect 111852 4020 111858 4072
rect 114278 4020 114284 4072
rect 114336 4060 114342 4072
rect 176746 4060 176752 4072
rect 114336 4032 176752 4060
rect 114336 4020 114342 4032
rect 176746 4020 176752 4032
rect 176804 4020 176810 4072
rect 383286 4020 383292 4072
rect 383344 4060 383350 4072
rect 460106 4060 460112 4072
rect 383344 4032 460112 4060
rect 383344 4020 383350 4032
rect 460106 4020 460112 4032
rect 460164 4020 460170 4072
rect 103606 3952 103612 4004
rect 103664 3992 103670 4004
rect 167362 3992 167368 4004
rect 103664 3964 167368 3992
rect 103664 3952 103670 3964
rect 167362 3952 167368 3964
rect 167420 3952 167426 4004
rect 367922 3952 367928 4004
rect 367980 3992 367986 4004
rect 433518 3992 433524 4004
rect 367980 3964 433524 3992
rect 367980 3952 367986 3964
rect 433518 3952 433524 3964
rect 433576 3952 433582 4004
rect 93026 3884 93032 3936
rect 93084 3924 93090 3936
rect 165522 3924 165528 3936
rect 93084 3896 165528 3924
rect 93084 3884 93090 3896
rect 165522 3884 165528 3896
rect 165580 3884 165586 3936
rect 172790 3884 172796 3936
rect 172848 3924 172854 3936
rect 216812 3924 216818 3936
rect 172848 3896 216818 3924
rect 172848 3884 172854 3896
rect 216812 3884 216818 3896
rect 216870 3884 216876 3936
rect 268562 3884 268568 3936
rect 268620 3924 268626 3936
rect 272196 3924 272202 3936
rect 268620 3896 272202 3924
rect 268620 3884 268626 3896
rect 272196 3884 272202 3896
rect 272254 3884 272260 3936
rect 273898 3884 273904 3936
rect 273956 3924 273962 3936
rect 275324 3924 275330 3936
rect 273956 3896 275330 3924
rect 273956 3884 273962 3896
rect 275324 3884 275330 3896
rect 275382 3884 275388 3936
rect 281488 3884 281494 3936
rect 281546 3924 281552 3936
rect 284570 3924 284576 3936
rect 281546 3896 284576 3924
rect 281546 3884 281552 3896
rect 284570 3884 284576 3896
rect 284628 3884 284634 3936
rect 379928 3884 379934 3936
rect 379986 3924 379992 3936
rect 454770 3924 454776 3936
rect 379986 3896 454776 3924
rect 379986 3884 379992 3896
rect 454770 3884 454776 3896
rect 454828 3884 454834 3936
rect 82354 3816 82360 3868
rect 82412 3856 82418 3868
rect 156506 3856 156512 3868
rect 82412 3828 156512 3856
rect 82412 3816 82418 3828
rect 156506 3816 156512 3828
rect 156564 3816 156570 3868
rect 188798 3816 188804 3868
rect 188856 3856 188862 3868
rect 225782 3856 225788 3868
rect 188856 3828 225788 3856
rect 188856 3816 188862 3828
rect 225782 3816 225788 3828
rect 225840 3816 225846 3868
rect 361390 3816 361396 3868
rect 361448 3856 361454 3868
rect 422846 3856 422852 3868
rect 361448 3828 422852 3856
rect 361448 3816 361454 3828
rect 422846 3816 422852 3828
rect 422904 3816 422910 3868
rect 427814 3816 427820 3868
rect 427872 3856 427878 3868
rect 555878 3856 555884 3868
rect 427872 3828 555884 3856
rect 427872 3816 427878 3828
rect 555878 3816 555884 3828
rect 555936 3816 555942 3868
rect 87690 3748 87696 3800
rect 87748 3788 87754 3800
rect 162762 3788 162768 3800
rect 87748 3760 162768 3788
rect 87748 3748 87754 3760
rect 162762 3748 162768 3760
rect 162820 3748 162826 3800
rect 183462 3748 183468 3800
rect 183520 3788 183526 3800
rect 222654 3788 222660 3800
rect 183520 3760 222660 3788
rect 183520 3748 183526 3760
rect 222654 3748 222660 3760
rect 222712 3748 222718 3800
rect 371050 3748 371056 3800
rect 371108 3788 371114 3800
rect 438854 3788 438860 3800
rect 371108 3760 438860 3788
rect 371108 3748 371114 3760
rect 438854 3748 438860 3760
rect 438912 3748 438918 3800
rect 444190 3788 444196 3800
rect 441586 3760 444196 3788
rect 77018 3680 77024 3732
rect 77076 3720 77082 3732
rect 153102 3720 153108 3732
rect 77076 3692 153108 3720
rect 77076 3680 77082 3692
rect 153102 3680 153108 3692
rect 153160 3680 153166 3732
rect 178126 3680 178132 3732
rect 178184 3720 178190 3732
rect 219618 3720 219624 3732
rect 178184 3692 219624 3720
rect 178184 3680 178190 3692
rect 219618 3680 219624 3692
rect 219676 3680 219682 3732
rect 373902 3680 373908 3732
rect 373960 3720 373966 3732
rect 441586 3720 441614 3760
rect 444190 3748 444196 3760
rect 444248 3748 444254 3800
rect 454678 3748 454684 3800
rect 454736 3788 454742 3800
rect 534626 3788 534632 3800
rect 454736 3760 534632 3788
rect 454736 3748 454742 3760
rect 534626 3748 534632 3760
rect 534684 3748 534690 3800
rect 373960 3692 441614 3720
rect 373960 3680 373966 3692
rect 443730 3680 443736 3732
rect 443788 3720 443794 3732
rect 539962 3720 539968 3732
rect 443788 3692 539968 3720
rect 443788 3680 443794 3692
rect 539962 3680 539968 3692
rect 540020 3680 540026 3732
rect 71682 3612 71688 3664
rect 71740 3652 71746 3664
rect 149146 3652 149152 3664
rect 71740 3624 149152 3652
rect 71740 3612 71746 3624
rect 149146 3612 149152 3624
rect 149204 3612 149210 3664
rect 167454 3612 167460 3664
rect 167512 3652 167518 3664
rect 213454 3652 213460 3664
rect 167512 3624 213460 3652
rect 167512 3612 167518 3624
rect 213454 3612 213460 3624
rect 213512 3612 213518 3664
rect 324866 3612 324872 3664
rect 324924 3652 324930 3664
rect 358998 3652 359004 3664
rect 324924 3624 359004 3652
rect 324924 3612 324930 3624
rect 358998 3612 359004 3624
rect 359056 3612 359062 3664
rect 386322 3612 386328 3664
rect 386380 3652 386386 3664
rect 465442 3652 465448 3664
rect 386380 3624 465448 3652
rect 386380 3612 386386 3624
rect 465442 3612 465448 3624
rect 465500 3612 465506 3664
rect 66438 3544 66444 3596
rect 66496 3584 66502 3596
rect 146110 3584 146116 3596
rect 66496 3556 146116 3584
rect 66496 3544 66502 3556
rect 146110 3544 146116 3556
rect 146168 3544 146174 3596
rect 162210 3544 162216 3596
rect 162268 3584 162274 3596
rect 210326 3584 210332 3596
rect 162268 3556 210332 3584
rect 162268 3544 162274 3556
rect 210326 3544 210332 3556
rect 210384 3544 210390 3596
rect 318702 3544 318708 3596
rect 318760 3584 318766 3596
rect 348418 3584 348424 3596
rect 318760 3556 348424 3584
rect 318760 3544 318766 3556
rect 348418 3544 348424 3556
rect 348476 3544 348482 3596
rect 389082 3544 389088 3596
rect 389140 3584 389146 3596
rect 470778 3584 470784 3596
rect 389140 3556 470784 3584
rect 389140 3544 389146 3556
rect 470778 3544 470784 3556
rect 470836 3544 470842 3596
rect 55950 3476 55956 3528
rect 56008 3516 56014 3528
rect 118050 3516 118056 3528
rect 56008 3488 118056 3516
rect 56008 3476 56014 3488
rect 118050 3476 118056 3488
rect 118108 3476 118114 3528
rect 151538 3476 151544 3528
rect 151596 3516 151602 3528
rect 204254 3516 204260 3528
rect 151596 3488 204260 3516
rect 151596 3476 151602 3488
rect 204254 3476 204260 3488
rect 204312 3476 204318 3528
rect 343358 3476 343364 3528
rect 343416 3516 343422 3528
rect 390922 3516 390928 3528
rect 343416 3488 390928 3516
rect 343416 3476 343422 3488
rect 390922 3476 390928 3488
rect 390980 3476 390986 3528
rect 392578 3476 392584 3528
rect 392636 3516 392642 3528
rect 476114 3516 476120 3528
rect 392636 3488 476120 3516
rect 392636 3476 392642 3488
rect 476114 3476 476120 3488
rect 476172 3476 476178 3528
rect 98362 3408 98368 3460
rect 98420 3448 98426 3460
rect 173434 3448 173440 3460
rect 98420 3420 173440 3448
rect 98420 3408 98426 3420
rect 173434 3408 173440 3420
rect 173492 3408 173498 3460
rect 337194 3408 337200 3460
rect 337252 3448 337258 3460
rect 380342 3448 380348 3460
rect 337252 3420 380348 3448
rect 337252 3408 337258 3420
rect 380342 3408 380348 3420
rect 380400 3408 380406 3460
rect 395614 3408 395620 3460
rect 395672 3448 395678 3460
rect 481450 3448 481456 3460
rect 395672 3420 481456 3448
rect 395672 3408 395678 3420
rect 481450 3408 481456 3420
rect 481508 3408 481514 3460
rect 522942 3408 522948 3460
rect 523000 3448 523006 3460
rect 566550 3448 566556 3460
rect 523000 3420 566556 3448
rect 523000 3408 523006 3420
rect 566550 3408 566556 3420
rect 566608 3408 566614 3460
rect 42610 3340 42616 3392
rect 42668 3380 42674 3392
rect 117590 3380 117596 3392
rect 42668 3352 117596 3380
rect 42668 3340 42674 3352
rect 117590 3340 117596 3352
rect 117648 3340 117654 3392
rect 119706 3340 119712 3392
rect 119764 3380 119770 3392
rect 130657 3383 130715 3389
rect 130657 3380 130669 3383
rect 119764 3352 130669 3380
rect 119764 3340 119770 3352
rect 130657 3349 130669 3352
rect 130703 3349 130715 3383
rect 130657 3343 130715 3349
rect 146202 3340 146208 3392
rect 146260 3380 146266 3392
rect 201126 3380 201132 3392
rect 146260 3352 201132 3380
rect 146260 3340 146266 3352
rect 201126 3340 201132 3352
rect 201184 3340 201190 3392
rect 204714 3340 204720 3392
rect 204772 3380 204778 3392
rect 234982 3380 234988 3392
rect 204772 3352 234988 3380
rect 204772 3340 204778 3352
rect 234982 3340 234988 3352
rect 235040 3340 235046 3392
rect 247402 3340 247408 3392
rect 247460 3380 247466 3392
rect 259638 3380 259644 3392
rect 247460 3352 259644 3380
rect 247460 3340 247466 3352
rect 259638 3340 259644 3352
rect 259696 3340 259702 3392
rect 309502 3340 309508 3392
rect 309560 3380 309566 3392
rect 332410 3380 332416 3392
rect 309560 3352 332416 3380
rect 309560 3340 309566 3352
rect 332410 3340 332416 3352
rect 332468 3340 332474 3392
rect 352558 3340 352564 3392
rect 352616 3380 352622 3392
rect 404817 3383 404875 3389
rect 404817 3380 404829 3383
rect 352616 3352 404829 3380
rect 352616 3340 352622 3352
rect 404817 3349 404829 3352
rect 404863 3349 404875 3383
rect 404817 3343 404875 3349
rect 404906 3340 404912 3392
rect 404964 3380 404970 3392
rect 407669 3383 407727 3389
rect 407669 3380 407681 3383
rect 404964 3352 407681 3380
rect 404964 3340 404970 3352
rect 407669 3349 407681 3352
rect 407715 3349 407727 3383
rect 407669 3343 407727 3349
rect 407758 3340 407764 3392
rect 407816 3380 407822 3392
rect 486694 3380 486700 3392
rect 407816 3352 486700 3380
rect 407816 3340 407822 3352
rect 486694 3340 486700 3352
rect 486752 3340 486758 3392
rect 29178 3272 29184 3324
rect 29236 3312 29242 3324
rect 136634 3312 136640 3324
rect 29236 3284 136640 3312
rect 29236 3272 29242 3284
rect 136634 3272 136640 3284
rect 136692 3272 136698 3324
rect 140866 3272 140872 3324
rect 140924 3312 140930 3324
rect 198090 3312 198096 3324
rect 140924 3284 198096 3312
rect 140924 3272 140930 3284
rect 198090 3272 198096 3284
rect 198148 3272 198154 3324
rect 199378 3272 199384 3324
rect 199436 3312 199442 3324
rect 231946 3312 231952 3324
rect 199436 3284 231952 3312
rect 199436 3272 199442 3284
rect 231946 3272 231952 3284
rect 232004 3272 232010 3324
rect 358722 3272 358728 3324
rect 358780 3312 358786 3324
rect 417326 3312 417332 3324
rect 358780 3284 417332 3312
rect 358780 3272 358786 3284
rect 417326 3272 417332 3284
rect 417384 3272 417390 3324
rect 417421 3315 417479 3321
rect 417421 3281 417433 3315
rect 417467 3312 417479 3315
rect 492030 3312 492036 3324
rect 417467 3284 492036 3312
rect 417467 3281 417479 3284
rect 417421 3275 417479 3281
rect 492030 3272 492036 3284
rect 492088 3272 492094 3324
rect 518618 3272 518624 3324
rect 518676 3312 518682 3324
rect 520550 3312 520556 3324
rect 518676 3284 520556 3312
rect 518676 3272 518682 3284
rect 520550 3272 520556 3284
rect 520608 3272 520614 3324
rect 23842 3204 23848 3256
rect 23900 3244 23906 3256
rect 133414 3244 133420 3256
rect 23900 3216 133420 3244
rect 23900 3204 23906 3216
rect 133414 3204 133420 3216
rect 133472 3204 133478 3256
rect 135530 3204 135536 3256
rect 135588 3244 135594 3256
rect 194962 3244 194968 3256
rect 135588 3216 194968 3244
rect 135588 3204 135594 3216
rect 194962 3204 194968 3216
rect 195020 3204 195026 3256
rect 226058 3204 226064 3256
rect 226116 3244 226122 3256
rect 247310 3244 247316 3256
rect 226116 3216 247316 3244
rect 226116 3204 226122 3216
rect 247310 3204 247316 3216
rect 247368 3204 247374 3256
rect 306190 3204 306196 3256
rect 306248 3244 306254 3256
rect 327074 3244 327080 3256
rect 306248 3216 327080 3244
rect 306248 3204 306254 3216
rect 327074 3204 327080 3216
rect 327132 3204 327138 3256
rect 331030 3204 331036 3256
rect 331088 3244 331094 3256
rect 369670 3244 369676 3256
rect 331088 3216 369676 3244
rect 331088 3204 331094 3216
rect 369670 3204 369676 3216
rect 369728 3204 369734 3256
rect 398742 3204 398748 3256
rect 398800 3244 398806 3256
rect 407758 3244 407764 3256
rect 398800 3216 407764 3244
rect 398800 3204 398806 3216
rect 407758 3204 407764 3216
rect 407816 3204 407822 3256
rect 407853 3247 407911 3253
rect 407853 3213 407865 3247
rect 407899 3244 407911 3247
rect 497366 3244 497372 3256
rect 407899 3216 497372 3244
rect 407899 3213 407911 3216
rect 407853 3207 407911 3213
rect 497366 3204 497372 3216
rect 497424 3204 497430 3256
rect 18506 3136 18512 3188
rect 18564 3176 18570 3188
rect 130378 3176 130384 3188
rect 18564 3148 130384 3176
rect 18564 3136 18570 3148
rect 130378 3136 130384 3148
rect 130436 3136 130442 3188
rect 191926 3176 191932 3188
rect 130488 3148 191932 3176
rect 13170 3068 13176 3120
rect 13228 3108 13234 3120
rect 127250 3108 127256 3120
rect 13228 3080 127256 3108
rect 13228 3068 13234 3080
rect 127250 3068 127256 3080
rect 127308 3068 127314 3120
rect 130286 3068 130292 3120
rect 130344 3108 130350 3120
rect 130488 3108 130516 3148
rect 191926 3136 191932 3148
rect 191984 3136 191990 3188
rect 215386 3136 215392 3188
rect 215444 3176 215450 3188
rect 241146 3176 241152 3188
rect 215444 3148 241152 3176
rect 215444 3136 215450 3148
rect 241146 3136 241152 3148
rect 241204 3136 241210 3188
rect 333882 3136 333888 3188
rect 333940 3176 333946 3188
rect 375006 3176 375012 3188
rect 333940 3148 375012 3176
rect 333940 3136 333946 3148
rect 375006 3136 375012 3148
rect 375064 3136 375070 3188
rect 404817 3179 404875 3185
rect 404817 3145 404829 3179
rect 404863 3176 404875 3179
rect 406930 3176 406936 3188
rect 404863 3148 406936 3176
rect 404863 3145 404875 3148
rect 404817 3139 404875 3145
rect 406930 3136 406936 3148
rect 406988 3136 406994 3188
rect 407393 3179 407451 3185
rect 407393 3145 407405 3179
rect 407439 3176 407451 3179
rect 417421 3179 417479 3185
rect 417421 3176 417433 3179
rect 407439 3148 417433 3176
rect 407439 3145 407451 3148
rect 407393 3139 407451 3145
rect 417421 3145 417433 3148
rect 417467 3145 417479 3179
rect 417421 3139 417479 3145
rect 417513 3179 417571 3185
rect 417513 3145 417525 3179
rect 417559 3176 417571 3179
rect 502610 3176 502616 3188
rect 417559 3148 502616 3176
rect 417559 3145 417571 3148
rect 417513 3139 417571 3145
rect 502610 3136 502616 3148
rect 502668 3136 502674 3188
rect 189074 3108 189080 3120
rect 130344 3080 130516 3108
rect 130580 3080 189080 3108
rect 130344 3068 130350 3080
rect 7834 3000 7840 3052
rect 7892 3040 7898 3052
rect 124214 3040 124220 3052
rect 7892 3012 124220 3040
rect 7892 3000 7898 3012
rect 124214 3000 124220 3012
rect 124272 3000 124278 3052
rect 2590 2932 2596 2984
rect 2648 2972 2654 2984
rect 121454 2972 121460 2984
rect 2648 2944 121460 2972
rect 2648 2932 2654 2944
rect 121454 2932 121460 2944
rect 121512 2932 121518 2984
rect 124950 2932 124956 2984
rect 125008 2972 125014 2984
rect 130580 2972 130608 3080
rect 189074 3068 189080 3080
rect 189132 3068 189138 3120
rect 210050 3068 210056 3120
rect 210108 3108 210114 3120
rect 238018 3108 238024 3120
rect 210108 3080 238024 3108
rect 210108 3068 210114 3080
rect 238018 3068 238024 3080
rect 238076 3068 238082 3120
rect 241974 3068 241980 3120
rect 242032 3108 242038 3120
rect 256602 3108 256608 3120
rect 242032 3080 256608 3108
rect 242032 3068 242038 3080
rect 256602 3068 256608 3080
rect 256660 3068 256666 3120
rect 321462 3068 321468 3120
rect 321520 3108 321526 3120
rect 353754 3108 353760 3120
rect 321520 3080 353760 3108
rect 321520 3068 321526 3080
rect 353754 3068 353760 3080
rect 353812 3068 353818 3120
rect 364886 3068 364892 3120
rect 364944 3108 364950 3120
rect 428182 3108 428188 3120
rect 364944 3080 428188 3108
rect 364944 3068 364950 3080
rect 428182 3068 428188 3080
rect 428240 3068 428246 3120
rect 438670 3068 438676 3120
rect 438728 3108 438734 3120
rect 550542 3108 550548 3120
rect 438728 3080 550548 3108
rect 438728 3068 438734 3080
rect 550542 3068 550548 3080
rect 550600 3068 550606 3120
rect 185762 3040 185768 3052
rect 132466 3012 185768 3040
rect 125008 2944 130608 2972
rect 130657 2975 130715 2981
rect 125008 2932 125014 2944
rect 130657 2941 130669 2975
rect 130703 2972 130715 2975
rect 132466 2972 132494 3012
rect 185762 3000 185768 3012
rect 185820 3000 185826 3052
rect 231302 3000 231308 3052
rect 231360 3040 231366 3052
rect 250346 3040 250352 3052
rect 231360 3012 250352 3040
rect 231360 3000 231366 3012
rect 250346 3000 250352 3012
rect 250404 3000 250410 3052
rect 257982 3000 257988 3052
rect 258040 3040 258046 3052
rect 265710 3040 265716 3052
rect 258040 3012 265716 3040
rect 258040 3000 258046 3012
rect 265710 3000 265716 3012
rect 265768 3000 265774 3052
rect 312538 3000 312544 3052
rect 312596 3040 312602 3052
rect 337746 3040 337752 3052
rect 312596 3012 337752 3040
rect 312596 3000 312602 3012
rect 337746 3000 337752 3012
rect 337804 3000 337810 3052
rect 340230 3000 340236 3052
rect 340288 3040 340294 3052
rect 385678 3040 385684 3052
rect 340288 3012 385684 3040
rect 340288 3000 340294 3012
rect 385678 3000 385684 3012
rect 385736 3000 385742 3052
rect 401410 3000 401416 3052
rect 401468 3040 401474 3052
rect 407393 3043 407451 3049
rect 407393 3040 407405 3043
rect 401468 3012 407405 3040
rect 401468 3000 401474 3012
rect 407393 3009 407405 3012
rect 407439 3009 407451 3043
rect 407393 3003 407451 3009
rect 407942 3000 407948 3052
rect 408000 3040 408006 3052
rect 417513 3043 417571 3049
rect 417513 3040 417525 3043
rect 408000 3012 417525 3040
rect 408000 3000 408006 3012
rect 417513 3009 417525 3012
rect 417559 3009 417571 3043
rect 417513 3003 417571 3009
rect 423306 3000 423312 3052
rect 423364 3040 423370 3052
rect 561214 3040 561220 3052
rect 423364 3012 561220 3040
rect 423364 3000 423370 3012
rect 561214 3000 561220 3012
rect 561272 3000 561278 3052
rect 130703 2944 132494 2972
rect 130703 2941 130715 2944
rect 130657 2935 130715 2941
rect 156874 2932 156880 2984
rect 156932 2972 156938 2984
rect 207290 2972 207296 2984
rect 156932 2944 207296 2972
rect 156932 2932 156938 2944
rect 207290 2932 207296 2944
rect 207348 2932 207354 2984
rect 220722 2932 220728 2984
rect 220780 2972 220786 2984
rect 244274 2972 244280 2984
rect 220780 2944 244280 2972
rect 220780 2932 220786 2944
rect 244274 2932 244280 2944
rect 244332 2932 244338 2984
rect 252646 2932 252652 2984
rect 252704 2972 252710 2984
rect 262674 2972 262680 2984
rect 252704 2944 262680 2972
rect 252704 2932 252710 2944
rect 262674 2932 262680 2944
rect 262732 2932 262738 2984
rect 315666 2932 315672 2984
rect 315724 2972 315730 2984
rect 343082 2972 343088 2984
rect 315724 2944 343088 2972
rect 315724 2932 315730 2944
rect 343082 2932 343088 2944
rect 343140 2932 343146 2984
rect 346302 2932 346308 2984
rect 346360 2972 346366 2984
rect 396258 2972 396264 2984
rect 346360 2944 396264 2972
rect 346360 2932 346366 2944
rect 396258 2932 396264 2944
rect 396316 2932 396322 2984
rect 426342 2932 426348 2984
rect 426400 2972 426406 2984
rect 571886 2972 571892 2984
rect 426400 2944 571892 2972
rect 426400 2932 426406 2944
rect 571886 2932 571892 2944
rect 571944 2932 571950 2984
rect 45094 2864 45100 2916
rect 45152 2904 45158 2916
rect 50338 2904 50344 2916
rect 45152 2876 50344 2904
rect 45152 2864 45158 2876
rect 50338 2864 50344 2876
rect 50396 2864 50402 2916
rect 52362 2864 52368 2916
rect 52420 2904 52426 2916
rect 522114 2904 522120 2916
rect 52420 2876 522120 2904
rect 52420 2864 52426 2876
rect 522114 2864 522120 2876
rect 522172 2864 522178 2916
rect 34514 2796 34520 2848
rect 34572 2836 34578 2848
rect 44174 2836 44180 2848
rect 34572 2808 44180 2836
rect 34572 2796 34578 2808
rect 44174 2796 44180 2808
rect 44232 2796 44238 2848
rect 108942 2796 108948 2848
rect 109000 2836 109006 2848
rect 179598 2836 179604 2848
rect 109000 2808 179604 2836
rect 109000 2796 109006 2808
rect 179598 2796 179604 2808
rect 179656 2796 179662 2848
rect 194134 2796 194140 2848
rect 194192 2836 194198 2848
rect 229094 2836 229100 2848
rect 194192 2808 229100 2836
rect 194192 2796 194198 2808
rect 229094 2796 229100 2808
rect 229152 2796 229158 2848
rect 236638 2796 236644 2848
rect 236696 2836 236702 2848
rect 236696 2808 248414 2836
rect 236696 2796 236702 2808
rect 19242 2728 19248 2780
rect 19300 2768 19306 2780
rect 106182 2768 106188 2780
rect 19300 2740 106188 2768
rect 19300 2728 19306 2740
rect 106182 2728 106188 2740
rect 106240 2728 106246 2780
rect 111794 2728 111800 2780
rect 111852 2768 111858 2780
rect 151998 2768 152004 2780
rect 111852 2740 152004 2768
rect 111852 2728 111858 2740
rect 151998 2728 152004 2740
rect 152056 2728 152062 2780
rect 153102 2728 153108 2780
rect 153160 2768 153166 2780
rect 161106 2768 161112 2780
rect 153160 2740 161112 2768
rect 153160 2728 153166 2740
rect 161106 2728 161112 2740
rect 161164 2728 161170 2780
rect 164234 2768 164240 2780
rect 161216 2740 164240 2768
rect 28902 2660 28908 2712
rect 28960 2700 28966 2712
rect 119338 2700 119344 2712
rect 28960 2672 119344 2700
rect 28960 2660 28966 2672
rect 119338 2660 119344 2672
rect 119396 2660 119402 2712
rect 156506 2660 156512 2712
rect 156564 2700 156570 2712
rect 161216 2700 161244 2740
rect 164234 2728 164240 2740
rect 164292 2728 164298 2780
rect 165522 2728 165528 2780
rect 165580 2768 165586 2780
rect 170398 2768 170404 2780
rect 165580 2740 170404 2768
rect 165580 2728 165586 2740
rect 170398 2728 170404 2740
rect 170456 2728 170462 2780
rect 176746 2728 176752 2780
rect 176804 2768 176810 2780
rect 182634 2768 182640 2780
rect 176804 2740 182640 2768
rect 176804 2728 176810 2740
rect 182634 2728 182640 2740
rect 182692 2728 182698 2780
rect 248386 2768 248414 2808
rect 263226 2796 263232 2848
rect 263284 2836 263290 2848
rect 289630 2836 289636 2848
rect 263284 2808 267734 2836
rect 263284 2796 263290 2808
rect 253474 2768 253480 2780
rect 248386 2740 253480 2768
rect 253474 2728 253480 2740
rect 253532 2728 253538 2780
rect 267706 2768 267734 2808
rect 287026 2808 289636 2836
rect 269114 2768 269120 2780
rect 267706 2740 269120 2768
rect 269114 2728 269120 2740
rect 269172 2728 269178 2780
rect 284846 2728 284852 2780
rect 284904 2768 284910 2780
rect 287026 2768 287054 2808
rect 289630 2796 289636 2808
rect 289688 2796 289694 2848
rect 295150 2836 295156 2848
rect 289740 2808 295156 2836
rect 284904 2740 287054 2768
rect 284904 2728 284910 2740
rect 287974 2728 287980 2780
rect 288032 2768 288038 2780
rect 289740 2768 289768 2808
rect 295150 2796 295156 2808
rect 295208 2796 295214 2848
rect 303338 2796 303344 2848
rect 303396 2836 303402 2848
rect 321830 2836 321836 2848
rect 303396 2808 321836 2836
rect 303396 2796 303402 2808
rect 321830 2796 321836 2808
rect 321888 2796 321894 2848
rect 327902 2796 327908 2848
rect 327960 2836 327966 2848
rect 364334 2836 364340 2848
rect 327960 2808 364340 2836
rect 327960 2796 327966 2808
rect 364334 2796 364340 2808
rect 364392 2796 364398 2848
rect 377214 2796 377220 2848
rect 377272 2836 377278 2848
rect 449526 2836 449532 2848
rect 377272 2808 449532 2836
rect 377272 2796 377278 2808
rect 449526 2796 449532 2808
rect 449584 2796 449590 2848
rect 484302 2796 484308 2848
rect 484360 2836 484366 2848
rect 523954 2836 523960 2848
rect 484360 2808 523960 2836
rect 484360 2796 484366 2808
rect 523954 2796 523960 2808
rect 524012 2796 524018 2848
rect 288032 2740 289768 2768
rect 288032 2728 288038 2740
rect 417142 2728 417148 2780
rect 417200 2768 417206 2780
rect 454678 2768 454684 2780
rect 417200 2740 454684 2768
rect 417200 2728 417206 2740
rect 454678 2728 454684 2740
rect 454736 2728 454742 2780
rect 156564 2672 161244 2700
rect 156564 2660 156570 2672
rect 162762 2660 162768 2712
rect 162820 2700 162826 2712
rect 167270 2700 167276 2712
rect 162820 2672 167276 2700
rect 162820 2660 162826 2672
rect 167270 2660 167276 2672
rect 167328 2660 167334 2712
rect 167362 2660 167368 2712
rect 167420 2700 167426 2712
rect 176654 2700 176660 2712
rect 167420 2672 176660 2700
rect 167420 2660 167426 2672
rect 176654 2660 176660 2672
rect 176712 2660 176718 2712
rect 420270 2660 420276 2712
rect 420328 2700 420334 2712
rect 427814 2700 427820 2712
rect 420328 2672 427820 2700
rect 420328 2660 420334 2672
rect 427814 2660 427820 2672
rect 427872 2660 427878 2712
rect 435634 2660 435640 2712
rect 435692 2700 435698 2712
rect 443730 2700 443736 2712
rect 435692 2672 443736 2700
rect 435692 2660 435698 2672
rect 443730 2660 443736 2672
rect 443788 2660 443794 2712
rect 1302 2592 1308 2644
rect 1360 2632 1366 2644
rect 58618 2632 58624 2644
rect 1360 2604 58624 2632
rect 1360 2592 1366 2604
rect 58618 2592 58624 2604
rect 58676 2592 58682 2644
rect 75822 2592 75828 2644
rect 75880 2632 75886 2644
rect 499666 2632 499672 2644
rect 75880 2604 499672 2632
rect 75880 2592 75886 2604
rect 499666 2592 499672 2604
rect 499724 2592 499730 2644
rect 5994 2524 6000 2576
rect 6052 2564 6058 2576
rect 48222 2564 48228 2576
rect 6052 2536 48228 2564
rect 6052 2524 6058 2536
rect 48222 2524 48228 2536
rect 48280 2524 48286 2576
rect 68922 2524 68928 2576
rect 68980 2564 68986 2576
rect 490374 2564 490380 2576
rect 68980 2536 490380 2564
rect 68980 2524 68986 2536
rect 490374 2524 490380 2536
rect 490432 2524 490438 2576
rect 89346 2456 89352 2508
rect 89404 2496 89410 2508
rect 502702 2496 502708 2508
rect 89404 2468 502708 2496
rect 89404 2456 89410 2468
rect 502702 2456 502708 2468
rect 502760 2456 502766 2508
rect 92382 2388 92388 2440
rect 92440 2428 92446 2440
rect 505738 2428 505744 2440
rect 92440 2400 505744 2428
rect 92440 2388 92446 2400
rect 505738 2388 505744 2400
rect 505796 2388 505802 2440
rect 108850 2320 108856 2372
rect 108908 2360 108914 2372
rect 520642 2360 520648 2372
rect 108908 2332 520648 2360
rect 108908 2320 108914 2332
rect 520642 2320 520648 2332
rect 520700 2320 520706 2372
rect 112622 2252 112628 2304
rect 112680 2292 112686 2304
rect 520366 2292 520372 2304
rect 112680 2264 520372 2292
rect 112680 2252 112686 2264
rect 520366 2252 520372 2264
rect 520424 2252 520430 2304
rect 105998 2184 106004 2236
rect 106056 2224 106062 2236
rect 511994 2224 512000 2236
rect 106056 2196 512000 2224
rect 106056 2184 106062 2196
rect 511994 2184 512000 2196
rect 512052 2184 512058 2236
rect 22646 2116 22652 2168
rect 22704 2156 22710 2168
rect 108301 2159 108359 2165
rect 108301 2156 108313 2159
rect 22704 2128 108313 2156
rect 22704 2116 22710 2128
rect 108301 2125 108313 2128
rect 108347 2125 108359 2159
rect 108301 2119 108359 2125
rect 113818 2116 113824 2168
rect 113876 2156 113882 2168
rect 114370 2156 114376 2168
rect 113876 2128 114376 2156
rect 113876 2116 113882 2128
rect 114370 2116 114376 2128
rect 114428 2116 114434 2168
rect 115290 2116 115296 2168
rect 115348 2156 115354 2168
rect 115348 2128 115520 2156
rect 115348 2116 115354 2128
rect 32582 2048 32588 2100
rect 32640 2088 32646 2100
rect 115382 2088 115388 2100
rect 32640 2060 115388 2088
rect 32640 2048 32646 2060
rect 115382 2048 115388 2060
rect 115440 2048 115446 2100
rect 115492 2088 115520 2128
rect 119522 2116 119528 2168
rect 119580 2156 119586 2168
rect 515030 2156 515036 2168
rect 119580 2128 515036 2156
rect 119580 2116 119586 2128
rect 515030 2116 515036 2128
rect 515088 2116 515094 2168
rect 508866 2088 508872 2100
rect 115492 2060 508872 2088
rect 508866 2048 508872 2060
rect 508924 2048 508930 2100
rect 44174 1980 44180 2032
rect 44232 2020 44238 2032
rect 432138 2020 432144 2032
rect 44232 1992 432144 2020
rect 44232 1980 44238 1992
rect 432138 1980 432144 1992
rect 432196 1980 432202 2032
rect 9306 1912 9312 1964
rect 9364 1952 9370 1964
rect 114002 1952 114008 1964
rect 9364 1924 114008 1952
rect 9364 1912 9370 1924
rect 114002 1912 114008 1924
rect 114060 1912 114066 1964
rect 114094 1912 114100 1964
rect 114152 1952 114158 1964
rect 114152 1924 115704 1952
rect 114152 1912 114158 1924
rect 108301 1887 108359 1893
rect 108301 1853 108313 1887
rect 108347 1884 108359 1887
rect 115566 1884 115572 1896
rect 108347 1856 115572 1884
rect 108347 1853 108359 1856
rect 108301 1847 108359 1853
rect 115566 1844 115572 1856
rect 115624 1844 115630 1896
rect 99282 1776 99288 1828
rect 99340 1816 99346 1828
rect 114186 1816 114192 1828
rect 99340 1788 114192 1816
rect 99340 1776 99346 1788
rect 114186 1776 114192 1788
rect 114244 1776 114250 1828
rect 114370 1776 114376 1828
rect 114428 1816 114434 1828
rect 115477 1819 115535 1825
rect 115477 1816 115489 1819
rect 114428 1788 115489 1816
rect 114428 1776 114434 1788
rect 115477 1785 115489 1788
rect 115523 1785 115535 1819
rect 115676 1816 115704 1924
rect 116578 1912 116584 1964
rect 116636 1952 116642 1964
rect 496814 1952 496820 1964
rect 116636 1924 496820 1952
rect 116636 1912 116642 1924
rect 496814 1912 496820 1924
rect 496872 1912 496878 1964
rect 115753 1887 115811 1893
rect 115753 1853 115765 1887
rect 115799 1884 115811 1887
rect 493410 1884 493416 1896
rect 115799 1856 493416 1884
rect 115799 1853 115811 1856
rect 115753 1847 115811 1853
rect 493410 1844 493416 1856
rect 493468 1844 493474 1896
rect 487338 1816 487344 1828
rect 115676 1788 487344 1816
rect 115477 1779 115535 1785
rect 487338 1776 487344 1788
rect 487396 1776 487402 1828
rect 39758 1708 39764 1760
rect 39816 1748 39822 1760
rect 139578 1748 139584 1760
rect 39816 1720 139584 1748
rect 39816 1708 39822 1720
rect 139578 1708 139584 1720
rect 139636 1708 139642 1760
rect 149146 1708 149152 1760
rect 149204 1748 149210 1760
rect 158070 1748 158076 1760
rect 149204 1720 158076 1748
rect 149204 1708 149210 1720
rect 158070 1708 158076 1720
rect 158128 1708 158134 1760
rect 278682 1708 278688 1760
rect 278740 1748 278746 1760
rect 279234 1748 279240 1760
rect 278740 1720 279240 1748
rect 278740 1708 278746 1720
rect 279234 1708 279240 1720
rect 279292 1708 279298 1760
rect 291010 1708 291016 1760
rect 291068 1748 291074 1760
rect 300486 1748 300492 1760
rect 291068 1720 300492 1748
rect 291068 1708 291074 1720
rect 300486 1708 300492 1720
rect 300544 1708 300550 1760
rect 316494 1748 316500 1760
rect 303172 1720 316500 1748
rect 50338 1640 50344 1692
rect 50396 1680 50402 1692
rect 142706 1680 142712 1692
rect 50396 1652 142712 1680
rect 50396 1640 50402 1652
rect 142706 1640 142712 1652
rect 142764 1640 142770 1692
rect 146110 1640 146116 1692
rect 146168 1680 146174 1692
rect 154942 1680 154948 1692
rect 146168 1652 154948 1680
rect 146168 1640 146174 1652
rect 154942 1640 154948 1652
rect 155000 1640 155006 1692
rect 300210 1640 300216 1692
rect 300268 1680 300274 1692
rect 303172 1680 303200 1720
rect 316494 1708 316500 1720
rect 316552 1708 316558 1760
rect 349522 1708 349528 1760
rect 349580 1748 349586 1760
rect 401594 1748 401600 1760
rect 349580 1720 401600 1748
rect 349580 1708 349586 1720
rect 401594 1708 401600 1720
rect 401652 1708 401658 1760
rect 410978 1708 410984 1760
rect 411036 1748 411042 1760
rect 513374 1748 513380 1760
rect 411036 1720 513380 1748
rect 411036 1708 411042 1720
rect 513374 1708 513380 1720
rect 513432 1708 513438 1760
rect 311158 1680 311164 1692
rect 300268 1652 303200 1680
rect 306346 1652 311164 1680
rect 300268 1640 300274 1652
rect 50430 1572 50436 1624
rect 50488 1612 50494 1624
rect 145742 1612 145748 1624
rect 50488 1584 145748 1612
rect 50488 1572 50494 1584
rect 145742 1572 145748 1584
rect 145800 1572 145806 1624
rect 293862 1572 293868 1624
rect 293920 1612 293926 1624
rect 305822 1612 305828 1624
rect 293920 1584 305828 1612
rect 293920 1572 293926 1584
rect 305822 1572 305828 1584
rect 305880 1572 305886 1624
rect 55766 1504 55772 1556
rect 55824 1544 55830 1556
rect 149054 1544 149060 1556
rect 55824 1516 149060 1544
rect 55824 1504 55830 1516
rect 149054 1504 149060 1516
rect 149112 1504 149118 1556
rect 297174 1504 297180 1556
rect 297232 1544 297238 1556
rect 306346 1544 306374 1652
rect 311158 1640 311164 1652
rect 311216 1640 311222 1692
rect 355594 1640 355600 1692
rect 355652 1680 355658 1692
rect 412266 1680 412272 1692
rect 355652 1652 412272 1680
rect 355652 1640 355658 1652
rect 412266 1640 412272 1652
rect 412324 1640 412330 1692
rect 429102 1640 429108 1692
rect 429160 1680 429166 1692
rect 508038 1680 508044 1692
rect 429160 1652 508044 1680
rect 429160 1640 429166 1652
rect 508038 1640 508044 1652
rect 508096 1640 508102 1692
rect 413922 1572 413928 1624
rect 413980 1612 413986 1624
rect 484302 1612 484308 1624
rect 413980 1584 484308 1612
rect 413980 1572 413986 1584
rect 484302 1572 484308 1584
rect 484360 1572 484366 1624
rect 297232 1516 306374 1544
rect 297232 1504 297238 1516
rect 15930 1436 15936 1488
rect 15988 1476 15994 1488
rect 520826 1476 520832 1488
rect 15988 1448 520832 1476
rect 15988 1436 15994 1448
rect 520826 1436 520832 1448
rect 520884 1436 520890 1488
rect 25958 1368 25964 1420
rect 26016 1408 26022 1420
rect 468846 1408 468852 1420
rect 26016 1380 468852 1408
rect 26016 1368 26022 1380
rect 468846 1368 468852 1380
rect 468904 1368 468910 1420
rect 39298 1300 39304 1352
rect 39356 1340 39362 1352
rect 478046 1340 478052 1352
rect 39356 1312 478052 1340
rect 39356 1300 39362 1312
rect 478046 1300 478052 1312
rect 478104 1300 478110 1352
rect 116762 1232 116768 1284
rect 116820 1272 116826 1284
rect 459646 1272 459652 1284
rect 116820 1244 459652 1272
rect 116820 1232 116826 1244
rect 459646 1232 459652 1244
rect 459704 1232 459710 1284
rect 116854 1164 116860 1216
rect 116912 1204 116918 1216
rect 453482 1204 453488 1216
rect 116912 1176 453488 1204
rect 116912 1164 116918 1176
rect 453482 1164 453488 1176
rect 453540 1164 453546 1216
rect 119890 1096 119896 1148
rect 119948 1136 119954 1148
rect 441154 1136 441160 1148
rect 119948 1108 441160 1136
rect 119948 1096 119954 1108
rect 441154 1096 441160 1108
rect 441212 1096 441218 1148
<< via1 >>
rect 38476 158924 38528 158976
rect 145288 158924 145340 158976
rect 34520 158856 34572 158908
rect 142804 158856 142856 158908
rect 30656 158788 30708 158840
rect 140136 158788 140188 158840
rect 26792 158720 26844 158772
rect 137468 158720 137520 158772
rect 11152 158652 11204 158704
rect 127072 158652 127124 158704
rect 22836 158584 22888 158636
rect 134892 158584 134944 158636
rect 70584 158516 70636 158568
rect 167276 158516 167328 158568
rect 66720 158448 66772 158500
rect 164240 158448 164292 158500
rect 62856 158380 62908 158432
rect 161664 158380 161716 158432
rect 55220 158312 55272 158364
rect 156328 158312 156380 158364
rect 18972 158244 19024 158296
rect 132592 158244 132644 158296
rect 104716 158176 104768 158228
rect 189632 158176 189684 158228
rect 90088 158108 90140 158160
rect 179880 158108 179932 158160
rect 58900 158040 58952 158092
rect 158996 158040 159048 158092
rect 51080 157972 51132 158024
rect 153752 157972 153804 158024
rect 47216 157904 47268 157956
rect 151176 157904 151228 157956
rect 43352 157836 43404 157888
rect 148508 157836 148560 157888
rect 148600 157836 148652 157888
rect 218888 157836 218940 157888
rect 15016 157768 15068 157820
rect 129740 157768 129792 157820
rect 132040 157768 132092 157820
rect 207756 157768 207808 157820
rect 144736 157700 144788 157752
rect 216220 157700 216272 157752
rect 129096 157632 129148 157684
rect 205824 157632 205876 157684
rect 117412 157564 117464 157616
rect 198004 157564 198056 157616
rect 108672 157496 108724 157548
rect 192116 157496 192168 157548
rect 100852 157428 100904 157480
rect 186964 157428 187016 157480
rect 119436 157360 119488 157412
rect 510160 157360 510212 157412
rect 84292 157292 84344 157344
rect 82268 157224 82320 157276
rect 77484 157156 77536 157208
rect 171416 157156 171468 157208
rect 174544 157292 174596 157344
rect 181076 157224 181128 157276
rect 173900 157156 173952 157208
rect 190460 157292 190512 157344
rect 201224 157292 201276 157344
rect 253940 157292 253992 157344
rect 426256 157292 426308 157344
rect 458548 157292 458600 157344
rect 472440 157292 472492 157344
rect 527732 157292 527784 157344
rect 191564 157224 191616 157276
rect 193404 157224 193456 157276
rect 248696 157224 248748 157276
rect 428924 157224 428976 157276
rect 462504 157224 462556 157276
rect 473728 157224 473780 157276
rect 529756 157224 529808 157276
rect 189080 157156 189132 157208
rect 189540 157156 189592 157208
rect 246120 157156 246172 157208
rect 442540 157156 442592 157208
rect 482928 157156 482980 157208
rect 484952 157156 485004 157208
rect 540428 157156 540480 157208
rect 76472 157088 76524 157140
rect 170680 157088 170732 157140
rect 173808 157088 173860 157140
rect 69664 157020 69716 157072
rect 166080 157020 166132 157072
rect 169760 157020 169812 157072
rect 177856 157088 177908 157140
rect 238392 157088 238444 157140
rect 251916 157088 251968 157140
rect 287796 157088 287848 157140
rect 434628 157088 434680 157140
rect 471244 157088 471296 157140
rect 474464 157088 474516 157140
rect 530676 157088 530728 157140
rect 236000 157020 236052 157072
rect 244096 157020 244148 157072
rect 282552 157020 282604 157072
rect 436652 157020 436704 157072
rect 474188 157020 474240 157072
rect 476028 157020 476080 157072
rect 533620 157020 533672 157072
rect 68652 156952 68704 157004
rect 165620 156952 165672 157004
rect 168104 156952 168156 157004
rect 231860 156952 231912 157004
rect 240232 156952 240284 157004
rect 280252 156952 280304 157004
rect 437388 156952 437440 157004
rect 475108 156952 475160 157004
rect 476948 156952 477000 157004
rect 534632 156952 534684 157004
rect 54024 156884 54076 156936
rect 155960 156884 156012 156936
rect 166172 156884 166224 156936
rect 230572 156884 230624 156936
rect 236276 156884 236328 156936
rect 277584 156884 277636 156936
rect 439964 156884 440016 156936
rect 479064 156884 479116 156936
rect 480076 156884 480128 156936
rect 539508 156884 539560 156936
rect 46204 156816 46256 156868
rect 150624 156816 150676 156868
rect 158352 156816 158404 156868
rect 225328 156816 225380 156868
rect 233424 156816 233476 156868
rect 275376 156816 275428 156868
rect 441528 156816 441580 156868
rect 481916 156816 481968 156868
rect 484216 156816 484268 156868
rect 545304 156816 545356 156868
rect 33600 156748 33652 156800
rect 142252 156748 142304 156800
rect 146668 156748 146720 156800
rect 228548 156748 228600 156800
rect 272156 156748 272208 156800
rect 442816 156748 442868 156800
rect 483940 156748 483992 156800
rect 486700 156748 486752 156800
rect 549168 156748 549220 156800
rect 17960 156680 18012 156732
rect 131672 156680 131724 156732
rect 134984 156680 135036 156732
rect 212908 156680 212960 156732
rect 261760 156680 261812 156732
rect 447048 156680 447100 156732
rect 489736 156680 489788 156732
rect 490656 156680 490708 156732
rect 555056 156680 555108 156732
rect 6276 156612 6328 156664
rect 123852 156612 123904 156664
rect 131028 156612 131080 156664
rect 207020 156612 207072 156664
rect 207112 156612 207164 156664
rect 258080 156612 258132 156664
rect 263600 156612 263652 156664
rect 295524 156612 295576 156664
rect 415860 156612 415912 156664
rect 443000 156612 443052 156664
rect 448428 156612 448480 156664
rect 491668 156612 491720 156664
rect 491944 156612 491996 156664
rect 556988 156612 557040 156664
rect 92020 156544 92072 156596
rect 175740 156544 175792 156596
rect 225972 156544 226024 156596
rect 420736 156544 420788 156596
rect 450728 156544 450780 156596
rect 469864 156544 469916 156596
rect 523868 156544 523920 156596
rect 99840 156476 99892 156528
rect 186412 156476 186464 156528
rect 196716 156476 196768 156528
rect 197360 156476 197412 156528
rect 205088 156476 205140 156528
rect 256700 156476 256752 156528
rect 467196 156476 467248 156528
rect 520004 156476 520056 156528
rect 103796 156408 103848 156460
rect 182088 156408 182140 156460
rect 105728 156340 105780 156392
rect 186320 156408 186372 156460
rect 199384 156340 199436 156392
rect 209872 156408 209924 156460
rect 217508 156408 217560 156460
rect 254584 156408 254636 156460
rect 462688 156408 462740 156460
rect 513104 156408 513156 156460
rect 239036 156340 239088 156392
rect 456524 156340 456576 156392
rect 504364 156340 504416 156392
rect 107660 156272 107712 156324
rect 228548 156272 228600 156324
rect 452568 156272 452620 156324
rect 498568 156272 498620 156324
rect 115480 156204 115532 156256
rect 233792 156204 233844 156256
rect 449072 156204 449124 156256
rect 492680 156204 492732 156256
rect 119344 156136 119396 156188
rect 194968 156136 195020 156188
rect 112536 156068 112588 156120
rect 128084 156068 128136 156120
rect 204812 156068 204864 156120
rect 247224 156136 247276 156188
rect 453580 156136 453632 156188
rect 499488 156136 499540 156188
rect 241612 156068 241664 156120
rect 450360 156068 450412 156120
rect 494612 156068 494664 156120
rect 96896 156000 96948 156052
rect 155868 156000 155920 156052
rect 158720 156000 158772 156052
rect 14096 155864 14148 155916
rect 129004 155932 129056 155984
rect 44272 155864 44324 155916
rect 140688 155864 140740 155916
rect 140780 155864 140832 155916
rect 149612 155864 149664 155916
rect 155408 155932 155460 155984
rect 156604 155932 156656 155984
rect 218152 156000 218204 156052
rect 220636 156000 220688 156052
rect 259828 156000 259880 156052
rect 286968 156043 287020 156052
rect 286968 156009 286977 156043
rect 286977 156009 287011 156043
rect 287011 156009 287020 156043
rect 286968 156000 287020 156009
rect 445116 156000 445168 156052
rect 486792 156000 486844 156052
rect 220820 155932 220872 155984
rect 222108 155932 222160 155984
rect 265072 155932 265124 155984
rect 158904 155864 158956 155916
rect 163228 155864 163280 155916
rect 179420 155864 179472 155916
rect 180800 155864 180852 155916
rect 186596 155864 186648 155916
rect 190552 155864 190604 155916
rect 197360 155864 197412 155916
rect 201960 155864 202012 155916
rect 5264 155796 5316 155848
rect 102140 155796 102192 155848
rect 110604 155796 110656 155848
rect 113180 155796 113232 155848
rect 118332 155796 118384 155848
rect 200028 155796 200080 155848
rect 200212 155796 200264 155848
rect 202788 155796 202840 155848
rect 242164 155864 242216 155916
rect 208492 155796 208544 155848
rect 255412 155864 255464 155916
rect 257804 155864 257856 155916
rect 252928 155796 252980 155848
rect 287060 155932 287112 155984
rect 286968 155864 287020 155916
rect 289912 155864 289964 155916
rect 309140 155864 309192 155916
rect 309416 155864 309468 155916
rect 315304 155864 315356 155916
rect 329748 155864 329800 155916
rect 329932 155864 329984 155916
rect 336464 155864 336516 155916
rect 338672 155864 338724 155916
rect 344192 155864 344244 155916
rect 354220 155864 354272 155916
rect 355968 155864 356020 155916
rect 388168 155864 388220 155916
rect 393228 155864 393280 155916
rect 401692 155864 401744 155916
rect 403992 155864 404044 155916
rect 404820 155864 404872 155916
rect 407856 155864 407908 155916
rect 287980 155796 288032 155848
rect 293040 155796 293092 155848
rect 294788 155796 294840 155848
rect 55956 155728 56008 155780
rect 153476 155728 153528 155780
rect 159272 155728 159324 155780
rect 169760 155728 169812 155780
rect 173808 155728 173860 155780
rect 175924 155728 175976 155780
rect 40408 155660 40460 155712
rect 137192 155660 137244 155712
rect 172980 155660 173032 155712
rect 235080 155728 235132 155780
rect 229376 155660 229428 155712
rect 237012 155660 237064 155712
rect 237288 155660 237340 155712
rect 246028 155728 246080 155780
rect 280712 155728 280764 155780
rect 281172 155728 281224 155780
rect 286692 155728 286744 155780
rect 246948 155660 247000 155712
rect 247040 155660 247092 155712
rect 31668 155592 31720 155644
rect 156512 155592 156564 155644
rect 160284 155592 160336 155644
rect 224040 155592 224092 155644
rect 249064 155592 249116 155644
rect 250904 155592 250956 155644
rect 277400 155592 277452 155644
rect 282092 155660 282144 155712
rect 300676 155728 300728 155780
rect 316040 155796 316092 155848
rect 320180 155796 320232 155848
rect 307300 155728 307352 155780
rect 309232 155728 309284 155780
rect 312360 155728 312412 155780
rect 326804 155728 326856 155780
rect 328920 155796 328972 155848
rect 334440 155796 334492 155848
rect 334808 155796 334860 155848
rect 340788 155796 340840 155848
rect 353300 155796 353352 155848
rect 355416 155796 355468 155848
rect 365076 155796 365128 155848
rect 365996 155796 366048 155848
rect 403440 155796 403492 155848
rect 406936 155796 406988 155848
rect 412548 155864 412600 155916
rect 412640 155864 412692 155916
rect 506940 155932 506992 155984
rect 428372 155864 428424 155916
rect 430212 155864 430264 155916
rect 464436 155864 464488 155916
rect 464988 155864 465040 155916
rect 517060 155864 517112 155916
rect 574560 155864 574612 155916
rect 425428 155796 425480 155848
rect 427636 155796 427688 155848
rect 460480 155796 460532 155848
rect 467748 155796 467800 155848
rect 520924 155796 520976 155848
rect 333244 155728 333296 155780
rect 380900 155728 380952 155780
rect 384488 155728 384540 155780
rect 414664 155728 414716 155780
rect 429292 155728 429344 155780
rect 430488 155728 430540 155780
rect 465356 155728 465408 155780
rect 473084 155728 473136 155780
rect 528744 155728 528796 155780
rect 313740 155660 313792 155712
rect 314292 155660 314344 155712
rect 328184 155660 328236 155712
rect 333796 155660 333848 155712
rect 339408 155660 339460 155712
rect 342536 155660 342588 155712
rect 348240 155660 348292 155712
rect 404176 155660 404228 155712
rect 409696 155660 409748 155712
rect 434168 155660 434220 155712
rect 435364 155660 435416 155712
rect 472164 155660 472216 155712
rect 478328 155660 478380 155712
rect 536564 155660 536616 155712
rect 280160 155592 280212 155644
rect 291752 155592 291804 155644
rect 291844 155592 291896 155644
rect 304540 155592 304592 155644
rect 311992 155592 312044 155644
rect 35532 155524 35584 155576
rect 140780 155524 140832 155576
rect 141792 155524 141844 155576
rect 143816 155524 143868 155576
rect 153108 155524 153160 155576
rect 155316 155524 155368 155576
rect 162768 155524 162820 155576
rect 164148 155524 164200 155576
rect 225604 155524 225656 155576
rect 229376 155524 229428 155576
rect 229468 155524 229520 155576
rect 264980 155524 265032 155576
rect 266544 155524 266596 155576
rect 288992 155524 289044 155576
rect 293868 155524 293920 155576
rect 29644 155456 29696 155508
rect 31668 155456 31720 155508
rect 32588 155456 32640 155508
rect 132776 155456 132828 155508
rect 12164 155388 12216 155440
rect 25504 155388 25556 155440
rect 27712 155388 27764 155440
rect 133972 155456 134024 155508
rect 139860 155456 139912 155508
rect 132960 155388 133012 155440
rect 23848 155320 23900 155372
rect 9220 155252 9272 155304
rect 125232 155320 125284 155372
rect 130108 155320 130160 155372
rect 4344 155184 4396 155236
rect 11520 155184 11572 155236
rect 16028 155184 16080 155236
rect 132960 155252 133012 155304
rect 136548 155320 136600 155372
rect 143632 155388 143684 155440
rect 135168 155252 135220 155304
rect 52092 155116 52144 155168
rect 144828 155320 144880 155372
rect 145656 155456 145708 155508
rect 147588 155456 147640 155508
rect 156604 155456 156656 155508
rect 156696 155456 156748 155508
rect 221740 155456 221792 155508
rect 281540 155456 281592 155508
rect 284024 155456 284076 155508
rect 284116 155456 284168 155508
rect 306932 155524 306984 155576
rect 313096 155524 313148 155576
rect 308036 155456 308088 155508
rect 206468 155388 206520 155440
rect 211896 155388 211948 155440
rect 211988 155388 212040 155440
rect 146484 155320 146536 155372
rect 149060 155320 149112 155372
rect 151544 155320 151596 155372
rect 158720 155320 158772 155372
rect 217784 155388 217836 155440
rect 222108 155388 222160 155440
rect 226524 155388 226576 155440
rect 226616 155388 226668 155440
rect 269396 155388 269448 155440
rect 269488 155388 269540 155440
rect 229284 155320 229336 155372
rect 258724 155320 258776 155372
rect 260564 155320 260616 155372
rect 260656 155320 260708 155372
rect 265532 155320 265584 155372
rect 272800 155320 272852 155372
rect 277124 155320 277176 155372
rect 277492 155388 277544 155440
rect 279148 155388 279200 155440
rect 279240 155388 279292 155440
rect 298744 155388 298796 155440
rect 290004 155320 290056 155372
rect 290924 155320 290976 155372
rect 308588 155388 308640 155440
rect 310428 155456 310480 155508
rect 321652 155592 321704 155644
rect 322112 155592 322164 155644
rect 334624 155592 334676 155644
rect 337660 155592 337712 155644
rect 342720 155592 342772 155644
rect 344560 155592 344612 155644
rect 349528 155592 349580 155644
rect 385868 155592 385920 155644
rect 389364 155592 389416 155644
rect 406108 155592 406160 155644
rect 319168 155524 319220 155576
rect 332600 155524 332652 155576
rect 335728 155524 335780 155576
rect 340972 155524 341024 155576
rect 358176 155524 358228 155576
rect 358820 155524 358872 155576
rect 379612 155524 379664 155576
rect 382556 155524 382608 155576
rect 385960 155524 386012 155576
rect 390284 155524 390336 155576
rect 411996 155524 412048 155576
rect 437112 155592 437164 155644
rect 438676 155592 438728 155644
rect 477040 155592 477092 155644
rect 479616 155592 479668 155644
rect 538496 155592 538548 155644
rect 413836 155524 413888 155576
rect 416688 155524 416740 155576
rect 430304 155524 430356 155576
rect 433064 155524 433116 155576
rect 469312 155524 469364 155576
rect 482192 155524 482244 155576
rect 542360 155524 542412 155576
rect 575480 155524 575532 155576
rect 576492 155524 576544 155576
rect 578424 155524 578476 155576
rect 313280 155456 313332 155508
rect 328368 155456 328420 155508
rect 330852 155456 330904 155508
rect 336556 155456 336608 155508
rect 378140 155456 378192 155508
rect 380624 155456 380676 155508
rect 382372 155456 382424 155508
rect 385500 155456 385552 155508
rect 386788 155456 386840 155508
rect 391296 155456 391348 155508
rect 404268 155456 404320 155508
rect 405924 155456 405976 155508
rect 407764 155456 407816 155508
rect 412456 155456 412508 155508
rect 438124 155456 438176 155508
rect 311164 155388 311216 155440
rect 311348 155388 311400 155440
rect 326712 155388 326764 155440
rect 327908 155388 327960 155440
rect 338488 155388 338540 155440
rect 398564 155388 398616 155440
rect 318984 155320 319036 155372
rect 321100 155320 321152 155372
rect 334164 155320 334216 155372
rect 382280 155320 382332 155372
rect 386420 155320 386472 155372
rect 401600 155320 401652 155372
rect 404912 155320 404964 155372
rect 411168 155388 411220 155440
rect 436100 155388 436152 155440
rect 438032 155388 438084 155440
rect 476120 155456 476172 155508
rect 484768 155456 484820 155508
rect 546316 155456 546368 155508
rect 441252 155388 441304 155440
rect 480996 155388 481048 155440
rect 483572 155388 483624 155440
rect 544292 155388 544344 155440
rect 417608 155320 417660 155372
rect 417976 155320 418028 155372
rect 444932 155320 444984 155372
rect 445668 155320 445720 155372
rect 484860 155320 484912 155372
rect 488356 155320 488408 155372
rect 552112 155320 552164 155372
rect 203156 155252 203208 155304
rect 220636 155252 220688 155304
rect 223672 155252 223724 155304
rect 269028 155252 269080 155304
rect 270408 155252 270460 155304
rect 202236 155184 202288 155236
rect 209044 155184 209096 155236
rect 210976 155184 211028 155236
rect 185584 155116 185636 155168
rect 240232 155116 240284 155168
rect 39396 155048 39448 155100
rect 124128 155048 124180 155100
rect 202880 155048 202932 155100
rect 209964 155048 210016 155100
rect 243452 155048 243504 155100
rect 244832 155048 244884 155100
rect 252652 155184 252704 155236
rect 253848 155184 253900 155236
rect 275284 155252 275336 155304
rect 300124 155252 300176 155304
rect 301596 155252 301648 155304
rect 308496 155252 308548 155304
rect 324412 155252 324464 155304
rect 331864 155252 331916 155304
rect 337936 155252 337988 155304
rect 402244 155252 402296 155304
rect 422484 155252 422536 155304
rect 424968 155252 425020 155304
rect 456616 155252 456668 155304
rect 456708 155252 456760 155304
rect 502432 155252 502484 155304
rect 502984 155252 503036 155304
rect 569684 155252 569736 155304
rect 296904 155184 296956 155236
rect 304908 155184 304960 155236
rect 305552 155184 305604 155236
rect 322848 155184 322900 155236
rect 323032 155184 323084 155236
rect 334072 155184 334124 155236
rect 343548 155184 343600 155236
rect 349068 155184 349120 155236
rect 384856 155184 384908 155236
rect 388352 155184 388404 155236
rect 401508 155184 401560 155236
rect 421564 155184 421616 155236
rect 422024 155184 422076 155236
rect 452752 155184 452804 155236
rect 454868 155184 454920 155236
rect 501420 155184 501472 155236
rect 502248 155184 502300 155236
rect 572628 155184 572680 155236
rect 249984 155116 250036 155168
rect 281448 155116 281500 155168
rect 297916 155116 297968 155168
rect 316408 155116 316460 155168
rect 259368 155048 259420 155100
rect 285036 155048 285088 155100
rect 302240 155048 302292 155100
rect 314660 155048 314712 155100
rect 320088 155116 320140 155168
rect 324044 155116 324096 155168
rect 333980 155116 334032 155168
rect 355232 155116 355284 155168
rect 356704 155116 356756 155168
rect 405924 155116 405976 155168
rect 409788 155116 409840 155168
rect 426348 155116 426400 155168
rect 428280 155116 428332 155168
rect 86224 154980 86276 155032
rect 74540 154912 74592 154964
rect 167000 154980 167052 155032
rect 167092 154980 167144 155032
rect 171232 154980 171284 155032
rect 182088 154980 182140 155032
rect 187608 154980 187660 155032
rect 242256 154980 242308 155032
rect 480 154844 532 154896
rect 1308 154844 1360 154896
rect 97908 154844 97960 154896
rect 169760 154844 169812 154896
rect 175832 154844 175884 154896
rect 176844 154844 176896 154896
rect 177948 154844 178000 154896
rect 194232 154844 194284 154896
rect 94964 154776 95016 154828
rect 193128 154776 193180 154828
rect 194416 154844 194468 154896
rect 241152 154844 241204 154896
rect 195520 154776 195572 154828
rect 78404 154708 78456 154760
rect 110420 154708 110472 154760
rect 113548 154708 113600 154760
rect 56968 154640 57020 154692
rect 116768 154640 116820 154692
rect 120724 154708 120776 154760
rect 178040 154708 178092 154760
rect 178776 154708 178828 154760
rect 186320 154708 186372 154760
rect 121276 154640 121328 154692
rect 182088 154640 182140 154692
rect 182732 154640 182784 154692
rect 194968 154708 195020 154760
rect 195336 154708 195388 154760
rect 245108 154912 245160 154964
rect 277492 154980 277544 155032
rect 285680 154980 285732 155032
rect 268476 154912 268528 154964
rect 276296 154912 276348 154964
rect 297732 154980 297784 155032
rect 302608 154912 302660 154964
rect 307484 154980 307536 155032
rect 317236 155048 317288 155100
rect 326896 155048 326948 155100
rect 326988 155048 327040 155100
rect 338028 155048 338080 155100
rect 356244 155048 356296 155100
rect 357440 155048 357492 155100
rect 400312 155048 400364 155100
rect 402060 155048 402112 155100
rect 321560 154980 321612 155032
rect 325056 154980 325108 155032
rect 336648 154980 336700 155032
rect 399576 154980 399628 155032
rect 418620 155048 418672 155100
rect 413744 154980 413796 155032
rect 424416 155048 424468 155100
rect 425612 155048 425664 155100
rect 457628 155048 457680 155100
rect 255320 154844 255372 154896
rect 199292 154708 199344 154760
rect 246948 154776 247000 154828
rect 247040 154776 247092 154828
rect 247408 154776 247460 154828
rect 248972 154776 249024 154828
rect 254860 154776 254912 154828
rect 262864 154844 262916 154896
rect 270408 154844 270460 154896
rect 291108 154844 291160 154896
rect 292856 154844 292908 154896
rect 306288 154844 306340 154896
rect 319628 154912 319680 154964
rect 325976 154912 326028 154964
rect 337200 154912 337252 154964
rect 345480 154912 345532 154964
rect 347596 154912 347648 154964
rect 357164 154912 357216 154964
rect 357992 154912 358044 154964
rect 384212 154912 384264 154964
rect 387432 154912 387484 154964
rect 400220 154912 400272 154964
rect 402980 154912 403032 154964
rect 404728 154912 404780 154964
rect 413652 154912 413704 154964
rect 419448 154980 419500 155032
rect 448796 154980 448848 155032
rect 464620 155116 464672 155168
rect 516048 155116 516100 155168
rect 463332 155048 463384 155100
rect 514116 155048 514168 155100
rect 461492 154980 461544 155032
rect 462044 154980 462096 155032
rect 512184 154980 512236 155032
rect 415216 154912 415268 154964
rect 423036 154912 423088 154964
rect 453672 154912 453724 154964
rect 460112 154912 460164 154964
rect 509240 154912 509292 154964
rect 561680 154912 561732 154964
rect 563796 154912 563848 154964
rect 316592 154844 316644 154896
rect 191472 154640 191524 154692
rect 198280 154640 198332 154692
rect 89168 154572 89220 154624
rect 120172 154572 120224 154624
rect 122288 154572 122340 154624
rect 75460 154504 75512 154556
rect 167000 154504 167052 154556
rect 183008 154504 183060 154556
rect 183652 154572 183704 154624
rect 196348 154572 196400 154624
rect 206100 154640 206152 154692
rect 213920 154572 213972 154624
rect 219256 154572 219308 154624
rect 219624 154640 219676 154692
rect 252560 154640 252612 154692
rect 273260 154776 273312 154828
rect 273352 154776 273404 154828
rect 262864 154708 262916 154760
rect 256792 154640 256844 154692
rect 222108 154572 222160 154624
rect 222660 154572 222712 154624
rect 263600 154640 263652 154692
rect 264612 154708 264664 154760
rect 279332 154708 279384 154760
rect 275928 154572 275980 154624
rect 201500 154504 201552 154556
rect 202788 154504 202840 154556
rect 71596 154436 71648 154488
rect 59912 154368 59964 154420
rect 159640 154368 159692 154420
rect 64788 154300 64840 154352
rect 162860 154300 162912 154352
rect 164056 154436 164108 154488
rect 172612 154436 172664 154488
rect 175924 154436 175976 154488
rect 192760 154436 192812 154488
rect 192852 154436 192904 154488
rect 248052 154436 248104 154488
rect 249984 154436 250036 154488
rect 252560 154504 252612 154556
rect 262404 154504 262456 154556
rect 264980 154504 265032 154556
rect 272800 154504 272852 154556
rect 277216 154640 277268 154692
rect 283104 154776 283156 154828
rect 286048 154776 286100 154828
rect 298008 154708 298060 154760
rect 306564 154776 306616 154828
rect 317328 154776 317380 154828
rect 321744 154776 321796 154828
rect 303620 154708 303672 154760
rect 322204 154708 322256 154760
rect 332784 154844 332836 154896
rect 338672 154844 338724 154896
rect 400956 154844 401008 154896
rect 420552 154844 420604 154896
rect 341616 154776 341668 154828
rect 347504 154776 347556 154828
rect 395988 154776 396040 154828
rect 407028 154776 407080 154828
rect 420460 154776 420512 154828
rect 449808 154844 449860 154896
rect 459468 154844 459520 154896
rect 508228 154844 508280 154896
rect 289728 154640 289780 154692
rect 299572 154640 299624 154692
rect 299664 154640 299716 154692
rect 282368 154572 282420 154624
rect 285864 154572 285916 154624
rect 288440 154504 288492 154556
rect 291568 154504 291620 154556
rect 293960 154504 294012 154556
rect 305920 154572 305972 154624
rect 306472 154572 306524 154624
rect 309876 154504 309928 154556
rect 253296 154436 253348 154488
rect 255320 154436 255372 154488
rect 267832 154436 267884 154488
rect 271788 154436 271840 154488
rect 273352 154436 273404 154488
rect 279332 154436 279384 154488
rect 293592 154436 293644 154488
rect 304632 154436 304684 154488
rect 318156 154640 318208 154692
rect 324320 154504 324372 154556
rect 320916 154436 320968 154488
rect 340604 154708 340656 154760
rect 339684 154640 339736 154692
rect 346308 154640 346360 154692
rect 336740 154572 336792 154624
rect 330668 154504 330720 154556
rect 344376 154504 344428 154556
rect 406752 154708 406804 154760
rect 417792 154708 417844 154760
rect 445852 154776 445904 154828
rect 460664 154776 460716 154828
rect 510252 154776 510304 154828
rect 441988 154708 442040 154760
rect 457536 154708 457588 154760
rect 505376 154708 505428 154760
rect 352288 154640 352340 154692
rect 353392 154640 353444 154692
rect 409420 154640 409472 154692
rect 433248 154640 433300 154692
rect 468300 154640 468352 154692
rect 346492 154572 346544 154624
rect 347044 154504 347096 154556
rect 331956 154436 332008 154488
rect 340972 154436 341024 154488
rect 343732 154436 343784 154488
rect 184296 154368 184348 154420
rect 184664 154368 184716 154420
rect 167460 154300 167512 154352
rect 169760 154300 169812 154352
rect 184940 154300 184992 154352
rect 188528 154368 188580 154420
rect 245660 154368 245712 154420
rect 249064 154368 249116 154420
rect 261116 154368 261168 154420
rect 262680 154368 262732 154420
rect 294880 154368 294932 154420
rect 303620 154368 303672 154420
rect 242900 154300 242952 154352
rect 243176 154300 243228 154352
rect 281908 154300 281960 154352
rect 291108 154300 291160 154352
rect 303988 154300 304040 154352
rect 53104 154232 53156 154284
rect 155040 154232 155092 154284
rect 155868 154232 155920 154284
rect 162768 154232 162820 154284
rect 177212 154232 177264 154284
rect 177948 154232 178000 154284
rect 237656 154232 237708 154284
rect 239220 154232 239272 154284
rect 279332 154232 279384 154284
rect 284484 154232 284536 154284
rect 285680 154232 285732 154284
rect 301412 154232 301464 154284
rect 306288 154232 306340 154284
rect 315028 154232 315080 154284
rect 348424 154572 348476 154624
rect 349344 154572 349396 154624
rect 350356 154572 350408 154624
rect 351368 154572 351420 154624
rect 354128 154504 354180 154556
rect 361488 154504 361540 154556
rect 362040 154504 362092 154556
rect 362592 154504 362644 154556
rect 363052 154504 363104 154556
rect 365628 154504 365680 154556
rect 367928 154572 367980 154624
rect 366456 154504 366508 154556
rect 368848 154572 368900 154624
rect 353484 154436 353536 154488
rect 362868 154436 362920 154488
rect 363972 154436 364024 154488
rect 367008 154436 367060 154488
rect 369860 154436 369912 154488
rect 352840 154368 352892 154420
rect 367744 154368 367796 154420
rect 370872 154572 370924 154624
rect 374920 154504 374972 154556
rect 381544 154572 381596 154624
rect 375196 154436 375248 154488
rect 379612 154436 379664 154488
rect 376208 154368 376260 154420
rect 383476 154572 383528 154624
rect 387708 154504 387760 154556
rect 401048 154572 401100 154624
rect 414572 154572 414624 154624
rect 440976 154572 441028 154624
rect 511172 154640 511224 154692
rect 410708 154504 410760 154556
rect 435180 154504 435232 154556
rect 461400 154504 461452 154556
rect 500132 154572 500184 154624
rect 503352 154572 503404 154624
rect 471796 154504 471848 154556
rect 526812 154504 526864 154556
rect 390468 154436 390520 154488
rect 401600 154436 401652 154488
rect 408316 154436 408368 154488
rect 432236 154436 432288 154488
rect 432604 154436 432656 154488
rect 480904 154436 480956 154488
rect 484952 154436 485004 154488
rect 487068 154436 487120 154488
rect 550180 154436 550232 154488
rect 383292 154368 383344 154420
rect 394240 154368 394292 154420
rect 395068 154368 395120 154420
rect 352104 154300 352156 154352
rect 368388 154300 368440 154352
rect 371792 154300 371844 154352
rect 384028 154300 384080 154352
rect 395160 154300 395212 154352
rect 410800 154368 410852 154420
rect 413928 154368 413980 154420
rect 440056 154368 440108 154420
rect 491208 154368 491260 154420
rect 556068 154368 556120 154420
rect 411812 154300 411864 154352
rect 413284 154300 413336 154352
rect 439044 154300 439096 154352
rect 493968 154300 494020 154352
rect 559932 154300 559984 154352
rect 350816 154232 350868 154284
rect 369676 154232 369728 154284
rect 373724 154232 373776 154284
rect 381452 154232 381504 154284
rect 386788 154232 386840 154284
rect 393044 154232 393096 154284
rect 408868 154232 408920 154284
rect 494612 154232 494664 154284
rect 560944 154232 560996 154284
rect 48228 154164 48280 154216
rect 36544 154096 36596 154148
rect 24768 154028 24820 154080
rect 136180 154028 136232 154080
rect 20904 153960 20956 154012
rect 133880 153960 133932 154012
rect 135168 153960 135220 154012
rect 136548 153960 136600 154012
rect 137836 154096 137888 154148
rect 140872 154096 140924 154148
rect 144828 154096 144880 154148
rect 140964 154028 141016 154080
rect 156512 154164 156564 154216
rect 170036 154164 170088 154216
rect 152004 154096 152056 154148
rect 160100 154096 160152 154148
rect 164792 154096 164844 154148
rect 165160 154096 165212 154148
rect 169024 154096 169076 154148
rect 232504 154164 232556 154216
rect 235356 154164 235408 154216
rect 276664 154164 276716 154216
rect 298836 154164 298888 154216
rect 302240 154164 302292 154216
rect 312452 154164 312504 154216
rect 347596 154164 347648 154216
rect 350172 154164 350224 154216
rect 372988 154164 373040 154216
rect 378600 154164 378652 154216
rect 382096 154164 382148 154216
rect 392308 154164 392360 154216
rect 394424 154164 394476 154216
rect 395712 154164 395764 154216
rect 412548 154164 412600 154216
rect 419172 154164 419224 154216
rect 447876 154164 447928 154216
rect 496544 154164 496596 154216
rect 561680 154164 561732 154216
rect 229836 154096 229888 154148
rect 231492 154096 231544 154148
rect 154580 154028 154632 154080
rect 155316 154028 155368 154080
rect 156972 154028 157024 154080
rect 157340 154028 157392 154080
rect 224960 154028 225012 154080
rect 227536 154028 227588 154080
rect 271512 154028 271564 154080
rect 273260 154096 273312 154148
rect 285772 154096 285824 154148
rect 291752 154096 291804 154148
rect 306656 154096 306708 154148
rect 372344 154096 372396 154148
rect 377680 154096 377732 154148
rect 384948 154096 385000 154148
rect 397184 154096 397236 154148
rect 397276 154096 397328 154148
rect 415676 154096 415728 154148
rect 421748 154096 421800 154148
rect 451740 154096 451792 154148
rect 497832 154096 497884 154148
rect 565728 154096 565780 154148
rect 274088 154028 274140 154080
rect 281448 154028 281500 154080
rect 296168 154028 296220 154080
rect 304908 154028 304960 154080
rect 317696 154028 317748 154080
rect 386236 154028 386288 154080
rect 398748 154028 398800 154080
rect 400128 154028 400180 154080
rect 419540 154028 419592 154080
rect 426900 154028 426952 154080
rect 459560 154028 459612 154080
rect 499120 154028 499172 154080
rect 567752 154028 567804 154080
rect 17040 153892 17092 153944
rect 131120 153892 131172 153944
rect 131304 153892 131356 153944
rect 144000 153960 144052 154012
rect 149244 153960 149296 154012
rect 216864 153960 216916 154012
rect 219716 153960 219768 154012
rect 266360 153960 266412 154012
rect 276020 153960 276072 154012
rect 291200 153960 291252 154012
rect 293040 153960 293092 154012
rect 311900 153960 311952 154012
rect 311992 153960 312044 154012
rect 322940 153960 322992 154012
rect 347780 153960 347832 154012
rect 351460 153960 351512 154012
rect 373908 153960 373960 154012
rect 378140 153960 378192 154012
rect 389824 153960 389876 154012
rect 401692 153960 401744 154012
rect 405464 153960 405516 154012
rect 427360 153960 427412 154012
rect 429568 153960 429620 154012
rect 463424 153960 463476 154012
rect 500868 153960 500920 154012
rect 570696 153960 570748 154012
rect 1400 153824 1452 153876
rect 120632 153824 120684 153876
rect 120724 153824 120776 153876
rect 125784 153824 125836 153876
rect 130384 153824 130436 153876
rect 131212 153824 131264 153876
rect 132960 153824 133012 153876
rect 133052 153824 133104 153876
rect 135536 153824 135588 153876
rect 138112 153892 138164 153944
rect 138204 153892 138256 153944
rect 140688 153892 140740 153944
rect 140780 153892 140832 153944
rect 143540 153892 143592 153944
rect 143632 153892 143684 153944
rect 146576 153892 146628 153944
rect 211620 153892 211672 153944
rect 215852 153892 215904 153944
rect 203892 153824 203944 153876
rect 204168 153824 204220 153876
rect 255872 153824 255924 153876
rect 263600 153892 263652 153944
rect 270500 153892 270552 153944
rect 278228 153892 278280 153944
rect 305276 153892 305328 153944
rect 309140 153892 309192 153944
rect 320272 153892 320324 153944
rect 334440 153892 334492 153944
rect 339132 153892 339184 153944
rect 376484 153892 376536 153944
rect 380900 153892 380952 153944
rect 382740 153892 382792 153944
rect 388168 153892 388220 153944
rect 391204 153892 391256 153944
rect 404268 153892 404320 153944
rect 408040 153892 408092 153944
rect 431224 153892 431276 153944
rect 431776 153892 431828 153944
rect 467288 153892 467340 153944
rect 503076 153892 503128 153944
rect 573548 153892 573600 153944
rect 263692 153824 263744 153876
rect 83280 153756 83332 153808
rect 175280 153756 175332 153808
rect 179420 153756 179472 153808
rect 211160 153756 211212 153808
rect 260564 153756 260616 153808
rect 292580 153824 292632 153876
rect 295800 153824 295852 153876
rect 317052 153824 317104 153876
rect 336464 153824 336516 153876
rect 339776 153824 339828 153876
rect 340788 153824 340840 153876
rect 342996 153824 343048 153876
rect 373632 153824 373684 153876
rect 379428 153824 379480 153876
rect 389088 153824 389140 153876
rect 400220 153824 400272 153876
rect 402704 153824 402756 153876
rect 423496 153824 423548 153876
rect 456248 153824 456300 153876
rect 500132 153824 500184 153876
rect 501696 153824 501748 153876
rect 571616 153824 571668 153876
rect 270408 153756 270460 153808
rect 280620 153756 280672 153808
rect 287060 153756 287112 153808
rect 289084 153756 289136 153808
rect 290004 153756 290056 153808
rect 291660 153756 291712 153808
rect 326804 153756 326856 153808
rect 328092 153756 328144 153808
rect 328184 153756 328236 153808
rect 329380 153756 329432 153808
rect 339408 153756 339460 153808
rect 342352 153756 342404 153808
rect 377496 153756 377548 153808
rect 382372 153756 382424 153808
rect 385776 153756 385828 153808
rect 398104 153756 398156 153808
rect 398288 153756 398340 153808
rect 413836 153756 413888 153808
rect 416504 153756 416556 153808
rect 443920 153756 443972 153808
rect 470324 153756 470376 153808
rect 524880 153756 524932 153808
rect 93032 153688 93084 153740
rect 91100 153620 91152 153672
rect 180432 153688 180484 153740
rect 185584 153688 185636 153740
rect 213920 153688 213972 153740
rect 262220 153688 262272 153740
rect 265624 153688 265676 153740
rect 273352 153688 273404 153740
rect 283196 153688 283248 153740
rect 327080 153688 327132 153740
rect 331312 153688 331364 153740
rect 378784 153688 378836 153740
rect 384212 153688 384264 153740
rect 391848 153688 391900 153740
rect 403440 153688 403492 153740
rect 424324 153688 424376 153740
rect 455604 153688 455656 153740
rect 469128 153688 469180 153740
rect 522856 153688 522908 153740
rect 178040 153620 178092 153672
rect 195428 153620 195480 153672
rect 195520 153620 195572 153672
rect 219624 153620 219676 153672
rect 260932 153620 260984 153672
rect 263048 153620 263100 153672
rect 269396 153620 269448 153672
rect 270868 153620 270920 153672
rect 321744 153620 321796 153672
rect 326712 153620 326764 153672
rect 327448 153620 327500 153672
rect 336556 153620 336608 153672
rect 340420 153620 340472 153672
rect 370964 153620 371016 153672
rect 375748 153620 375800 153672
rect 380072 153620 380124 153672
rect 385868 153620 385920 153672
rect 388536 153620 388588 153672
rect 400312 153620 400364 153672
rect 403532 153620 403584 153672
rect 413652 153620 413704 153672
rect 466184 153620 466236 153672
rect 518992 153620 519044 153672
rect 98920 153552 98972 153604
rect 185676 153552 185728 153604
rect 193128 153552 193180 153604
rect 208400 153552 208452 153604
rect 208492 153552 208544 153604
rect 214288 153552 214340 153604
rect 321652 153552 321704 153604
rect 327080 153552 327132 153604
rect 337936 153552 337988 153604
rect 341064 153552 341116 153604
rect 369032 153552 369084 153604
rect 372804 153552 372856 153604
rect 378048 153552 378100 153604
rect 382280 153552 382332 153604
rect 393780 153552 393832 153604
rect 405924 153552 405976 153604
rect 417148 153552 417200 153604
rect 417976 153552 418028 153604
rect 443828 153552 443880 153604
rect 445668 153552 445720 153604
rect 455236 153552 455288 153604
rect 456708 153552 456760 153604
rect 463608 153552 463660 153604
rect 515128 153552 515180 153604
rect 1308 153484 1360 153536
rect 120080 153484 120132 153536
rect 193404 153484 193456 153536
rect 200120 153484 200172 153536
rect 200580 153484 200632 153536
rect 249800 153484 249852 153536
rect 257160 153484 257212 153536
rect 259368 153484 259420 153536
rect 260472 153484 260524 153536
rect 284300 153484 284352 153536
rect 286416 153484 286468 153536
rect 291568 153484 291620 153536
rect 297548 153484 297600 153536
rect 297916 153484 297968 153536
rect 299480 153484 299532 153536
rect 322848 153484 322900 153536
rect 323492 153484 323544 153536
rect 344192 153484 344244 153536
rect 345664 153484 345716 153536
rect 370320 153484 370372 153536
rect 374736 153484 374788 153536
rect 380716 153484 380768 153536
rect 385960 153484 386012 153536
rect 392492 153484 392544 153536
rect 404820 153484 404872 153536
rect 458088 153484 458140 153536
rect 171968 153416 172020 153468
rect 181720 153416 181772 153468
rect 182088 153416 182140 153468
rect 198740 153416 198792 153468
rect 271788 153416 271840 153468
rect 277952 153416 278004 153468
rect 299572 153416 299624 153468
rect 307300 153416 307352 153468
rect 320088 153416 320140 153468
rect 324872 153416 324924 153468
rect 326160 153416 326212 153468
rect 333980 153416 334032 153468
rect 335912 153416 335964 153468
rect 342720 153416 342772 153468
rect 345204 153416 345256 153468
rect 364156 153416 364208 153468
rect 365076 153416 365128 153468
rect 365168 153416 365220 153468
rect 366916 153416 366968 153468
rect 371608 153416 371660 153468
rect 376668 153416 376720 153468
rect 384672 153416 384724 153468
rect 396172 153416 396224 153468
rect 397000 153416 397052 153468
rect 407764 153416 407816 153468
rect 500408 153484 500460 153536
rect 502984 153484 503036 153536
rect 506296 153416 506348 153468
rect 511816 153416 511868 153468
rect 523040 153416 523092 153468
rect 74264 153348 74316 153400
rect 99288 153348 99340 153400
rect 102140 153348 102192 153400
rect 36912 153280 36964 153332
rect 110420 153280 110472 153332
rect 23112 153212 23164 153264
rect 75184 153212 75236 153264
rect 108948 153212 109000 153264
rect 113916 153212 113968 153264
rect 114192 153280 114244 153332
rect 120172 153348 120224 153400
rect 179420 153348 179472 153400
rect 179512 153348 179564 153400
rect 188252 153348 188304 153400
rect 246948 153348 247000 153400
rect 250720 153348 250772 153400
rect 268200 153348 268252 153400
rect 280712 153348 280764 153400
rect 283840 153348 283892 153400
rect 285864 153348 285916 153400
rect 287244 153348 287296 153400
rect 293960 153348 294012 153400
rect 296996 153348 297048 153400
rect 298008 153348 298060 153400
rect 302332 153348 302384 153400
rect 306564 153348 306616 153400
rect 307944 153348 307996 153400
rect 308036 153348 308088 153400
rect 310520 153348 310572 153400
rect 317328 153348 317380 153400
rect 318340 153348 318392 153400
rect 324412 153348 324464 153400
rect 325792 153348 325844 153400
rect 334072 153348 334124 153400
rect 335452 153348 335504 153400
rect 338672 153348 338724 153400
rect 341708 153348 341760 153400
rect 353392 153348 353444 153400
rect 354864 153348 354916 153400
rect 363880 153348 363932 153400
rect 364984 153348 365036 153400
rect 379428 153348 379480 153400
rect 384856 153348 384908 153400
rect 387248 153348 387300 153400
rect 400036 153348 400088 153400
rect 512736 153348 512788 153400
rect 123208 153280 123260 153332
rect 124128 153280 124180 153332
rect 115204 153212 115256 153264
rect 116768 153212 116820 153264
rect 157708 153280 157760 153332
rect 158812 153280 158864 153332
rect 162216 153280 162268 153332
rect 194784 153280 194836 153332
rect 197268 153280 197320 153332
rect 512828 153280 512880 153332
rect 520280 153280 520332 153332
rect 145932 153212 145984 153264
rect 149060 153212 149112 153264
rect 169392 153212 169444 153264
rect 171140 153212 171192 153264
rect 514116 153212 514168 153264
rect 515404 153212 515456 153264
rect 520464 153212 520516 153264
rect 60832 153144 60884 153196
rect 160284 153144 160336 153196
rect 170128 153144 170180 153196
rect 233240 153144 233292 153196
rect 471152 153144 471204 153196
rect 525800 153144 525852 153196
rect 49148 153076 49200 153128
rect 152464 153076 152516 153128
rect 158904 153076 158956 153128
rect 223580 153076 223632 153128
rect 423588 153076 423640 153128
rect 454684 153076 454736 153128
rect 475752 153076 475804 153128
rect 532608 153076 532660 153128
rect 45284 153008 45336 153060
rect 149888 153008 149940 153060
rect 153108 153008 153160 153060
rect 162308 153008 162360 153060
rect 227904 153008 227956 153060
rect 255780 153008 255832 153060
rect 290372 153008 290424 153060
rect 431500 153008 431552 153060
rect 466276 153008 466328 153060
rect 475108 153008 475160 153060
rect 531688 153008 531740 153060
rect 42340 152940 42392 152992
rect 147956 152940 148008 152992
rect 152556 152940 152608 152992
rect 221372 152940 221424 152992
rect 248144 152940 248196 152992
rect 285128 152940 285180 152992
rect 434076 152940 434128 152992
rect 470232 152940 470284 152992
rect 478788 152940 478840 152992
rect 537484 152940 537536 152992
rect 41328 152872 41380 152924
rect 147220 152872 147272 152924
rect 150532 152872 150584 152924
rect 220084 152872 220136 152924
rect 238300 152872 238352 152924
rect 278780 152872 278832 152924
rect 439320 152872 439372 152924
rect 478052 152872 478104 152924
rect 482836 152872 482888 152924
rect 543372 152872 543424 152924
rect 31668 152804 31720 152856
rect 139492 152804 139544 152856
rect 140780 152804 140832 152856
rect 141424 152804 141476 152856
rect 142712 152804 142764 152856
rect 214932 152804 214984 152856
rect 232412 152804 232464 152856
rect 274732 152804 274784 152856
rect 440608 152804 440660 152856
rect 479984 152804 480036 152856
rect 485504 152804 485556 152856
rect 547236 152804 547288 152856
rect 22100 152736 22152 152788
rect 11520 152668 11572 152720
rect 122840 152668 122892 152720
rect 124220 152668 124272 152720
rect 10140 152600 10192 152652
rect 126428 152600 126480 152652
rect 138940 152736 138992 152788
rect 212540 152736 212592 152788
rect 224592 152736 224644 152788
rect 269580 152736 269632 152788
rect 486148 152736 486200 152788
rect 548248 152736 548300 152788
rect 209136 152668 209188 152720
rect 259092 152668 259144 152720
rect 445668 152668 445720 152720
rect 487804 152668 487856 152720
rect 488080 152668 488132 152720
rect 551192 152668 551244 152720
rect 134248 152600 134300 152652
rect 135904 152600 135956 152652
rect 210332 152600 210384 152652
rect 211896 152600 211948 152652
rect 212448 152600 212500 152652
rect 216956 152600 217008 152652
rect 264336 152600 264388 152652
rect 271420 152600 271472 152652
rect 300860 152600 300912 152652
rect 446496 152600 446548 152652
rect 488816 152600 488868 152652
rect 489368 152600 489420 152652
rect 553124 152600 553176 152652
rect 7288 152532 7340 152584
rect 124496 152532 124548 152584
rect 127164 152532 127216 152584
rect 204536 152532 204588 152584
rect 2412 152464 2464 152516
rect 121460 152464 121512 152516
rect 123300 152464 123352 152516
rect 201868 152464 201920 152516
rect 203248 152464 203300 152516
rect 220728 152532 220780 152584
rect 266912 152532 266964 152584
rect 267556 152532 267608 152584
rect 298192 152532 298244 152584
rect 449716 152532 449768 152584
rect 208032 152464 208084 152516
rect 258448 152464 258500 152516
rect 259736 152464 259788 152516
rect 292948 152464 293000 152516
rect 418528 152464 418580 152516
rect 446864 152464 446916 152516
rect 452292 152464 452344 152516
rect 493324 152532 493376 152584
rect 558828 152532 558880 152584
rect 493692 152464 493744 152516
rect 498108 152464 498160 152516
rect 566740 152464 566792 152516
rect 57980 152396 58032 152448
rect 158352 152396 158404 152448
rect 215576 152396 215628 152448
rect 468576 152396 468628 152448
rect 521936 152396 521988 152448
rect 72608 152328 72660 152380
rect 168380 152328 168432 152380
rect 179788 152328 179840 152380
rect 239588 152328 239640 152380
rect 466000 152328 466052 152380
rect 517980 152328 518032 152380
rect 80336 152260 80388 152312
rect 173256 152260 173308 152312
rect 181812 152260 181864 152312
rect 240968 152260 241020 152312
rect 458824 152260 458876 152312
rect 507308 152260 507360 152312
rect 73528 152192 73580 152244
rect 169070 152192 169122 152244
rect 175832 152192 175884 152244
rect 85212 152124 85264 152176
rect 176890 152124 176942 152176
rect 178224 152192 178276 152244
rect 236690 152192 236742 152244
rect 453902 152192 453954 152244
rect 500500 152192 500552 152244
rect 88156 152056 88208 152108
rect 178822 152056 178874 152108
rect 185768 152124 185820 152176
rect 243866 152124 243918 152176
rect 450682 152124 450734 152176
rect 231446 152056 231498 152108
rect 451326 152056 451378 152108
rect 497556 152124 497608 152176
rect 95976 151988 96028 152040
rect 183652 151988 183704 152040
rect 197452 151988 197504 152040
rect 251364 151988 251416 152040
rect 447784 151988 447836 152040
rect 490748 151988 490800 152040
rect 495624 152056 495676 152108
rect 496452 152056 496504 152108
rect 111524 151920 111576 151972
rect 194048 151920 194100 151972
rect 202512 151920 202564 151972
rect 249340 151920 249392 151972
rect 444288 151920 444340 151972
rect 485688 151920 485740 151972
rect 75184 151895 75236 151904
rect 75184 151861 75193 151895
rect 75193 151861 75227 151895
rect 75227 151861 75236 151895
rect 75184 151852 75236 151861
rect 78128 151895 78180 151904
rect 78128 151861 78137 151895
rect 78137 151861 78171 151895
rect 78171 151861 78180 151895
rect 78128 151852 78180 151861
rect 88340 151895 88392 151904
rect 88340 151861 88349 151895
rect 88349 151861 88383 151895
rect 88383 151861 88392 151895
rect 88340 151852 88392 151861
rect 91928 151895 91980 151904
rect 91928 151861 91937 151895
rect 91937 151861 91971 151895
rect 91971 151861 91980 151895
rect 91928 151852 91980 151861
rect 95148 151895 95200 151904
rect 95148 151861 95157 151895
rect 95157 151861 95191 151895
rect 95191 151861 95200 151895
rect 95148 151852 95200 151861
rect 99288 151895 99340 151904
rect 99288 151861 99297 151895
rect 99297 151861 99331 151895
rect 99331 151861 99340 151895
rect 99288 151852 99340 151861
rect 112444 151852 112496 151904
rect 116400 151852 116452 151904
rect 197360 151852 197412 151904
rect 199108 151852 199160 151904
rect 244372 151852 244424 151904
rect 105636 151827 105688 151836
rect 105636 151793 105645 151827
rect 105645 151793 105679 151827
rect 105679 151793 105688 151827
rect 105636 151784 105688 151793
rect 146484 151784 146536 151836
rect 25504 151716 25556 151768
rect 127716 151716 127768 151768
rect 212448 151784 212500 151836
rect 252008 151784 252060 151836
rect 503628 151784 503680 151836
rect 520556 151784 520608 151836
rect 212908 151716 212960 151768
rect 64420 151648 64472 151700
rect 171140 151648 171192 151700
rect 505008 151648 505060 151700
rect 528560 151648 528612 151700
rect 50620 151580 50672 151632
rect 197268 151580 197320 151632
rect 506940 151623 506992 151632
rect 506940 151589 506949 151623
rect 506949 151589 506983 151623
rect 506983 151589 506992 151623
rect 506940 151580 506992 151589
rect 3056 151512 3108 151564
rect 117044 151512 117096 151564
rect 118332 151512 118384 151564
rect 3240 151444 3292 151496
rect 40132 151419 40184 151428
rect 40132 151385 40141 151419
rect 40141 151385 40175 151419
rect 40175 151385 40184 151419
rect 40132 151376 40184 151385
rect 43812 151376 43864 151428
rect 115388 151376 115440 151428
rect 117136 151444 117188 151496
rect 503720 151512 503772 151564
rect 505652 151512 505704 151564
rect 545120 151512 545172 151564
rect 575480 151444 575532 151496
rect 117320 151376 117372 151428
rect 118424 151376 118476 151428
rect 575572 151376 575624 151428
rect 3424 151308 3476 151360
rect 115020 151308 115072 151360
rect 116952 151308 117004 151360
rect 507768 151308 507820 151360
rect 508872 151351 508924 151360
rect 508872 151317 508881 151351
rect 508881 151317 508915 151351
rect 508915 151317 508924 151351
rect 508872 151308 508924 151317
rect 4804 151240 4856 151292
rect 112628 151240 112680 151292
rect 114008 151240 114060 151292
rect 515404 151308 515456 151360
rect 518624 151308 518676 151360
rect 519268 151308 519320 151360
rect 520372 151308 520424 151360
rect 520648 151240 520700 151292
rect 521752 151104 521804 151156
rect 5172 151036 5224 151088
rect 521844 150968 521896 151020
rect 522304 150900 522356 150952
rect 3884 150832 3936 150884
rect 112720 150832 112772 150884
rect 4160 150764 4212 150816
rect 114284 150764 114336 150816
rect 3700 150696 3752 150748
rect 114376 150696 114428 150748
rect 117320 150696 117372 150748
rect 118608 150696 118660 150748
rect 3424 150628 3476 150680
rect 115112 150628 115164 150680
rect 119528 150560 119580 150612
rect 113364 150492 113416 150544
rect 117228 150424 117280 150476
rect 3792 150356 3844 150408
rect 112536 150356 112588 150408
rect 4068 150288 4120 150340
rect 115848 150288 115900 150340
rect 3976 150220 4028 150272
rect 115756 150220 115808 150272
rect 3516 147636 3568 147688
rect 5172 147636 5224 147688
rect 113364 147568 113416 147620
rect 117320 147568 117372 147620
rect 3608 145936 3660 145988
rect 4160 145936 4212 145988
rect 3516 140768 3568 140820
rect 4804 140768 4856 140820
rect 115388 136552 115440 136604
rect 117688 136552 117740 136604
rect 115388 129752 115440 129804
rect 117320 129752 117372 129804
rect 114928 127984 114980 128036
rect 117780 127984 117832 128036
rect 115572 124176 115624 124228
rect 117320 124176 117372 124228
rect 114192 111800 114244 111852
rect 117872 111800 117924 111852
rect 115020 104796 115072 104848
rect 117504 104796 117556 104848
rect 112720 102756 112772 102808
rect 117688 102756 117740 102808
rect 116308 99424 116360 99476
rect 119712 99424 119764 99476
rect 112628 99288 112680 99340
rect 115112 99288 115164 99340
rect 115020 96568 115072 96620
rect 117504 96568 117556 96620
rect 115112 95140 115164 95192
rect 117872 95140 117924 95192
rect 114376 88816 114428 88868
rect 118608 88816 118660 88868
rect 115848 86912 115900 86964
rect 117320 86912 117372 86964
rect 112536 85008 112588 85060
rect 117780 85008 117832 85060
rect 115756 84124 115808 84176
rect 117320 84124 117372 84176
rect 114284 73108 114336 73160
rect 117320 73108 117372 73160
rect 112444 67532 112496 67584
rect 117320 67532 117372 67584
rect 116308 67396 116360 67448
rect 119896 67396 119948 67448
rect 115756 58828 115808 58880
rect 117872 58828 117924 58880
rect 115848 56176 115900 56228
rect 117320 56176 117372 56228
rect 115112 53796 115164 53848
rect 118608 53796 118660 53848
rect 522580 52368 522632 52420
rect 114284 48220 114336 48272
rect 117412 48288 117464 48340
rect 114468 46860 114520 46912
rect 117320 46928 117372 46980
rect 114376 45704 114428 45756
rect 117320 45704 117372 45756
rect 115020 39448 115072 39500
rect 118516 39448 118568 39500
rect 113732 37204 113784 37256
rect 117320 37272 117372 37324
rect 114836 34552 114888 34604
rect 117872 34552 117924 34604
rect 114928 34484 114980 34536
rect 117228 34484 117280 34536
rect 3700 33804 3752 33856
rect 4804 33804 4856 33856
rect 3792 31016 3844 31068
rect 4896 31016 4948 31068
rect 114744 30336 114796 30388
rect 117320 30336 117372 30388
rect 112536 29520 112588 29572
rect 114836 29520 114888 29572
rect 112444 29452 112496 29504
rect 114928 29452 114980 29504
rect 4068 28908 4120 28960
rect 4988 28908 5040 28960
rect 116492 20816 116544 20868
rect 119896 20816 119948 20868
rect 3976 20612 4028 20664
rect 5080 20612 5132 20664
rect 3424 19252 3476 19304
rect 5172 19252 5224 19304
rect 114836 16600 114888 16652
rect 117504 16600 117556 16652
rect 114744 13812 114796 13864
rect 117320 13812 117372 13864
rect 3516 11840 3568 11892
rect 5264 11840 5316 11892
rect 117964 11704 118016 11756
rect 118332 11704 118384 11756
rect 3608 11636 3660 11688
rect 3884 11636 3936 11688
rect 114652 11024 114704 11076
rect 117320 11024 117372 11076
rect 3332 9596 3384 9648
rect 5448 9596 5500 9648
rect 114560 7216 114612 7268
rect 117320 7216 117372 7268
rect 3516 6468 3568 6520
rect 4344 6468 4396 6520
rect 2872 5856 2924 5908
rect 118608 5856 118660 5908
rect 2964 5788 3016 5840
rect 118516 5788 118568 5840
rect 3700 5720 3752 5772
rect 117872 5720 117924 5772
rect 3148 5652 3200 5704
rect 117136 5652 117188 5704
rect 3884 5584 3936 5636
rect 117780 5584 117832 5636
rect 3056 5516 3108 5568
rect 114928 5516 114980 5568
rect 3424 5448 3476 5500
rect 114744 5448 114796 5500
rect 3240 5380 3292 5432
rect 114560 5380 114612 5432
rect 4804 5312 4856 5364
rect 115756 5312 115808 5364
rect 4068 5244 4120 5296
rect 114836 5244 114888 5296
rect 117044 5244 117096 5296
rect 520924 5244 520976 5296
rect 3976 5176 4028 5228
rect 114652 5176 114704 5228
rect 5172 5108 5224 5160
rect 115848 5108 115900 5160
rect 119896 5108 119948 5160
rect 576860 5108 576912 5160
rect 520740 5040 520792 5092
rect 521844 4972 521896 5024
rect 4896 4904 4948 4956
rect 115112 4904 115164 4956
rect 118700 4904 118752 4956
rect 577228 4904 577280 4956
rect 522028 4836 522080 4888
rect 522396 4768 522448 4820
rect 3608 4700 3660 4752
rect 113732 4700 113784 4752
rect 5080 4632 5132 4684
rect 114468 4632 114520 4684
rect 444380 4675 444432 4684
rect 444380 4641 444389 4675
rect 444389 4641 444423 4675
rect 444423 4641 444432 4675
rect 444380 4632 444432 4641
rect 463332 4675 463384 4684
rect 463332 4641 463341 4675
rect 463341 4641 463375 4675
rect 463375 4641 463384 4675
rect 463332 4632 463384 4641
rect 5264 4564 5316 4616
rect 114284 4564 114336 4616
rect 4344 4496 4396 4548
rect 114376 4496 114428 4548
rect 12164 4471 12216 4480
rect 12164 4437 12173 4471
rect 12173 4437 12207 4471
rect 12207 4437 12216 4471
rect 12164 4428 12216 4437
rect 48228 4428 48280 4480
rect 118424 4428 118476 4480
rect 62672 4403 62724 4412
rect 62672 4369 62681 4403
rect 62681 4369 62715 4403
rect 62715 4369 62724 4403
rect 62672 4360 62724 4369
rect 71964 4360 72016 4412
rect 74908 4360 74960 4412
rect 79324 4403 79376 4412
rect 79324 4369 79333 4403
rect 79333 4369 79367 4403
rect 79367 4369 79376 4403
rect 79324 4360 79376 4369
rect 82176 4360 82228 4412
rect 82820 4360 82872 4412
rect 85948 4360 86000 4412
rect 116676 4360 116728 4412
rect 81992 4292 82044 4344
rect 86408 4292 86460 4344
rect 95976 4335 96028 4344
rect 95976 4301 95985 4335
rect 95985 4301 96019 4335
rect 96019 4301 96028 4335
rect 95976 4292 96028 4301
rect 106188 4292 106240 4344
rect 118240 4292 118292 4344
rect 3332 4224 3384 4276
rect 112444 4224 112496 4276
rect 2964 4156 3016 4208
rect 117320 4156 117372 4208
rect 45928 4088 45980 4140
rect 522212 4088 522264 4140
rect 61108 4020 61160 4072
rect 111800 4020 111852 4072
rect 114284 4020 114336 4072
rect 176752 4020 176804 4072
rect 383292 4020 383344 4072
rect 460112 4020 460164 4072
rect 103612 3952 103664 4004
rect 167368 3952 167420 4004
rect 367928 3952 367980 4004
rect 433524 3952 433576 4004
rect 93032 3884 93084 3936
rect 165528 3884 165580 3936
rect 172796 3884 172848 3936
rect 216818 3884 216870 3936
rect 268568 3884 268620 3936
rect 272202 3884 272254 3936
rect 273904 3884 273956 3936
rect 275330 3884 275382 3936
rect 281494 3884 281546 3936
rect 284576 3884 284628 3936
rect 379934 3884 379986 3936
rect 454776 3884 454828 3936
rect 82360 3816 82412 3868
rect 156512 3816 156564 3868
rect 188804 3816 188856 3868
rect 225788 3816 225840 3868
rect 361396 3816 361448 3868
rect 422852 3816 422904 3868
rect 427820 3816 427872 3868
rect 555884 3816 555936 3868
rect 87696 3748 87748 3800
rect 162768 3748 162820 3800
rect 183468 3748 183520 3800
rect 222660 3748 222712 3800
rect 371056 3748 371108 3800
rect 438860 3748 438912 3800
rect 77024 3680 77076 3732
rect 153108 3680 153160 3732
rect 178132 3680 178184 3732
rect 219624 3680 219676 3732
rect 373908 3680 373960 3732
rect 444196 3748 444248 3800
rect 454684 3748 454736 3800
rect 534632 3748 534684 3800
rect 443736 3680 443788 3732
rect 539968 3680 540020 3732
rect 71688 3612 71740 3664
rect 149152 3612 149204 3664
rect 167460 3612 167512 3664
rect 213460 3612 213512 3664
rect 324872 3612 324924 3664
rect 359004 3612 359056 3664
rect 386328 3612 386380 3664
rect 465448 3612 465500 3664
rect 66444 3544 66496 3596
rect 146116 3544 146168 3596
rect 162216 3544 162268 3596
rect 210332 3544 210384 3596
rect 318708 3544 318760 3596
rect 348424 3544 348476 3596
rect 389088 3544 389140 3596
rect 470784 3544 470836 3596
rect 55956 3476 56008 3528
rect 118056 3476 118108 3528
rect 151544 3476 151596 3528
rect 204260 3476 204312 3528
rect 343364 3476 343416 3528
rect 390928 3476 390980 3528
rect 392584 3476 392636 3528
rect 476120 3476 476172 3528
rect 98368 3408 98420 3460
rect 173440 3408 173492 3460
rect 337200 3408 337252 3460
rect 380348 3408 380400 3460
rect 395620 3408 395672 3460
rect 481456 3408 481508 3460
rect 522948 3408 523000 3460
rect 566556 3408 566608 3460
rect 42616 3340 42668 3392
rect 117596 3340 117648 3392
rect 119712 3340 119764 3392
rect 146208 3340 146260 3392
rect 201132 3340 201184 3392
rect 204720 3340 204772 3392
rect 234988 3340 235040 3392
rect 247408 3340 247460 3392
rect 259644 3340 259696 3392
rect 309508 3340 309560 3392
rect 332416 3340 332468 3392
rect 352564 3340 352616 3392
rect 404912 3340 404964 3392
rect 407764 3340 407816 3392
rect 486700 3340 486752 3392
rect 29184 3272 29236 3324
rect 136640 3272 136692 3324
rect 140872 3272 140924 3324
rect 198096 3272 198148 3324
rect 199384 3272 199436 3324
rect 231952 3272 232004 3324
rect 358728 3272 358780 3324
rect 417332 3272 417384 3324
rect 492036 3272 492088 3324
rect 518624 3272 518676 3324
rect 520556 3272 520608 3324
rect 23848 3204 23900 3256
rect 133420 3204 133472 3256
rect 135536 3204 135588 3256
rect 194968 3204 195020 3256
rect 226064 3204 226116 3256
rect 247316 3204 247368 3256
rect 306196 3204 306248 3256
rect 327080 3204 327132 3256
rect 331036 3204 331088 3256
rect 369676 3204 369728 3256
rect 398748 3204 398800 3256
rect 407764 3204 407816 3256
rect 497372 3204 497424 3256
rect 18512 3136 18564 3188
rect 130384 3136 130436 3188
rect 13176 3068 13228 3120
rect 127256 3068 127308 3120
rect 130292 3068 130344 3120
rect 191932 3136 191984 3188
rect 215392 3136 215444 3188
rect 241152 3136 241204 3188
rect 333888 3136 333940 3188
rect 375012 3136 375064 3188
rect 406936 3136 406988 3188
rect 502616 3136 502668 3188
rect 7840 3000 7892 3052
rect 124220 3000 124272 3052
rect 2596 2932 2648 2984
rect 121460 2932 121512 2984
rect 124956 2932 125008 2984
rect 189080 3068 189132 3120
rect 210056 3068 210108 3120
rect 238024 3068 238076 3120
rect 241980 3068 242032 3120
rect 256608 3068 256660 3120
rect 321468 3068 321520 3120
rect 353760 3068 353812 3120
rect 364892 3068 364944 3120
rect 428188 3068 428240 3120
rect 438676 3068 438728 3120
rect 550548 3068 550600 3120
rect 185768 3000 185820 3052
rect 231308 3000 231360 3052
rect 250352 3000 250404 3052
rect 257988 3000 258040 3052
rect 265716 3000 265768 3052
rect 312544 3000 312596 3052
rect 337752 3000 337804 3052
rect 340236 3000 340288 3052
rect 385684 3000 385736 3052
rect 401416 3000 401468 3052
rect 407948 3000 408000 3052
rect 423312 3000 423364 3052
rect 561220 3000 561272 3052
rect 156880 2932 156932 2984
rect 207296 2932 207348 2984
rect 220728 2932 220780 2984
rect 244280 2932 244332 2984
rect 252652 2932 252704 2984
rect 262680 2932 262732 2984
rect 315672 2932 315724 2984
rect 343088 2932 343140 2984
rect 346308 2932 346360 2984
rect 396264 2932 396316 2984
rect 426348 2932 426400 2984
rect 571892 2932 571944 2984
rect 45100 2864 45152 2916
rect 50344 2864 50396 2916
rect 52368 2864 52420 2916
rect 522120 2864 522172 2916
rect 34520 2796 34572 2848
rect 44180 2796 44232 2848
rect 108948 2796 109000 2848
rect 179604 2796 179656 2848
rect 194140 2796 194192 2848
rect 229100 2796 229152 2848
rect 236644 2796 236696 2848
rect 19248 2728 19300 2780
rect 106188 2728 106240 2780
rect 111800 2728 111852 2780
rect 152004 2728 152056 2780
rect 153108 2728 153160 2780
rect 161112 2728 161164 2780
rect 28908 2660 28960 2712
rect 119344 2660 119396 2712
rect 156512 2660 156564 2712
rect 164240 2728 164292 2780
rect 165528 2728 165580 2780
rect 170404 2728 170456 2780
rect 176752 2728 176804 2780
rect 182640 2728 182692 2780
rect 263232 2796 263284 2848
rect 253480 2728 253532 2780
rect 269120 2728 269172 2780
rect 284852 2728 284904 2780
rect 289636 2796 289688 2848
rect 287980 2728 288032 2780
rect 295156 2796 295208 2848
rect 303344 2796 303396 2848
rect 321836 2796 321888 2848
rect 327908 2796 327960 2848
rect 364340 2796 364392 2848
rect 377220 2796 377272 2848
rect 449532 2796 449584 2848
rect 484308 2796 484360 2848
rect 523960 2796 524012 2848
rect 417148 2728 417200 2780
rect 454684 2728 454736 2780
rect 162768 2660 162820 2712
rect 167276 2660 167328 2712
rect 167368 2660 167420 2712
rect 176660 2660 176712 2712
rect 420276 2660 420328 2712
rect 427820 2660 427872 2712
rect 435640 2660 435692 2712
rect 443736 2660 443788 2712
rect 1308 2592 1360 2644
rect 58624 2592 58676 2644
rect 75828 2592 75880 2644
rect 499672 2592 499724 2644
rect 6000 2524 6052 2576
rect 48228 2524 48280 2576
rect 68928 2524 68980 2576
rect 490380 2524 490432 2576
rect 89352 2456 89404 2508
rect 502708 2456 502760 2508
rect 92388 2388 92440 2440
rect 505744 2388 505796 2440
rect 108856 2320 108908 2372
rect 520648 2320 520700 2372
rect 112628 2252 112680 2304
rect 520372 2252 520424 2304
rect 106004 2184 106056 2236
rect 512000 2184 512052 2236
rect 22652 2116 22704 2168
rect 113824 2116 113876 2168
rect 114376 2116 114428 2168
rect 115296 2116 115348 2168
rect 32588 2048 32640 2100
rect 115388 2048 115440 2100
rect 119528 2116 119580 2168
rect 515036 2116 515088 2168
rect 508872 2048 508924 2100
rect 44180 1980 44232 2032
rect 432144 1980 432196 2032
rect 9312 1912 9364 1964
rect 114008 1912 114060 1964
rect 114100 1912 114152 1964
rect 115572 1844 115624 1896
rect 99288 1776 99340 1828
rect 114192 1776 114244 1828
rect 114376 1776 114428 1828
rect 116584 1912 116636 1964
rect 496820 1912 496872 1964
rect 493416 1844 493468 1896
rect 487344 1776 487396 1828
rect 39764 1708 39816 1760
rect 139584 1708 139636 1760
rect 149152 1708 149204 1760
rect 158076 1708 158128 1760
rect 278688 1708 278740 1760
rect 279240 1708 279292 1760
rect 291016 1708 291068 1760
rect 300492 1708 300544 1760
rect 50344 1640 50396 1692
rect 142712 1640 142764 1692
rect 146116 1640 146168 1692
rect 154948 1640 155000 1692
rect 300216 1640 300268 1692
rect 316500 1708 316552 1760
rect 349528 1708 349580 1760
rect 401600 1708 401652 1760
rect 410984 1708 411036 1760
rect 513380 1708 513432 1760
rect 50436 1572 50488 1624
rect 145748 1572 145800 1624
rect 293868 1572 293920 1624
rect 305828 1572 305880 1624
rect 55772 1504 55824 1556
rect 149060 1504 149112 1556
rect 297180 1504 297232 1556
rect 311164 1640 311216 1692
rect 355600 1640 355652 1692
rect 412272 1640 412324 1692
rect 429108 1640 429160 1692
rect 508044 1640 508096 1692
rect 413928 1572 413980 1624
rect 484308 1572 484360 1624
rect 15936 1436 15988 1488
rect 520832 1436 520884 1488
rect 25964 1368 26016 1420
rect 468852 1368 468904 1420
rect 39304 1300 39356 1352
rect 478052 1300 478104 1352
rect 116768 1232 116820 1284
rect 459652 1232 459704 1284
rect 116860 1164 116912 1216
rect 453488 1164 453540 1216
rect 119896 1096 119948 1148
rect 441160 1096 441212 1148
<< metal2 >>
rect 478 159200 534 160000
rect 1398 159200 1454 160000
rect 2410 159200 2466 160000
rect 3330 159200 3386 160000
rect 4342 159200 4398 160000
rect 5262 159200 5318 160000
rect 6274 159200 6330 160000
rect 7286 159200 7342 160000
rect 8206 159200 8262 160000
rect 9218 159200 9274 160000
rect 10138 159200 10194 160000
rect 11150 159200 11206 160000
rect 12162 159200 12218 160000
rect 13082 159200 13138 160000
rect 14094 159200 14150 160000
rect 15014 159200 15070 160000
rect 16026 159200 16082 160000
rect 17038 159200 17094 160000
rect 17958 159200 18014 160000
rect 18970 159200 19026 160000
rect 19890 159200 19946 160000
rect 20902 159200 20958 160000
rect 21914 159200 21970 160000
rect 22834 159200 22890 160000
rect 23846 159200 23902 160000
rect 24766 159200 24822 160000
rect 25778 159200 25834 160000
rect 26790 159200 26846 160000
rect 27710 159200 27766 160000
rect 28722 159200 28778 160000
rect 29642 159200 29698 160000
rect 30654 159200 30710 160000
rect 31666 159200 31722 160000
rect 32586 159200 32642 160000
rect 33598 159200 33654 160000
rect 34518 159200 34574 160000
rect 35530 159200 35586 160000
rect 36542 159200 36598 160000
rect 37462 159200 37518 160000
rect 38474 159200 38530 160000
rect 39394 159200 39450 160000
rect 40406 159200 40462 160000
rect 41326 159200 41382 160000
rect 42338 159200 42394 160000
rect 43350 159200 43406 160000
rect 44270 159200 44326 160000
rect 45282 159200 45338 160000
rect 46202 159200 46258 160000
rect 47214 159200 47270 160000
rect 48226 159200 48282 160000
rect 49146 159200 49202 160000
rect 50158 159200 50214 160000
rect 51078 159200 51134 160000
rect 52090 159200 52146 160000
rect 53102 159200 53158 160000
rect 54022 159200 54078 160000
rect 55034 159200 55090 160000
rect 55954 159200 56010 160000
rect 56966 159200 57022 160000
rect 57978 159200 58034 160000
rect 58898 159200 58954 160000
rect 59910 159200 59966 160000
rect 60830 159200 60886 160000
rect 61842 159200 61898 160000
rect 62854 159200 62910 160000
rect 63774 159200 63830 160000
rect 64786 159200 64842 160000
rect 65706 159200 65762 160000
rect 66718 159200 66774 160000
rect 67730 159200 67786 160000
rect 68650 159200 68706 160000
rect 69662 159200 69718 160000
rect 70582 159200 70638 160000
rect 71594 159200 71650 160000
rect 72606 159200 72662 160000
rect 73526 159200 73582 160000
rect 74538 159200 74594 160000
rect 75458 159200 75514 160000
rect 76470 159200 76526 160000
rect 77482 159200 77538 160000
rect 78402 159200 78458 160000
rect 79414 159200 79470 160000
rect 80334 159200 80390 160000
rect 81346 159200 81402 160000
rect 82266 159200 82322 160000
rect 83278 159200 83334 160000
rect 84290 159200 84346 160000
rect 85210 159200 85266 160000
rect 86222 159200 86278 160000
rect 87142 159200 87198 160000
rect 88154 159200 88210 160000
rect 89166 159200 89222 160000
rect 90086 159200 90142 160000
rect 91098 159200 91154 160000
rect 92018 159200 92074 160000
rect 93030 159200 93086 160000
rect 94042 159200 94098 160000
rect 94962 159200 95018 160000
rect 95974 159200 96030 160000
rect 96894 159200 96950 160000
rect 97906 159200 97962 160000
rect 98918 159200 98974 160000
rect 99838 159200 99894 160000
rect 100850 159200 100906 160000
rect 101770 159200 101826 160000
rect 102782 159200 102838 160000
rect 103794 159200 103850 160000
rect 104714 159200 104770 160000
rect 105726 159200 105782 160000
rect 106646 159200 106702 160000
rect 107658 159200 107714 160000
rect 108670 159200 108726 160000
rect 109590 159200 109646 160000
rect 110602 159200 110658 160000
rect 111522 159200 111578 160000
rect 112534 159200 112590 160000
rect 113546 159200 113602 160000
rect 114466 159200 114522 160000
rect 115478 159200 115534 160000
rect 116398 159200 116454 160000
rect 117410 159200 117466 160000
rect 118330 159200 118386 160000
rect 119342 159200 119398 160000
rect 120354 159200 120410 160000
rect 121274 159200 121330 160000
rect 122286 159200 122342 160000
rect 123206 159200 123262 160000
rect 124218 159200 124274 160000
rect 125230 159200 125286 160000
rect 126150 159200 126206 160000
rect 127162 159200 127218 160000
rect 128082 159200 128138 160000
rect 129094 159200 129150 160000
rect 130106 159200 130162 160000
rect 131026 159200 131082 160000
rect 132038 159200 132094 160000
rect 132958 159200 133014 160000
rect 133970 159200 134026 160000
rect 134982 159200 135038 160000
rect 135902 159200 135958 160000
rect 136914 159202 136970 160000
rect 137020 159310 137232 159338
rect 137020 159202 137048 159310
rect 136914 159200 137048 159202
rect 492 154902 520 159200
rect 480 154896 532 154902
rect 480 154838 532 154844
rect 1308 154896 1360 154902
rect 1308 154838 1360 154844
rect 1320 153542 1348 154838
rect 1412 153882 1440 159200
rect 1400 153876 1452 153882
rect 1400 153818 1452 153824
rect 1308 153536 1360 153542
rect 1308 153478 1360 153484
rect 1320 2650 1348 153478
rect 2424 152522 2452 159200
rect 3344 156641 3372 159200
rect 3422 157584 3478 157593
rect 3422 157519 3478 157528
rect 3330 156632 3386 156641
rect 3330 156567 3386 156576
rect 2412 152516 2464 152522
rect 2412 152458 2464 152464
rect 3056 151564 3108 151570
rect 3056 151506 3108 151512
rect 3068 148481 3096 151506
rect 3240 151496 3292 151502
rect 3240 151438 3292 151444
rect 3054 148472 3110 148481
rect 3054 148407 3110 148416
rect 3252 139369 3280 151438
rect 3436 151366 3464 157519
rect 4356 155242 4384 159200
rect 5276 155854 5304 159200
rect 6288 156670 6316 159200
rect 6276 156664 6328 156670
rect 6276 156606 6328 156612
rect 5264 155848 5316 155854
rect 5264 155790 5316 155796
rect 4344 155236 4396 155242
rect 4344 155178 4396 155184
rect 5998 153232 6054 153241
rect 5998 153167 6054 153176
rect 3514 152960 3570 152969
rect 3514 152895 3570 152904
rect 3528 152289 3556 152895
rect 3514 152280 3570 152289
rect 3514 152215 3570 152224
rect 6012 151994 6040 153167
rect 7300 152590 7328 159200
rect 8220 155281 8248 159200
rect 9232 155310 9260 159200
rect 9220 155304 9272 155310
rect 8206 155272 8262 155281
rect 9220 155246 9272 155252
rect 8206 155207 8262 155216
rect 10152 152658 10180 159200
rect 11164 158710 11192 159200
rect 11152 158704 11204 158710
rect 11152 158646 11204 158652
rect 12176 155446 12204 159200
rect 12164 155440 12216 155446
rect 12164 155382 12216 155388
rect 11520 155236 11572 155242
rect 11520 155178 11572 155184
rect 11532 152726 11560 155178
rect 13096 154329 13124 159200
rect 14108 155922 14136 159200
rect 15028 157826 15056 159200
rect 15016 157820 15068 157826
rect 15016 157762 15068 157768
rect 14096 155916 14148 155922
rect 14096 155858 14148 155864
rect 16040 155242 16068 159200
rect 16028 155236 16080 155242
rect 16028 155178 16080 155184
rect 13082 154320 13138 154329
rect 13082 154255 13138 154264
rect 17052 153950 17080 159200
rect 17972 156738 18000 159200
rect 18984 158302 19012 159200
rect 18972 158296 19024 158302
rect 18972 158238 19024 158244
rect 17960 156732 18012 156738
rect 17960 156674 18012 156680
rect 19904 155417 19932 159200
rect 19890 155408 19946 155417
rect 19890 155343 19946 155352
rect 20916 154018 20944 159200
rect 21928 154714 21956 159200
rect 22848 158642 22876 159200
rect 22836 158636 22888 158642
rect 22836 158578 22888 158584
rect 23860 155378 23888 159200
rect 23848 155372 23900 155378
rect 23848 155314 23900 155320
rect 21928 154686 22140 154714
rect 20904 154012 20956 154018
rect 20904 153954 20956 153960
rect 17040 153944 17092 153950
rect 17040 153886 17092 153892
rect 22112 152794 22140 154686
rect 24780 154086 24808 159200
rect 25792 156777 25820 159200
rect 26804 158778 26832 159200
rect 26792 158772 26844 158778
rect 26792 158714 26844 158720
rect 25778 156768 25834 156777
rect 25778 156703 25834 156712
rect 27724 155446 27752 159200
rect 25504 155440 25556 155446
rect 25504 155382 25556 155388
rect 27712 155440 27764 155446
rect 27712 155382 27764 155388
rect 24768 154080 24820 154086
rect 24768 154022 24820 154028
rect 23112 153264 23164 153270
rect 23112 153206 23164 153212
rect 22100 152788 22152 152794
rect 22100 152730 22152 152736
rect 11520 152720 11572 152726
rect 11520 152662 11572 152668
rect 10140 152652 10192 152658
rect 10140 152594 10192 152600
rect 7288 152584 7340 152590
rect 7288 152526 7340 152532
rect 23124 151994 23152 153206
rect 5704 151966 6040 151994
rect 22816 151966 23152 151994
rect 25516 151774 25544 155382
rect 28736 154465 28764 159200
rect 29656 155514 29684 159200
rect 30668 158846 30696 159200
rect 30656 158840 30708 158846
rect 30656 158782 30708 158788
rect 31680 155650 31708 159200
rect 31668 155644 31720 155650
rect 31668 155586 31720 155592
rect 32600 155514 32628 159200
rect 33612 156806 33640 159200
rect 34532 158914 34560 159200
rect 34520 158908 34572 158914
rect 34520 158850 34572 158856
rect 33600 156800 33652 156806
rect 33600 156742 33652 156748
rect 35544 155582 35572 159200
rect 35532 155576 35584 155582
rect 35532 155518 35584 155524
rect 29644 155508 29696 155514
rect 29644 155450 29696 155456
rect 31668 155508 31720 155514
rect 31668 155450 31720 155456
rect 32588 155508 32640 155514
rect 32588 155450 32640 155456
rect 28722 154456 28778 154465
rect 28722 154391 28778 154400
rect 30010 153504 30066 153513
rect 30010 153439 30066 153448
rect 26606 153368 26662 153377
rect 26606 153303 26662 153312
rect 26620 151994 26648 153303
rect 30024 151994 30052 153439
rect 31680 152862 31708 155450
rect 36556 154154 36584 159200
rect 36544 154148 36596 154154
rect 36544 154090 36596 154096
rect 36912 153332 36964 153338
rect 36912 153274 36964 153280
rect 31668 152856 31720 152862
rect 31668 152798 31720 152804
rect 33506 152008 33562 152017
rect 26312 151966 26648 151994
rect 29716 151966 30052 151994
rect 33212 151966 33506 151994
rect 36924 151994 36952 153274
rect 37476 152561 37504 159200
rect 38488 158982 38516 159200
rect 38476 158976 38528 158982
rect 38476 158918 38528 158924
rect 39408 155106 39436 159200
rect 40420 155718 40448 159200
rect 40408 155712 40460 155718
rect 40408 155654 40460 155660
rect 39396 155100 39448 155106
rect 39396 155042 39448 155048
rect 41340 152930 41368 159200
rect 42352 152998 42380 159200
rect 43364 157894 43392 159200
rect 43352 157888 43404 157894
rect 43352 157830 43404 157836
rect 44284 155922 44312 159200
rect 44272 155916 44324 155922
rect 44272 155858 44324 155864
rect 45296 153066 45324 159200
rect 46216 156874 46244 159200
rect 47228 157962 47256 159200
rect 47216 157956 47268 157962
rect 47216 157898 47268 157904
rect 46204 156868 46256 156874
rect 46204 156810 46256 156816
rect 48240 154222 48268 159200
rect 48228 154216 48280 154222
rect 48228 154158 48280 154164
rect 49160 153134 49188 159200
rect 49148 153128 49200 153134
rect 49148 153070 49200 153076
rect 45284 153060 45336 153066
rect 45284 153002 45336 153008
rect 42340 152992 42392 152998
rect 42340 152934 42392 152940
rect 41328 152924 41380 152930
rect 41328 152866 41380 152872
rect 50172 152697 50200 159200
rect 51092 158030 51120 159200
rect 51080 158024 51132 158030
rect 51080 157966 51132 157972
rect 52104 155174 52132 159200
rect 52092 155168 52144 155174
rect 52092 155110 52144 155116
rect 53116 154290 53144 159200
rect 54036 156942 54064 159200
rect 55048 158522 55076 159200
rect 55048 158494 55260 158522
rect 55232 158370 55260 158494
rect 55220 158364 55272 158370
rect 55220 158306 55272 158312
rect 54024 156936 54076 156942
rect 54024 156878 54076 156884
rect 55968 155786 55996 159200
rect 55956 155780 56008 155786
rect 55956 155722 56008 155728
rect 56980 154698 57008 159200
rect 56968 154692 57020 154698
rect 56968 154634 57020 154640
rect 53104 154284 53156 154290
rect 53104 154226 53156 154232
rect 57518 153640 57574 153649
rect 57518 153575 57574 153584
rect 50158 152688 50214 152697
rect 50158 152623 50214 152632
rect 37462 152552 37518 152561
rect 37462 152487 37518 152496
rect 57532 151994 57560 153575
rect 57992 152454 58020 159200
rect 58912 158098 58940 159200
rect 58900 158092 58952 158098
rect 58900 158034 58952 158040
rect 59924 154426 59952 159200
rect 59912 154420 59964 154426
rect 59912 154362 59964 154368
rect 60844 153202 60872 159200
rect 61856 156913 61884 159200
rect 62868 158438 62896 159200
rect 62856 158432 62908 158438
rect 62856 158374 62908 158380
rect 61842 156904 61898 156913
rect 61842 156839 61898 156848
rect 63788 155553 63816 159200
rect 63774 155544 63830 155553
rect 63774 155479 63830 155488
rect 64800 154358 64828 159200
rect 64788 154352 64840 154358
rect 64788 154294 64840 154300
rect 60832 153196 60884 153202
rect 60832 153138 60884 153144
rect 65720 152833 65748 159200
rect 66732 158506 66760 159200
rect 66720 158500 66772 158506
rect 66720 158442 66772 158448
rect 67744 155689 67772 159200
rect 68664 157010 68692 159200
rect 69676 157078 69704 159200
rect 70596 158574 70624 159200
rect 70584 158568 70636 158574
rect 70584 158510 70636 158516
rect 69664 157072 69716 157078
rect 69664 157014 69716 157020
rect 68652 157004 68704 157010
rect 68652 156946 68704 156952
rect 67730 155680 67786 155689
rect 67730 155615 67786 155624
rect 71608 154494 71636 159200
rect 71596 154488 71648 154494
rect 71596 154430 71648 154436
rect 65706 152824 65762 152833
rect 65706 152759 65762 152768
rect 57980 152448 58032 152454
rect 57980 152390 58032 152396
rect 72620 152386 72648 159200
rect 72608 152380 72660 152386
rect 72608 152322 72660 152328
rect 73540 152250 73568 159200
rect 74552 154970 74580 159200
rect 74540 154964 74592 154970
rect 74540 154906 74592 154912
rect 75472 154562 75500 159200
rect 76484 157146 76512 159200
rect 77496 157214 77524 159200
rect 77484 157208 77536 157214
rect 77484 157150 77536 157156
rect 76472 157140 76524 157146
rect 76472 157082 76524 157088
rect 78416 154766 78444 159200
rect 79428 155961 79456 159200
rect 79414 155952 79470 155961
rect 79414 155887 79470 155896
rect 78404 154760 78456 154766
rect 78404 154702 78456 154708
rect 75460 154556 75512 154562
rect 75460 154498 75512 154504
rect 74264 153400 74316 153406
rect 74264 153342 74316 153348
rect 73528 152244 73580 152250
rect 73528 152186 73580 152192
rect 67500 152144 67556 152153
rect 67500 152079 67556 152088
rect 36616 151966 36952 151994
rect 57224 151966 57560 151994
rect 67514 151980 67542 152079
rect 33506 151943 33562 151952
rect 25504 151768 25556 151774
rect 74276 151722 74304 153342
rect 75184 153264 75236 153270
rect 75184 153206 75236 153212
rect 75196 151910 75224 153206
rect 80348 152318 80376 159200
rect 81360 157049 81388 159200
rect 82280 157282 82308 159200
rect 82268 157276 82320 157282
rect 82268 157218 82320 157224
rect 81346 157040 81402 157049
rect 81346 156975 81402 156984
rect 83292 153814 83320 159200
rect 84304 157350 84332 159200
rect 84292 157344 84344 157350
rect 84292 157286 84344 157292
rect 85026 153912 85082 153921
rect 85026 153847 85082 153856
rect 83280 153808 83332 153814
rect 81162 153776 81218 153785
rect 83280 153750 83332 153756
rect 81162 153711 81218 153720
rect 80336 152312 80388 152318
rect 80336 152254 80388 152260
rect 75184 151904 75236 151910
rect 78128 151904 78180 151910
rect 75184 151846 75236 151852
rect 77832 151852 78128 151858
rect 77832 151846 78180 151852
rect 77832 151830 78168 151846
rect 81176 151722 81204 153711
rect 85040 151994 85068 153847
rect 85224 152182 85252 159200
rect 86236 155038 86264 159200
rect 87156 155825 87184 159200
rect 87142 155816 87198 155825
rect 87142 155751 87198 155760
rect 86224 155032 86276 155038
rect 86224 154974 86276 154980
rect 85212 152176 85264 152182
rect 85212 152118 85264 152124
rect 88168 152114 88196 159200
rect 89180 154630 89208 159200
rect 90100 158166 90128 159200
rect 90088 158160 90140 158166
rect 90088 158102 90140 158108
rect 89168 154624 89220 154630
rect 89168 154566 89220 154572
rect 91112 153678 91140 159200
rect 92032 156602 92060 159200
rect 92020 156596 92072 156602
rect 92020 156538 92072 156544
rect 93044 153746 93072 159200
rect 93032 153740 93084 153746
rect 93032 153682 93084 153688
rect 91100 153672 91152 153678
rect 91100 153614 91152 153620
rect 94056 152969 94084 159200
rect 94976 154834 95004 159200
rect 94964 154828 95016 154834
rect 94964 154770 95016 154776
rect 94042 152960 94098 152969
rect 94042 152895 94098 152904
rect 88156 152108 88208 152114
rect 88156 152050 88208 152056
rect 95988 152046 96016 159200
rect 96908 156058 96936 159200
rect 96896 156052 96948 156058
rect 96896 155994 96948 156000
rect 97920 154902 97948 159200
rect 97908 154896 97960 154902
rect 97908 154838 97960 154844
rect 98826 154048 98882 154057
rect 98826 153983 98882 153992
rect 84732 151966 85068 151994
rect 95976 152040 96028 152046
rect 98840 151994 98868 153983
rect 98932 153610 98960 159200
rect 99852 156534 99880 159200
rect 100864 157486 100892 159200
rect 100852 157480 100904 157486
rect 100852 157422 100904 157428
rect 101784 157185 101812 159200
rect 101770 157176 101826 157185
rect 101770 157111 101826 157120
rect 99840 156528 99892 156534
rect 99840 156470 99892 156476
rect 102140 155848 102192 155854
rect 102140 155790 102192 155796
rect 98920 153604 98972 153610
rect 98920 153546 98972 153552
rect 102152 153406 102180 155790
rect 102796 154873 102824 159200
rect 103808 156466 103836 159200
rect 104728 158234 104756 159200
rect 104716 158228 104768 158234
rect 104716 158170 104768 158176
rect 103796 156460 103848 156466
rect 103796 156402 103848 156408
rect 105740 156398 105768 159200
rect 105728 156392 105780 156398
rect 105728 156334 105780 156340
rect 106660 155145 106688 159200
rect 107672 156330 107700 159200
rect 108684 157554 108712 159200
rect 108672 157548 108724 157554
rect 108672 157490 108724 157496
rect 107660 156324 107712 156330
rect 107660 156266 107712 156272
rect 106646 155136 106702 155145
rect 106646 155071 106702 155080
rect 102782 154864 102838 154873
rect 102782 154799 102838 154808
rect 109604 154737 109632 159200
rect 110616 155854 110644 159200
rect 110604 155848 110656 155854
rect 110604 155790 110656 155796
rect 110420 154760 110472 154766
rect 109590 154728 109646 154737
rect 110420 154702 110472 154708
rect 109590 154663 109646 154672
rect 99288 153400 99340 153406
rect 99288 153342 99340 153348
rect 102140 153400 102192 153406
rect 102140 153342 102192 153348
rect 95976 151982 96028 151988
rect 98532 151966 98868 151994
rect 99300 151910 99328 153342
rect 110432 153338 110460 154702
rect 110420 153332 110472 153338
rect 110420 153274 110472 153280
rect 108948 153264 109000 153270
rect 108948 153206 109000 153212
rect 108960 151994 108988 153206
rect 108836 151966 108988 151994
rect 111536 151978 111564 159200
rect 112548 156126 112576 159200
rect 112536 156120 112588 156126
rect 112536 156062 112588 156068
rect 113180 155848 113232 155854
rect 113180 155790 113232 155796
rect 113192 154578 113220 155790
rect 113560 154766 113588 159200
rect 114480 155009 114508 159200
rect 115492 156262 115520 159200
rect 115480 156256 115532 156262
rect 115480 156198 115532 156204
rect 114466 155000 114522 155009
rect 114466 154935 114522 154944
rect 113548 154760 113600 154766
rect 113548 154702 113600 154708
rect 113192 154550 114048 154578
rect 112534 154184 112590 154193
rect 112534 154119 112590 154128
rect 112548 151994 112576 154119
rect 114020 153320 114048 154550
rect 114192 153332 114244 153338
rect 114020 153292 114192 153320
rect 114192 153274 114244 153280
rect 113916 153264 113968 153270
rect 113916 153206 113968 153212
rect 115204 153264 115256 153270
rect 115204 153206 115256 153212
rect 113822 152144 113878 152153
rect 113822 152079 113878 152088
rect 111524 151972 111576 151978
rect 112240 151966 112576 151994
rect 111524 151914 111576 151920
rect 88340 151904 88392 151910
rect 88228 151852 88340 151858
rect 91928 151904 91980 151910
rect 88228 151846 88392 151852
rect 91632 151852 91928 151858
rect 95148 151904 95200 151910
rect 91632 151846 91980 151852
rect 95036 151852 95148 151858
rect 95036 151846 95200 151852
rect 99288 151904 99340 151910
rect 112444 151904 112496 151910
rect 102046 151872 102102 151881
rect 99288 151846 99340 151852
rect 88228 151830 88380 151846
rect 91632 151830 91968 151846
rect 95036 151830 95188 151846
rect 101936 151830 102046 151858
rect 105340 151842 105676 151858
rect 112444 151846 112496 151852
rect 105340 151836 105688 151842
rect 105340 151830 105636 151836
rect 102046 151807 102102 151816
rect 105636 151778 105688 151784
rect 25504 151710 25556 151716
rect 64124 151706 64460 151722
rect 64124 151700 64472 151706
rect 64124 151694 64420 151700
rect 74276 151694 74428 151722
rect 81176 151694 81328 151722
rect 64420 151642 64472 151648
rect 50620 151632 50672 151638
rect 50324 151580 50620 151586
rect 50324 151574 50672 151580
rect 50324 151558 50660 151574
rect 71318 151464 71374 151473
rect 40020 151434 40172 151450
rect 43516 151434 43852 151450
rect 40020 151428 40184 151434
rect 40020 151422 40132 151428
rect 43516 151428 43864 151434
rect 43516 151422 43812 151428
rect 40132 151370 40184 151376
rect 71024 151422 71318 151450
rect 71318 151399 71374 151408
rect 43812 151370 43864 151376
rect 3424 151360 3476 151366
rect 9402 151328 9458 151337
rect 3424 151302 3476 151308
rect 4804 151292 4856 151298
rect 9108 151286 9402 151314
rect 12806 151328 12862 151337
rect 12512 151286 12806 151314
rect 9402 151263 9458 151272
rect 16302 151328 16358 151337
rect 16008 151286 16302 151314
rect 12806 151263 12862 151272
rect 19706 151328 19762 151337
rect 19412 151286 19706 151314
rect 16302 151263 16358 151272
rect 47030 151328 47086 151337
rect 46920 151286 47030 151314
rect 19706 151263 19762 151272
rect 53930 151328 53986 151337
rect 53820 151286 53930 151314
rect 47030 151263 47086 151272
rect 60830 151328 60886 151337
rect 60720 151286 60830 151314
rect 53930 151263 53986 151272
rect 60830 151263 60886 151272
rect 4804 151234 4856 151240
rect 3884 150884 3936 150890
rect 3884 150826 3936 150832
rect 3700 150748 3752 150754
rect 3700 150690 3752 150696
rect 3424 150680 3476 150686
rect 3424 150622 3476 150628
rect 3330 149968 3386 149977
rect 3330 149903 3386 149912
rect 3238 139360 3294 139369
rect 3238 139295 3294 139304
rect 3344 134745 3372 149903
rect 3436 143857 3464 150622
rect 3516 147688 3568 147694
rect 3516 147630 3568 147636
rect 3422 143848 3478 143857
rect 3422 143783 3478 143792
rect 3528 142154 3556 147630
rect 3608 145988 3660 145994
rect 3608 145930 3660 145936
rect 3436 142126 3556 142154
rect 3330 134736 3386 134745
rect 3330 134671 3386 134680
rect 3436 98161 3464 142126
rect 3516 140820 3568 140826
rect 3516 140762 3568 140768
rect 3528 102785 3556 140762
rect 3620 107273 3648 145930
rect 3712 111897 3740 150690
rect 3792 150408 3844 150414
rect 3792 150350 3844 150356
rect 3804 116521 3832 150350
rect 3896 121009 3924 150826
rect 4160 150816 4212 150822
rect 4160 150758 4212 150764
rect 4068 150340 4120 150346
rect 4068 150282 4120 150288
rect 3976 150272 4028 150278
rect 3976 150214 4028 150220
rect 3988 125633 4016 150214
rect 4080 130121 4108 150282
rect 4172 145994 4200 150758
rect 4160 145988 4212 145994
rect 4160 145930 4212 145936
rect 4816 140826 4844 151234
rect 5172 151088 5224 151094
rect 5172 151030 5224 151036
rect 5184 147694 5212 151030
rect 5172 147688 5224 147694
rect 5172 147630 5224 147636
rect 4804 140820 4856 140826
rect 4804 140762 4856 140768
rect 4066 130112 4122 130121
rect 4066 130047 4122 130056
rect 3974 125624 4030 125633
rect 3974 125559 4030 125568
rect 3882 121000 3938 121009
rect 3882 120935 3938 120944
rect 3790 116512 3846 116521
rect 3790 116447 3846 116456
rect 3698 111888 3754 111897
rect 3698 111823 3754 111832
rect 3606 107264 3662 107273
rect 3606 107199 3662 107208
rect 3514 102776 3570 102785
rect 3514 102711 3570 102720
rect 3422 98152 3478 98161
rect 3422 98087 3478 98096
rect 3698 93664 3754 93673
rect 3698 93599 3754 93608
rect 3422 84416 3478 84425
rect 3422 84351 3478 84360
rect 3330 57080 3386 57089
rect 3330 57015 3386 57024
rect 3238 52456 3294 52465
rect 3238 52391 3294 52400
rect 3146 47968 3202 47977
rect 3146 47903 3202 47912
rect 3054 43344 3110 43353
rect 3054 43279 3110 43288
rect 2962 38720 3018 38729
rect 2962 38655 3018 38664
rect 2870 34232 2926 34241
rect 2870 34167 2926 34176
rect 2884 5914 2912 34167
rect 2872 5908 2924 5914
rect 2872 5850 2924 5856
rect 2976 5846 3004 38655
rect 2964 5840 3016 5846
rect 2964 5782 3016 5788
rect 3068 5574 3096 43279
rect 3160 5710 3188 47903
rect 3252 6914 3280 52391
rect 3344 9654 3372 57015
rect 3436 19310 3464 84351
rect 3514 70816 3570 70825
rect 3514 70751 3570 70760
rect 3424 19304 3476 19310
rect 3424 19246 3476 19252
rect 3422 15872 3478 15881
rect 3422 15807 3478 15816
rect 3332 9648 3384 9654
rect 3332 9590 3384 9596
rect 3252 6886 3372 6914
rect 3238 6760 3294 6769
rect 3238 6695 3294 6704
rect 3148 5704 3200 5710
rect 3148 5646 3200 5652
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 3252 5438 3280 6695
rect 3240 5432 3292 5438
rect 3240 5374 3292 5380
rect 3344 4282 3372 6886
rect 3436 5506 3464 15807
rect 3528 11898 3556 70751
rect 3606 66192 3662 66201
rect 3606 66127 3662 66136
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3620 11778 3648 66127
rect 3712 33862 3740 93599
rect 3790 89040 3846 89049
rect 3790 88975 3846 88984
rect 3700 33856 3752 33862
rect 3700 33798 3752 33804
rect 3804 31074 3832 88975
rect 4066 79928 4122 79937
rect 4066 79863 4122 79872
rect 3974 75304 4030 75313
rect 3974 75239 4030 75248
rect 3882 61568 3938 61577
rect 3882 61503 3938 61512
rect 3792 31068 3844 31074
rect 3792 31010 3844 31016
rect 3698 29608 3754 29617
rect 3698 29543 3754 29552
rect 3528 11750 3648 11778
rect 3528 6526 3556 11750
rect 3608 11688 3660 11694
rect 3608 11630 3660 11636
rect 3516 6520 3568 6526
rect 3516 6462 3568 6468
rect 3424 5500 3476 5506
rect 3424 5442 3476 5448
rect 3620 4758 3648 11630
rect 3712 5778 3740 29543
rect 3790 25120 3846 25129
rect 3790 25055 3846 25064
rect 3804 6914 3832 25055
rect 3896 11694 3924 61503
rect 3988 20670 4016 75239
rect 4080 28966 4108 79863
rect 112456 67590 112484 151846
rect 112628 151292 112680 151298
rect 112628 151234 112680 151240
rect 112536 150408 112588 150414
rect 112536 150350 112588 150356
rect 112548 85066 112576 150350
rect 112640 99346 112668 151234
rect 112720 150884 112772 150890
rect 112720 150826 112772 150832
rect 112732 102814 112760 150826
rect 113364 150544 113416 150550
rect 113364 150486 113416 150492
rect 113376 147626 113404 150486
rect 113364 147620 113416 147626
rect 113364 147562 113416 147568
rect 112720 102808 112772 102814
rect 112720 102750 112772 102756
rect 112628 99340 112680 99346
rect 112628 99282 112680 99288
rect 112536 85060 112588 85066
rect 112536 85002 112588 85008
rect 112444 67584 112496 67590
rect 112444 67526 112496 67532
rect 113732 37256 113784 37262
rect 113732 37198 113784 37204
rect 4804 33856 4856 33862
rect 4804 33798 4856 33804
rect 4068 28960 4120 28966
rect 4068 28902 4120 28908
rect 3976 20664 4028 20670
rect 3976 20606 4028 20612
rect 4066 20496 4122 20505
rect 4066 20431 4122 20440
rect 3884 11688 3936 11694
rect 3884 11630 3936 11636
rect 3974 11384 4030 11393
rect 3974 11319 4030 11328
rect 3804 6886 3924 6914
rect 3700 5772 3752 5778
rect 3700 5714 3752 5720
rect 3896 5642 3924 6886
rect 3884 5636 3936 5642
rect 3884 5578 3936 5584
rect 3988 5234 4016 11319
rect 4080 5302 4108 20431
rect 4344 6520 4396 6526
rect 4344 6462 4396 6468
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 3608 4752 3660 4758
rect 3608 4694 3660 4700
rect 4356 4554 4384 6462
rect 4816 5370 4844 33798
rect 4896 31068 4948 31074
rect 4896 31010 4948 31016
rect 4804 5364 4856 5370
rect 4804 5306 4856 5312
rect 4908 4962 4936 31010
rect 112536 29572 112588 29578
rect 112536 29514 112588 29520
rect 112444 29504 112496 29510
rect 112444 29446 112496 29452
rect 4988 28960 5040 28966
rect 4988 28902 5040 28908
rect 5000 6089 5028 28902
rect 5080 20664 5132 20670
rect 5080 20606 5132 20612
rect 4986 6080 5042 6089
rect 4986 6015 5042 6024
rect 4896 4956 4948 4962
rect 4896 4898 4948 4904
rect 5092 4690 5120 20606
rect 5172 19304 5224 19310
rect 5172 19246 5224 19252
rect 5184 5166 5212 19246
rect 5264 11892 5316 11898
rect 5264 11834 5316 11840
rect 5172 5160 5224 5166
rect 5172 5102 5224 5108
rect 5080 4684 5132 4690
rect 5080 4626 5132 4632
rect 5276 4622 5304 11834
rect 5448 9648 5500 9654
rect 5448 9590 5500 9596
rect 5460 5953 5488 9590
rect 5446 5944 5502 5953
rect 5446 5879 5502 5888
rect 5264 4616 5316 4622
rect 35806 4584 35862 4593
rect 5264 4558 5316 4564
rect 4344 4548 4396 4554
rect 35696 4542 35806 4570
rect 65982 4584 66038 4593
rect 65688 4542 65982 4570
rect 35806 4519 35862 4528
rect 65982 4519 66038 4528
rect 71962 4584 72018 4593
rect 72422 4584 72478 4593
rect 72312 4542 72422 4570
rect 71962 4519 72018 4528
rect 72422 4519 72478 4528
rect 74906 4584 74962 4593
rect 74906 4519 74962 4528
rect 81990 4584 82046 4593
rect 81990 4519 82046 4528
rect 82174 4584 82230 4593
rect 82634 4584 82690 4593
rect 82340 4542 82634 4570
rect 82174 4519 82230 4528
rect 82634 4519 82690 4528
rect 82818 4584 82874 4593
rect 82818 4519 82874 4528
rect 86406 4584 86462 4593
rect 102690 4584 102746 4593
rect 102396 4542 102690 4570
rect 86406 4519 86462 4528
rect 102690 4519 102746 4528
rect 4344 4490 4396 4496
rect 12164 4480 12216 4486
rect 48228 4480 48280 4486
rect 12216 4428 12328 4434
rect 12164 4422 12328 4428
rect 48228 4422 48280 4428
rect 12176 4406 12328 4422
rect 3332 4276 3384 4282
rect 3332 4218 3384 4224
rect 2964 4208 3016 4214
rect 2964 4150 3016 4156
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 1308 2644 1360 2650
rect 1308 2586 1360 2592
rect 2608 800 2636 2926
rect 2976 2281 3004 4150
rect 5704 4134 6040 4162
rect 9016 4134 9352 4162
rect 15640 4134 15976 4162
rect 18952 4134 19288 4162
rect 22356 4134 22692 4162
rect 25668 4134 26004 4162
rect 6012 2582 6040 4134
rect 7840 3052 7892 3058
rect 7840 2994 7892 3000
rect 6000 2576 6052 2582
rect 6000 2518 6052 2524
rect 2962 2272 3018 2281
rect 2962 2207 3018 2216
rect 7852 800 7880 2994
rect 9324 1970 9352 4134
rect 13176 3120 13228 3126
rect 13176 3062 13228 3068
rect 9312 1964 9364 1970
rect 9312 1906 9364 1912
rect 13188 800 13216 3062
rect 15948 1494 15976 4134
rect 18512 3188 18564 3194
rect 18512 3130 18564 3136
rect 15936 1488 15988 1494
rect 15936 1430 15988 1436
rect 18524 800 18552 3130
rect 19260 2786 19288 4134
rect 19248 2780 19300 2786
rect 19248 2722 19300 2728
rect 22664 2174 22692 4134
rect 23848 3256 23900 3262
rect 23848 3198 23900 3204
rect 22652 2168 22704 2174
rect 22652 2110 22704 2116
rect 23860 800 23888 3198
rect 25976 1426 26004 4134
rect 28966 3890 28994 4148
rect 32292 4134 32628 4162
rect 39008 4134 39344 4162
rect 42320 4134 42656 4162
rect 45632 4146 45968 4162
rect 45632 4140 45980 4146
rect 45632 4134 45928 4140
rect 28920 3862 28994 3890
rect 28920 2718 28948 3862
rect 29184 3324 29236 3330
rect 29184 3266 29236 3272
rect 28908 2712 28960 2718
rect 28908 2654 28960 2660
rect 25964 1420 26016 1426
rect 25964 1362 26016 1368
rect 29196 800 29224 3266
rect 32600 2106 32628 4134
rect 34520 2848 34572 2854
rect 34520 2790 34572 2796
rect 32588 2100 32640 2106
rect 32588 2042 32640 2048
rect 34532 800 34560 2790
rect 39316 1358 39344 4134
rect 42628 3398 42656 4134
rect 45928 4082 45980 4088
rect 42616 3392 42668 3398
rect 42616 3334 42668 3340
rect 45100 2916 45152 2922
rect 45100 2858 45152 2864
rect 44180 2848 44232 2854
rect 44180 2790 44232 2796
rect 44192 2038 44220 2790
rect 44180 2032 44232 2038
rect 44180 1974 44232 1980
rect 39764 1760 39816 1766
rect 39764 1702 39816 1708
rect 39304 1352 39356 1358
rect 39304 1294 39356 1300
rect 39776 800 39804 1702
rect 45112 800 45140 2858
rect 48240 2582 48268 4422
rect 62376 4418 62712 4434
rect 71976 4418 72004 4519
rect 74920 4418 74948 4519
rect 79028 4418 79364 4434
rect 62376 4412 62724 4418
rect 62376 4406 62672 4412
rect 62672 4354 62724 4360
rect 71964 4412 72016 4418
rect 71964 4354 72016 4360
rect 74908 4412 74960 4418
rect 79028 4412 79376 4418
rect 79028 4406 79324 4412
rect 74908 4354 74960 4360
rect 79324 4354 79376 4360
rect 82004 4350 82032 4519
rect 82188 4418 82216 4519
rect 82832 4418 82860 4519
rect 85652 4418 85988 4434
rect 82176 4412 82228 4418
rect 82176 4354 82228 4360
rect 82820 4412 82872 4418
rect 85652 4412 86000 4418
rect 85652 4406 85948 4412
rect 82820 4354 82872 4360
rect 85948 4354 86000 4360
rect 86420 4350 86448 4519
rect 81992 4344 82044 4350
rect 81992 4286 82044 4292
rect 86408 4344 86460 4350
rect 95976 4344 96028 4350
rect 86408 4286 86460 4292
rect 95680 4292 95976 4298
rect 95680 4286 96028 4292
rect 106188 4344 106240 4350
rect 106188 4286 106240 4292
rect 95680 4270 96016 4286
rect 49036 4134 49372 4162
rect 49344 2825 49372 4134
rect 52334 3890 52362 4148
rect 55660 4134 55996 4162
rect 52334 3862 52408 3890
rect 52380 2922 52408 3862
rect 55968 3534 55996 4134
rect 58636 4134 58972 4162
rect 55956 3528 56008 3534
rect 55956 3470 56008 3476
rect 50344 2916 50396 2922
rect 50344 2858 50396 2864
rect 52368 2916 52420 2922
rect 52368 2858 52420 2864
rect 49330 2816 49386 2825
rect 49330 2751 49386 2760
rect 48228 2576 48280 2582
rect 48228 2518 48280 2524
rect 50356 1698 50384 2858
rect 58636 2650 58664 4134
rect 61108 4072 61160 4078
rect 61108 4014 61160 4020
rect 58624 2644 58676 2650
rect 58624 2586 58676 2592
rect 50344 1692 50396 1698
rect 50344 1634 50396 1640
rect 50436 1624 50488 1630
rect 50436 1566 50488 1572
rect 50448 800 50476 1566
rect 55772 1556 55824 1562
rect 55772 1498 55824 1504
rect 55784 800 55812 1498
rect 61120 800 61148 4014
rect 68986 3890 69014 4148
rect 75716 4134 75868 4162
rect 89056 4134 89392 4162
rect 68940 3862 69014 3890
rect 66444 3596 66496 3602
rect 66444 3538 66496 3544
rect 66456 800 66484 3538
rect 68940 2582 68968 3862
rect 71688 3664 71740 3670
rect 71688 3606 71740 3612
rect 68928 2576 68980 2582
rect 68928 2518 68980 2524
rect 71700 800 71728 3606
rect 75840 2650 75868 4134
rect 82360 3868 82412 3874
rect 82360 3810 82412 3816
rect 77024 3732 77076 3738
rect 77024 3674 77076 3680
rect 75828 2644 75880 2650
rect 75828 2586 75880 2592
rect 77036 800 77064 3674
rect 82372 800 82400 3810
rect 87696 3800 87748 3806
rect 87696 3742 87748 3748
rect 87708 800 87736 3742
rect 89364 2514 89392 4134
rect 92354 3890 92382 4148
rect 98992 4134 99328 4162
rect 105708 4134 106044 4162
rect 93032 3936 93084 3942
rect 92354 3862 92428 3890
rect 93032 3878 93084 3884
rect 89352 2508 89404 2514
rect 89352 2450 89404 2456
rect 92400 2446 92428 3862
rect 92388 2440 92440 2446
rect 92388 2382 92440 2388
rect 93044 800 93072 3878
rect 98368 3460 98420 3466
rect 98368 3402 98420 3408
rect 98380 800 98408 3402
rect 99300 1834 99328 4134
rect 103612 4004 103664 4010
rect 103612 3946 103664 3952
rect 99288 1828 99340 1834
rect 99288 1770 99340 1776
rect 103624 800 103652 3946
rect 106016 2242 106044 4134
rect 106200 2786 106228 4286
rect 112456 4282 112484 29446
rect 112548 5953 112576 29514
rect 112534 5944 112590 5953
rect 112534 5879 112590 5888
rect 113744 4758 113772 37198
rect 113732 4752 113784 4758
rect 113732 4694 113784 4700
rect 112444 4276 112496 4282
rect 112444 4218 112496 4224
rect 108868 4134 109020 4162
rect 112332 4134 112668 4162
rect 106188 2780 106240 2786
rect 106188 2722 106240 2728
rect 108868 2378 108896 4134
rect 111800 4072 111852 4078
rect 111800 4014 111852 4020
rect 108948 2848 109000 2854
rect 108948 2790 109000 2796
rect 108856 2372 108908 2378
rect 108856 2314 108908 2320
rect 106004 2236 106056 2242
rect 106004 2178 106056 2184
rect 108960 800 108988 2790
rect 111812 2786 111840 4014
rect 111800 2780 111852 2786
rect 111800 2722 111852 2728
rect 112640 2310 112668 4134
rect 112628 2304 112680 2310
rect 112628 2246 112680 2252
rect 113836 2174 113864 152079
rect 113928 2961 113956 153206
rect 114926 152280 114982 152289
rect 114926 152215 114982 152224
rect 114098 151328 114154 151337
rect 114008 151292 114060 151298
rect 114098 151263 114154 151272
rect 114008 151234 114060 151240
rect 113914 2952 113970 2961
rect 113914 2887 113970 2896
rect 113824 2168 113876 2174
rect 113824 2110 113876 2116
rect 114020 1970 114048 151234
rect 114112 1970 114140 151263
rect 114284 150816 114336 150822
rect 114284 150758 114336 150764
rect 114192 111852 114244 111858
rect 114192 111794 114244 111800
rect 114008 1964 114060 1970
rect 114008 1906 114060 1912
rect 114100 1964 114152 1970
rect 114100 1906 114152 1912
rect 114204 1834 114232 111794
rect 114296 73166 114324 150758
rect 114376 150748 114428 150754
rect 114376 150690 114428 150696
rect 114388 88874 114416 150690
rect 114940 128042 114968 152215
rect 115020 151360 115072 151366
rect 115020 151302 115072 151308
rect 114928 128036 114980 128042
rect 114928 127978 114980 127984
rect 115032 104854 115060 151302
rect 115112 150680 115164 150686
rect 115112 150622 115164 150628
rect 115020 104848 115072 104854
rect 115020 104790 115072 104796
rect 115124 103514 115152 150622
rect 115032 103486 115152 103514
rect 115032 96626 115060 103486
rect 115112 99340 115164 99346
rect 115112 99282 115164 99288
rect 115020 96620 115072 96626
rect 115020 96562 115072 96568
rect 115124 95198 115152 99282
rect 115112 95192 115164 95198
rect 115112 95134 115164 95140
rect 114376 88868 114428 88874
rect 114376 88810 114428 88816
rect 114284 73160 114336 73166
rect 114284 73102 114336 73108
rect 115112 53848 115164 53854
rect 115112 53790 115164 53796
rect 114284 48272 114336 48278
rect 114284 48214 114336 48220
rect 114296 4622 114324 48214
rect 114468 46912 114520 46918
rect 114468 46854 114520 46860
rect 114376 45756 114428 45762
rect 114376 45698 114428 45704
rect 114284 4616 114336 4622
rect 114284 4558 114336 4564
rect 114388 4554 114416 45698
rect 114480 4690 114508 46854
rect 115020 39500 115072 39506
rect 115020 39442 115072 39448
rect 114836 34604 114888 34610
rect 114836 34546 114888 34552
rect 114744 30388 114796 30394
rect 114744 30330 114796 30336
rect 114756 26234 114784 30330
rect 114848 29578 114876 34546
rect 114928 34536 114980 34542
rect 114928 34478 114980 34484
rect 114836 29572 114888 29578
rect 114836 29514 114888 29520
rect 114940 29510 114968 34478
rect 114928 29504 114980 29510
rect 114928 29446 114980 29452
rect 114756 26206 114968 26234
rect 114836 16652 114888 16658
rect 114836 16594 114888 16600
rect 114744 13864 114796 13870
rect 114744 13806 114796 13812
rect 114652 11076 114704 11082
rect 114652 11018 114704 11024
rect 114560 7268 114612 7274
rect 114560 7210 114612 7216
rect 114572 5438 114600 7210
rect 114560 5432 114612 5438
rect 114560 5374 114612 5380
rect 114664 5234 114692 11018
rect 114756 5506 114784 13806
rect 114744 5500 114796 5506
rect 114744 5442 114796 5448
rect 114848 5302 114876 16594
rect 114940 5574 114968 26206
rect 115032 6089 115060 39442
rect 115018 6080 115074 6089
rect 115018 6015 115074 6024
rect 114928 5568 114980 5574
rect 114928 5510 114980 5516
rect 114836 5296 114888 5302
rect 114836 5238 114888 5244
rect 114652 5228 114704 5234
rect 114652 5170 114704 5176
rect 115124 4962 115152 53790
rect 115112 4956 115164 4962
rect 115112 4898 115164 4904
rect 114468 4684 114520 4690
rect 114468 4626 114520 4632
rect 114376 4548 114428 4554
rect 114376 4490 114428 4496
rect 114284 4072 114336 4078
rect 114284 4014 114336 4020
rect 114192 1828 114244 1834
rect 114192 1770 114244 1776
rect 114296 800 114324 4014
rect 115216 3097 115244 153206
rect 115478 152008 115534 152017
rect 115478 151943 115534 151952
rect 115294 151872 115350 151881
rect 115294 151807 115350 151816
rect 115202 3088 115258 3097
rect 115202 3023 115258 3032
rect 115308 2174 115336 151807
rect 115388 151428 115440 151434
rect 115388 151370 115440 151376
rect 115400 136610 115428 151370
rect 115388 136604 115440 136610
rect 115388 136546 115440 136552
rect 115388 129804 115440 129810
rect 115388 129746 115440 129752
rect 114376 2168 114428 2174
rect 114376 2110 114428 2116
rect 115296 2168 115348 2174
rect 115296 2110 115348 2116
rect 114388 1834 114416 2110
rect 115400 2106 115428 129746
rect 115492 2417 115520 151943
rect 116412 151910 116440 159200
rect 117424 157622 117452 159200
rect 117412 157616 117464 157622
rect 117412 157558 117464 157564
rect 118344 155854 118372 159200
rect 119356 156194 119384 159200
rect 119436 157412 119488 157418
rect 119436 157354 119488 157360
rect 119344 156188 119396 156194
rect 119344 156130 119396 156136
rect 118332 155848 118384 155854
rect 118332 155790 118384 155796
rect 116768 154692 116820 154698
rect 116768 154634 116820 154640
rect 116780 153270 116808 154634
rect 116768 153264 116820 153270
rect 116768 153206 116820 153212
rect 118238 152416 118294 152425
rect 118238 152351 118294 152360
rect 116400 151904 116452 151910
rect 116400 151846 116452 151852
rect 117044 151564 117096 151570
rect 117044 151506 117096 151512
rect 116582 151464 116638 151473
rect 116582 151399 116638 151408
rect 115662 150648 115718 150657
rect 115662 150583 115718 150592
rect 115572 124228 115624 124234
rect 115572 124170 115624 124176
rect 115478 2408 115534 2417
rect 115478 2343 115534 2352
rect 115388 2100 115440 2106
rect 115388 2042 115440 2048
rect 115584 1902 115612 124170
rect 115676 2009 115704 150583
rect 115848 150340 115900 150346
rect 115848 150282 115900 150288
rect 115756 150272 115808 150278
rect 115756 150214 115808 150220
rect 115768 84182 115796 150214
rect 115860 86970 115888 150282
rect 116306 100600 116362 100609
rect 116306 100535 116362 100544
rect 116320 99482 116348 100535
rect 116308 99476 116360 99482
rect 116308 99418 116360 99424
rect 115848 86964 115900 86970
rect 115848 86906 115900 86912
rect 115756 84176 115808 84182
rect 115756 84118 115808 84124
rect 116308 67448 116360 67454
rect 116308 67390 116360 67396
rect 116320 66473 116348 67390
rect 116306 66464 116362 66473
rect 116306 66399 116362 66408
rect 115756 58880 115808 58886
rect 115756 58822 115808 58828
rect 115768 5370 115796 58822
rect 115848 56228 115900 56234
rect 115848 56170 115900 56176
rect 115756 5364 115808 5370
rect 115756 5306 115808 5312
rect 115860 5166 115888 56170
rect 116490 20904 116546 20913
rect 116490 20839 116492 20848
rect 116544 20839 116546 20848
rect 116492 20810 116544 20816
rect 115848 5160 115900 5166
rect 115848 5102 115900 5108
rect 115662 2000 115718 2009
rect 116596 1970 116624 151399
rect 116952 151360 117004 151366
rect 116952 151302 117004 151308
rect 116674 141672 116730 141681
rect 116674 141607 116730 141616
rect 116688 4418 116716 141607
rect 116766 134736 116822 134745
rect 116766 134671 116822 134680
rect 116676 4412 116728 4418
rect 116676 4354 116728 4360
rect 115662 1935 115718 1944
rect 116584 1964 116636 1970
rect 116584 1906 116636 1912
rect 115572 1896 115624 1902
rect 115572 1838 115624 1844
rect 114376 1828 114428 1834
rect 114376 1770 114428 1776
rect 116780 1290 116808 134671
rect 116858 123312 116914 123321
rect 116858 123247 116914 123256
rect 116768 1284 116820 1290
rect 116768 1226 116820 1232
rect 116872 1222 116900 123247
rect 116964 112033 116992 151302
rect 116950 112024 117006 112033
rect 116950 111959 117006 111968
rect 116950 109848 117006 109857
rect 116950 109783 117006 109792
rect 116964 9625 116992 109783
rect 117056 98841 117084 151506
rect 117136 151496 117188 151502
rect 117136 151438 117188 151444
rect 117148 146169 117176 151438
rect 117320 151428 117372 151434
rect 117320 151370 117372 151376
rect 117332 150754 117360 151370
rect 118146 150784 118202 150793
rect 117320 150748 117372 150754
rect 118146 150719 118202 150728
rect 117320 150690 117372 150696
rect 117962 150512 118018 150521
rect 117228 150476 117280 150482
rect 117962 150447 118018 150456
rect 117228 150418 117280 150424
rect 117134 146160 117190 146169
rect 117134 146095 117190 146104
rect 117240 144809 117268 150418
rect 117870 150376 117926 150385
rect 117870 150311 117926 150320
rect 117320 147620 117372 147626
rect 117320 147562 117372 147568
rect 117332 147529 117360 147562
rect 117318 147520 117374 147529
rect 117318 147455 117374 147464
rect 117226 144800 117282 144809
rect 117226 144735 117282 144744
rect 117688 136604 117740 136610
rect 117688 136546 117740 136552
rect 117700 136513 117728 136546
rect 117686 136504 117742 136513
rect 117686 136439 117742 136448
rect 117594 132968 117650 132977
rect 117594 132903 117650 132912
rect 117318 130112 117374 130121
rect 117318 130047 117374 130056
rect 117332 129810 117360 130047
rect 117320 129804 117372 129810
rect 117320 129746 117372 129752
rect 117318 124264 117374 124273
rect 117318 124199 117320 124208
rect 117372 124199 117374 124208
rect 117320 124170 117372 124176
rect 117504 104848 117556 104854
rect 117504 104790 117556 104796
rect 117516 104689 117544 104790
rect 117502 104680 117558 104689
rect 117502 104615 117558 104624
rect 117042 98832 117098 98841
rect 117042 98767 117098 98776
rect 117504 96620 117556 96626
rect 117504 96562 117556 96568
rect 117516 95985 117544 96562
rect 117502 95976 117558 95985
rect 117502 95911 117558 95920
rect 117608 93854 117636 132903
rect 117780 128036 117832 128042
rect 117780 127978 117832 127984
rect 117792 103514 117820 127978
rect 117884 111858 117912 150311
rect 117872 111852 117924 111858
rect 117872 111794 117924 111800
rect 117792 103486 117912 103514
rect 117688 102808 117740 102814
rect 117688 102750 117740 102756
rect 117424 93826 117636 93854
rect 117424 89714 117452 93826
rect 117424 89686 117636 89714
rect 117320 86964 117372 86970
rect 117320 86906 117372 86912
rect 117332 86873 117360 86906
rect 117318 86864 117374 86873
rect 117318 86799 117374 86808
rect 117320 84176 117372 84182
rect 117320 84118 117372 84124
rect 117332 83881 117360 84118
rect 117318 83872 117374 83881
rect 117318 83807 117374 83816
rect 117320 73160 117372 73166
rect 117320 73102 117372 73108
rect 117332 72729 117360 73102
rect 117318 72720 117374 72729
rect 117318 72655 117374 72664
rect 117320 67584 117372 67590
rect 117320 67526 117372 67532
rect 117332 67017 117360 67526
rect 117318 67008 117374 67017
rect 117318 66943 117374 66952
rect 117318 57624 117374 57633
rect 117318 57559 117374 57568
rect 117332 56234 117360 57559
rect 117320 56228 117372 56234
rect 117320 56170 117372 56176
rect 117318 51776 117374 51785
rect 117318 51711 117374 51720
rect 117332 46986 117360 51711
rect 117410 48920 117466 48929
rect 117410 48855 117466 48864
rect 117424 48346 117452 48855
rect 117412 48340 117464 48346
rect 117412 48282 117464 48288
rect 117320 46980 117372 46986
rect 117320 46922 117372 46928
rect 117318 45928 117374 45937
rect 117318 45863 117374 45872
rect 117332 45762 117360 45863
rect 117320 45756 117372 45762
rect 117320 45698 117372 45704
rect 117318 43072 117374 43081
rect 117318 43007 117374 43016
rect 117332 37330 117360 43007
rect 117320 37324 117372 37330
rect 117320 37266 117372 37272
rect 117226 37224 117282 37233
rect 117226 37159 117282 37168
rect 117240 34542 117268 37159
rect 117228 34536 117280 34542
rect 117228 34478 117280 34484
rect 117134 34368 117190 34377
rect 117134 34303 117190 34312
rect 117042 32328 117098 32337
rect 117042 32263 117098 32272
rect 116950 9616 117006 9625
rect 116950 9551 117006 9560
rect 117056 5302 117084 32263
rect 117148 5710 117176 34303
rect 117318 31512 117374 31521
rect 117318 31447 117374 31456
rect 117332 30394 117360 31447
rect 117320 30388 117372 30394
rect 117320 30330 117372 30336
rect 117502 16960 117558 16969
rect 117502 16895 117558 16904
rect 117516 16658 117544 16895
rect 117504 16652 117556 16658
rect 117504 16594 117556 16600
rect 117318 14104 117374 14113
rect 117318 14039 117374 14048
rect 117332 13870 117360 14039
rect 117320 13864 117372 13870
rect 117320 13806 117372 13812
rect 117318 11112 117374 11121
rect 117318 11047 117320 11056
rect 117372 11047 117374 11056
rect 117320 11018 117372 11024
rect 117318 8256 117374 8265
rect 117318 8191 117374 8200
rect 117332 7274 117360 8191
rect 117320 7268 117372 7274
rect 117320 7210 117372 7216
rect 117136 5704 117188 5710
rect 117136 5646 117188 5652
rect 117318 5400 117374 5409
rect 117318 5335 117374 5344
rect 117044 5296 117096 5302
rect 117044 5238 117096 5244
rect 117332 4214 117360 5335
rect 117320 4208 117372 4214
rect 117320 4150 117372 4156
rect 117608 3398 117636 89686
rect 117700 81433 117728 102750
rect 117884 101833 117912 103486
rect 117870 101824 117926 101833
rect 117870 101759 117926 101768
rect 117872 95192 117924 95198
rect 117872 95134 117924 95140
rect 117780 85060 117832 85066
rect 117780 85002 117832 85008
rect 117686 81424 117742 81433
rect 117686 81359 117742 81368
rect 117792 80054 117820 85002
rect 117700 80026 117820 80054
rect 117700 78577 117728 80026
rect 117686 78568 117742 78577
rect 117686 78503 117742 78512
rect 117884 69873 117912 95134
rect 117870 69864 117926 69873
rect 117870 69799 117926 69808
rect 117870 63336 117926 63345
rect 117870 63271 117926 63280
rect 117884 58886 117912 63271
rect 117872 58880 117924 58886
rect 117872 58822 117924 58828
rect 117870 40216 117926 40225
rect 117870 40151 117926 40160
rect 117884 34610 117912 40151
rect 117872 34604 117924 34610
rect 117872 34546 117924 34552
rect 117870 22808 117926 22817
rect 117870 22743 117926 22752
rect 117778 19816 117834 19825
rect 117778 19751 117834 19760
rect 117792 5642 117820 19751
rect 117884 5778 117912 22743
rect 117976 11762 118004 150447
rect 118054 138816 118110 138825
rect 118054 138751 118110 138760
rect 117964 11756 118016 11762
rect 117964 11698 118016 11704
rect 117872 5772 117924 5778
rect 117872 5714 117924 5720
rect 117780 5636 117832 5642
rect 117780 5578 117832 5584
rect 118068 3534 118096 138751
rect 118056 3528 118108 3534
rect 118056 3470 118108 3476
rect 117596 3392 117648 3398
rect 117596 3334 117648 3340
rect 118160 2145 118188 150719
rect 118252 127945 118280 152351
rect 119448 151814 119476 157354
rect 120368 157321 120396 159200
rect 120354 157312 120410 157321
rect 120354 157247 120410 157256
rect 120724 154760 120776 154766
rect 120724 154702 120776 154708
rect 120172 154624 120224 154630
rect 120172 154566 120224 154572
rect 120080 153536 120132 153542
rect 120080 153478 120132 153484
rect 120092 151994 120120 153478
rect 120184 153406 120212 154566
rect 120736 153882 120764 154702
rect 121288 154698 121316 159200
rect 121918 156632 121974 156641
rect 121918 156567 121974 156576
rect 121276 154692 121328 154698
rect 121276 154634 121328 154640
rect 120632 153876 120684 153882
rect 120632 153818 120684 153824
rect 120724 153876 120776 153882
rect 120724 153818 120776 153824
rect 120172 153400 120224 153406
rect 120172 153342 120224 153348
rect 120644 151994 120672 153818
rect 121460 152516 121512 152522
rect 121460 152458 121512 152464
rect 121472 151994 121500 152458
rect 121932 151994 121960 156567
rect 122300 154630 122328 159200
rect 123220 155530 123248 159200
rect 123852 156664 123904 156670
rect 123852 156606 123904 156612
rect 123220 155502 123340 155530
rect 122288 154624 122340 154630
rect 122288 154566 122340 154572
rect 123208 153332 123260 153338
rect 123208 153274 123260 153280
rect 122840 152720 122892 152726
rect 122840 152662 122892 152668
rect 122852 151994 122880 152662
rect 123220 151994 123248 153274
rect 123312 152522 123340 155502
rect 123300 152516 123352 152522
rect 123300 152458 123352 152464
rect 123864 151994 123892 156606
rect 124128 155100 124180 155106
rect 124128 155042 124180 155048
rect 124140 153338 124168 155042
rect 124128 153332 124180 153338
rect 124128 153274 124180 153280
rect 124232 152726 124260 159200
rect 125244 155378 125272 159200
rect 125232 155372 125284 155378
rect 125232 155314 125284 155320
rect 125138 155272 125194 155281
rect 125138 155207 125194 155216
rect 124220 152720 124272 152726
rect 124220 152662 124272 152668
rect 124496 152584 124548 152590
rect 124496 152526 124548 152532
rect 124508 151994 124536 152526
rect 125152 151994 125180 155207
rect 126164 154601 126192 159200
rect 127072 158704 127124 158710
rect 127072 158646 127124 158652
rect 126150 154592 126206 154601
rect 126150 154527 126206 154536
rect 125784 153876 125836 153882
rect 125784 153818 125836 153824
rect 125796 151994 125824 153818
rect 126428 152652 126480 152658
rect 126428 152594 126480 152600
rect 126440 151994 126468 152594
rect 127084 151994 127112 158646
rect 127176 152590 127204 159200
rect 128096 156126 128124 159200
rect 129108 157690 129136 159200
rect 129740 157820 129792 157826
rect 129740 157762 129792 157768
rect 129096 157684 129148 157690
rect 129096 157626 129148 157632
rect 128084 156120 128136 156126
rect 128084 156062 128136 156068
rect 129004 155984 129056 155990
rect 129004 155926 129056 155932
rect 128358 154320 128414 154329
rect 128358 154255 128414 154264
rect 127164 152584 127216 152590
rect 127164 152526 127216 152532
rect 128372 151994 128400 154255
rect 129016 151994 129044 155926
rect 129752 151994 129780 157762
rect 130120 155378 130148 159200
rect 131040 156670 131068 159200
rect 132052 157826 132080 159200
rect 132592 158296 132644 158302
rect 132592 158238 132644 158244
rect 132040 157820 132092 157826
rect 132040 157762 132092 157768
rect 131672 156732 131724 156738
rect 131672 156674 131724 156680
rect 131028 156664 131080 156670
rect 131028 156606 131080 156612
rect 131210 155408 131266 155417
rect 130108 155372 130160 155378
rect 131210 155343 131266 155352
rect 130108 155314 130160 155320
rect 131120 153944 131172 153950
rect 131120 153886 131172 153892
rect 130384 153876 130436 153882
rect 130384 153818 130436 153824
rect 130396 151994 130424 153818
rect 131132 151994 131160 153886
rect 131224 153882 131252 155343
rect 131302 154592 131358 154601
rect 131302 154527 131358 154536
rect 131316 153950 131344 154527
rect 131304 153944 131356 153950
rect 131304 153886 131356 153892
rect 131212 153876 131264 153882
rect 131212 153818 131264 153824
rect 131684 151994 131712 156674
rect 132604 151994 132632 158238
rect 132776 155508 132828 155514
rect 132776 155450 132828 155456
rect 132788 155417 132816 155450
rect 132972 155446 133000 159200
rect 133984 155514 134012 159200
rect 134892 158636 134944 158642
rect 134892 158578 134944 158584
rect 133972 155508 134024 155514
rect 133972 155450 134024 155456
rect 132960 155440 133012 155446
rect 132774 155408 132830 155417
rect 132960 155382 133012 155388
rect 132774 155343 132830 155352
rect 132960 155304 133012 155310
rect 132960 155246 133012 155252
rect 132972 154034 133000 155246
rect 132972 154006 133092 154034
rect 133064 153882 133092 154006
rect 133880 154012 133932 154018
rect 133880 153954 133932 153960
rect 132960 153876 133012 153882
rect 132960 153818 133012 153824
rect 133052 153876 133104 153882
rect 133052 153818 133104 153824
rect 132972 151994 133000 153818
rect 133892 151994 133920 153954
rect 134248 152652 134300 152658
rect 134248 152594 134300 152600
rect 134260 151994 134288 152594
rect 134904 151994 134932 158578
rect 134996 156738 135024 159200
rect 134984 156732 135036 156738
rect 134984 156674 135036 156680
rect 135168 155304 135220 155310
rect 135168 155246 135220 155252
rect 135180 154018 135208 155246
rect 135168 154012 135220 154018
rect 135168 153954 135220 153960
rect 135536 153876 135588 153882
rect 135536 153818 135588 153824
rect 135548 151994 135576 153818
rect 135916 152658 135944 159200
rect 136928 159174 137048 159200
rect 136822 156768 136878 156777
rect 136822 156703 136878 156712
rect 136548 155372 136600 155378
rect 136548 155314 136600 155320
rect 136180 154080 136232 154086
rect 136180 154022 136232 154028
rect 135904 152652 135956 152658
rect 135904 152594 135956 152600
rect 136192 151994 136220 154022
rect 136560 154018 136588 155314
rect 136548 154012 136600 154018
rect 136548 153954 136600 153960
rect 136836 151994 136864 156703
rect 137204 155718 137232 159310
rect 137834 159200 137890 160000
rect 138846 159200 138902 160000
rect 139858 159200 139914 160000
rect 140778 159200 140834 160000
rect 141790 159200 141846 160000
rect 142710 159200 142766 160000
rect 143722 159200 143778 160000
rect 144734 159200 144790 160000
rect 145654 159200 145710 160000
rect 146666 159200 146722 160000
rect 147586 159200 147642 160000
rect 148598 159200 148654 160000
rect 149610 159200 149666 160000
rect 150530 159200 150586 160000
rect 151542 159200 151598 160000
rect 152462 159200 152518 160000
rect 153474 159200 153530 160000
rect 154486 159200 154542 160000
rect 155406 159200 155462 160000
rect 156418 159202 156474 160000
rect 156524 159310 156736 159338
rect 156524 159202 156552 159310
rect 156418 159200 156552 159202
rect 137468 158772 137520 158778
rect 137468 158714 137520 158720
rect 137192 155712 137244 155718
rect 137192 155654 137244 155660
rect 137480 151994 137508 158714
rect 137848 154154 137876 159200
rect 138202 155408 138258 155417
rect 138202 155343 138258 155352
rect 137836 154148 137888 154154
rect 137836 154090 137888 154096
rect 138216 153950 138244 155343
rect 138860 155122 138888 159200
rect 139872 155514 139900 159200
rect 140136 158840 140188 158846
rect 140136 158782 140188 158788
rect 139860 155508 139912 155514
rect 139860 155450 139912 155456
rect 138860 155094 138980 155122
rect 138846 154456 138902 154465
rect 138846 154391 138902 154400
rect 138112 153944 138164 153950
rect 138112 153886 138164 153892
rect 138204 153944 138256 153950
rect 138204 153886 138256 153892
rect 138124 151994 138152 153886
rect 138860 151994 138888 154391
rect 138952 152794 138980 155094
rect 139492 152856 139544 152862
rect 139492 152798 139544 152804
rect 138940 152788 138992 152794
rect 138940 152730 138992 152736
rect 139504 151994 139532 152798
rect 140148 151994 140176 158782
rect 140792 155922 140820 159200
rect 140688 155916 140740 155922
rect 140688 155858 140740 155864
rect 140780 155916 140832 155922
rect 140780 155858 140832 155864
rect 140700 155802 140728 155858
rect 140700 155774 140912 155802
rect 140780 155576 140832 155582
rect 140780 155518 140832 155524
rect 140792 153950 140820 155518
rect 140884 154154 140912 155774
rect 141804 155582 141832 159200
rect 142252 156800 142304 156806
rect 142252 156742 142304 156748
rect 141792 155576 141844 155582
rect 141792 155518 141844 155524
rect 140872 154148 140924 154154
rect 140872 154090 140924 154096
rect 140964 154080 141016 154086
rect 140964 154022 141016 154028
rect 140688 153944 140740 153950
rect 140688 153886 140740 153892
rect 140780 153944 140832 153950
rect 140780 153886 140832 153892
rect 140700 153762 140728 153886
rect 140700 153734 140820 153762
rect 140792 152862 140820 153734
rect 140780 152856 140832 152862
rect 140780 152798 140832 152804
rect 140976 151994 141004 154022
rect 141424 152856 141476 152862
rect 141424 152798 141476 152804
rect 141436 151994 141464 152798
rect 142264 151994 142292 156742
rect 142724 152862 142752 159200
rect 142804 158908 142856 158914
rect 142804 158850 142856 158856
rect 142712 152856 142764 152862
rect 142712 152798 142764 152804
rect 142816 151994 142844 158850
rect 143736 155564 143764 159200
rect 144748 157758 144776 159200
rect 145288 158976 145340 158982
rect 145288 158918 145340 158924
rect 144736 157752 144788 157758
rect 144736 157694 144788 157700
rect 143816 155576 143868 155582
rect 143736 155536 143816 155564
rect 143816 155518 143868 155524
rect 143632 155440 143684 155446
rect 143632 155382 143684 155388
rect 143644 153950 143672 155382
rect 144828 155372 144880 155378
rect 144828 155314 144880 155320
rect 144840 154154 144868 155314
rect 144828 154148 144880 154154
rect 144828 154090 144880 154096
rect 144000 154012 144052 154018
rect 144000 153954 144052 153960
rect 143540 153944 143592 153950
rect 143540 153886 143592 153892
rect 143632 153944 143684 153950
rect 143632 153886 143684 153892
rect 143552 151994 143580 153886
rect 144012 151994 144040 153954
rect 144918 152552 144974 152561
rect 144918 152487 144974 152496
rect 144932 151994 144960 152487
rect 145300 151994 145328 158918
rect 145668 155514 145696 159200
rect 146680 156806 146708 159200
rect 146668 156800 146720 156806
rect 146668 156742 146720 156748
rect 147600 155514 147628 159200
rect 148612 157894 148640 159200
rect 148508 157888 148560 157894
rect 148508 157830 148560 157836
rect 148600 157888 148652 157894
rect 148600 157830 148652 157836
rect 145656 155508 145708 155514
rect 145656 155450 145708 155456
rect 147588 155508 147640 155514
rect 147588 155450 147640 155456
rect 146484 155372 146536 155378
rect 146484 155314 146536 155320
rect 145932 153264 145984 153270
rect 145932 153206 145984 153212
rect 145944 151994 145972 153206
rect 120092 151966 120336 151994
rect 120644 151966 120980 151994
rect 121472 151966 121624 151994
rect 121932 151966 122268 151994
rect 122852 151966 122912 151994
rect 123220 151966 123556 151994
rect 123864 151966 124200 151994
rect 124508 151966 124844 151994
rect 125152 151966 125488 151994
rect 125796 151966 126132 151994
rect 126440 151966 126776 151994
rect 127084 151966 127420 151994
rect 128372 151966 128708 151994
rect 129016 151966 129352 151994
rect 129752 151966 130088 151994
rect 130396 151966 130732 151994
rect 131132 151966 131376 151994
rect 131684 151966 132020 151994
rect 132604 151966 132664 151994
rect 132972 151966 133308 151994
rect 133892 151966 133952 151994
rect 134260 151966 134596 151994
rect 134904 151966 135240 151994
rect 135548 151966 135884 151994
rect 136192 151966 136528 151994
rect 136836 151966 137172 151994
rect 137480 151966 137816 151994
rect 138124 151966 138460 151994
rect 138860 151966 139196 151994
rect 139504 151966 139840 151994
rect 140148 151966 140484 151994
rect 140976 151966 141128 151994
rect 141436 151966 141772 151994
rect 142264 151966 142416 151994
rect 142816 151966 143060 151994
rect 143552 151966 143704 151994
rect 144012 151966 144348 151994
rect 144932 151966 144992 151994
rect 145300 151966 145636 151994
rect 145944 151966 146280 151994
rect 119356 151786 119476 151814
rect 119894 151872 119950 151881
rect 146496 151842 146524 155314
rect 146576 153944 146628 153950
rect 146576 153886 146628 153892
rect 146588 151994 146616 153886
rect 147956 152992 148008 152998
rect 147956 152934 148008 152940
rect 147220 152924 147272 152930
rect 147220 152866 147272 152872
rect 147232 151994 147260 152866
rect 147968 151994 147996 152934
rect 148520 151994 148548 157830
rect 149624 155922 149652 159200
rect 149612 155916 149664 155922
rect 149612 155858 149664 155864
rect 149060 155372 149112 155378
rect 149060 155314 149112 155320
rect 149072 153270 149100 155314
rect 149244 154012 149296 154018
rect 149244 153954 149296 153960
rect 149060 153264 149112 153270
rect 149060 153206 149112 153212
rect 149256 151994 149284 153954
rect 149888 153060 149940 153066
rect 149888 153002 149940 153008
rect 149900 151994 149928 153002
rect 150544 152930 150572 159200
rect 151176 157956 151228 157962
rect 151176 157898 151228 157904
rect 150624 156868 150676 156874
rect 150624 156810 150676 156816
rect 150532 152924 150584 152930
rect 150532 152866 150584 152872
rect 150636 151994 150664 156810
rect 151188 151994 151216 157898
rect 151556 155378 151584 159200
rect 151544 155372 151596 155378
rect 151544 155314 151596 155320
rect 152004 154148 152056 154154
rect 152004 154090 152056 154096
rect 152016 151994 152044 154090
rect 152476 153218 152504 159200
rect 153488 155786 153516 159200
rect 153752 158024 153804 158030
rect 153752 157966 153804 157972
rect 153476 155780 153528 155786
rect 153476 155722 153528 155728
rect 153108 155576 153160 155582
rect 153108 155518 153160 155524
rect 152476 153190 152596 153218
rect 152464 153128 152516 153134
rect 152464 153070 152516 153076
rect 152476 151994 152504 153070
rect 152568 152998 152596 153190
rect 153120 153066 153148 155518
rect 153108 153060 153160 153066
rect 153108 153002 153160 153008
rect 152556 152992 152608 152998
rect 152556 152934 152608 152940
rect 153198 152688 153254 152697
rect 153198 152623 153254 152632
rect 153212 151994 153240 152623
rect 153764 151994 153792 157966
rect 154500 156641 154528 159200
rect 154486 156632 154542 156641
rect 154486 156567 154542 156576
rect 155420 155990 155448 159200
rect 156432 159174 156552 159200
rect 156328 158364 156380 158370
rect 156328 158306 156380 158312
rect 155960 156936 156012 156942
rect 155960 156878 156012 156884
rect 155868 156052 155920 156058
rect 155868 155994 155920 156000
rect 155408 155984 155460 155990
rect 155408 155926 155460 155932
rect 155316 155576 155368 155582
rect 155316 155518 155368 155524
rect 155040 154284 155092 154290
rect 155040 154226 155092 154232
rect 154580 154080 154632 154086
rect 154580 154022 154632 154028
rect 154592 151994 154620 154022
rect 155052 151994 155080 154226
rect 155328 154086 155356 155518
rect 155880 154290 155908 155994
rect 155868 154284 155920 154290
rect 155868 154226 155920 154232
rect 155316 154080 155368 154086
rect 155316 154022 155368 154028
rect 155972 151994 156000 156878
rect 156340 151994 156368 158306
rect 156604 155984 156656 155990
rect 156604 155926 156656 155932
rect 156512 155644 156564 155650
rect 156512 155586 156564 155592
rect 156524 154222 156552 155586
rect 156616 155514 156644 155926
rect 156708 155514 156736 159310
rect 157338 159200 157394 160000
rect 158350 159200 158406 160000
rect 159270 159200 159326 160000
rect 160282 159200 160338 160000
rect 161294 159200 161350 160000
rect 162214 159200 162270 160000
rect 163226 159200 163282 160000
rect 164146 159200 164202 160000
rect 165158 159200 165214 160000
rect 166170 159200 166226 160000
rect 167090 159200 167146 160000
rect 168102 159200 168158 160000
rect 169022 159200 169078 160000
rect 170034 159200 170090 160000
rect 171046 159200 171102 160000
rect 171966 159200 172022 160000
rect 172978 159200 173034 160000
rect 173898 159200 173954 160000
rect 174910 159200 174966 160000
rect 175922 159200 175978 160000
rect 176842 159200 176898 160000
rect 177854 159200 177910 160000
rect 178774 159200 178830 160000
rect 179786 159200 179842 160000
rect 180798 159200 180854 160000
rect 181718 159200 181774 160000
rect 182730 159200 182786 160000
rect 183650 159200 183706 160000
rect 184662 159200 184718 160000
rect 185674 159200 185730 160000
rect 186594 159200 186650 160000
rect 187606 159200 187662 160000
rect 188526 159200 188582 160000
rect 189538 159200 189594 160000
rect 190550 159200 190606 160000
rect 191470 159200 191526 160000
rect 192482 159202 192538 160000
rect 192588 159310 192892 159338
rect 192588 159202 192616 159310
rect 192482 159200 192616 159202
rect 156604 155508 156656 155514
rect 156604 155450 156656 155456
rect 156696 155508 156748 155514
rect 156696 155450 156748 155456
rect 156512 154216 156564 154222
rect 156512 154158 156564 154164
rect 157352 154086 157380 159200
rect 158364 156874 158392 159200
rect 158996 158092 159048 158098
rect 158996 158034 159048 158040
rect 158352 156868 158404 156874
rect 158352 156810 158404 156816
rect 158720 156052 158772 156058
rect 158720 155994 158772 156000
rect 158732 155378 158760 155994
rect 158904 155916 158956 155922
rect 158904 155858 158956 155864
rect 158810 155544 158866 155553
rect 158810 155479 158866 155488
rect 158720 155372 158772 155378
rect 158720 155314 158772 155320
rect 156972 154080 157024 154086
rect 156972 154022 157024 154028
rect 157340 154080 157392 154086
rect 157340 154022 157392 154028
rect 156984 151994 157012 154022
rect 158824 153338 158852 155479
rect 157708 153332 157760 153338
rect 157708 153274 157760 153280
rect 158812 153332 158864 153338
rect 158812 153274 158864 153280
rect 157720 151994 157748 153274
rect 158916 153134 158944 155858
rect 158904 153128 158956 153134
rect 158904 153070 158956 153076
rect 158352 152448 158404 152454
rect 158352 152390 158404 152396
rect 158364 151994 158392 152390
rect 159008 151994 159036 158034
rect 159284 155786 159312 159200
rect 159272 155780 159324 155786
rect 159272 155722 159324 155728
rect 160098 155680 160154 155689
rect 160296 155650 160324 159200
rect 160926 156904 160982 156913
rect 160926 156839 160982 156848
rect 160098 155615 160154 155624
rect 160284 155644 160336 155650
rect 159640 154420 159692 154426
rect 159640 154362 159692 154368
rect 159652 151994 159680 154362
rect 160112 154154 160140 155615
rect 160284 155586 160336 155592
rect 160100 154148 160152 154154
rect 160100 154090 160152 154096
rect 160284 153196 160336 153202
rect 160284 153138 160336 153144
rect 160296 151994 160324 153138
rect 160940 151994 160968 156839
rect 161308 155281 161336 159200
rect 161664 158432 161716 158438
rect 161664 158374 161716 158380
rect 161294 155272 161350 155281
rect 161294 155207 161350 155216
rect 161676 151994 161704 158374
rect 162228 153490 162256 159200
rect 163240 155922 163268 159200
rect 164054 155952 164110 155961
rect 163228 155916 163280 155922
rect 164054 155887 164110 155896
rect 163228 155858 163280 155864
rect 162768 155576 162820 155582
rect 162768 155518 162820 155524
rect 162780 154290 162808 155518
rect 164068 154494 164096 155887
rect 164160 155582 164188 159200
rect 164240 158500 164292 158506
rect 164240 158442 164292 158448
rect 164148 155576 164200 155582
rect 164148 155518 164200 155524
rect 164056 154488 164108 154494
rect 164056 154430 164108 154436
rect 162860 154352 162912 154358
rect 162860 154294 162912 154300
rect 162768 154284 162820 154290
rect 162768 154226 162820 154232
rect 162228 153462 162348 153490
rect 162216 153332 162268 153338
rect 162216 153274 162268 153280
rect 162228 151994 162256 153274
rect 162320 153066 162348 153462
rect 162308 153060 162360 153066
rect 162308 153002 162360 153008
rect 162872 151994 162900 154294
rect 163502 152824 163558 152833
rect 163502 152759 163558 152768
rect 163516 151994 163544 152759
rect 164252 151994 164280 158442
rect 165172 154154 165200 159200
rect 166080 157072 166132 157078
rect 166080 157014 166132 157020
rect 165620 157004 165672 157010
rect 165620 156946 165672 156952
rect 164792 154148 164844 154154
rect 164792 154090 164844 154096
rect 165160 154148 165212 154154
rect 165160 154090 165212 154096
rect 164804 151994 164832 154090
rect 165632 151994 165660 156946
rect 166092 151994 166120 157014
rect 166184 156942 166212 159200
rect 166172 156936 166224 156942
rect 166172 156878 166224 156884
rect 167104 155038 167132 159200
rect 167276 158568 167328 158574
rect 167276 158510 167328 158516
rect 167000 155032 167052 155038
rect 167000 154974 167052 154980
rect 167092 155032 167144 155038
rect 167092 154974 167144 154980
rect 167012 154562 167040 154974
rect 167000 154556 167052 154562
rect 167000 154498 167052 154504
rect 146588 151966 146924 151994
rect 147232 151966 147568 151994
rect 147968 151966 148304 151994
rect 148520 151966 148948 151994
rect 149256 151966 149592 151994
rect 149900 151966 150236 151994
rect 150636 151966 150880 151994
rect 151188 151966 151524 151994
rect 152016 151966 152168 151994
rect 152476 151966 152812 151994
rect 153212 151966 153456 151994
rect 153764 151966 154100 151994
rect 154592 151966 154744 151994
rect 155052 151966 155388 151994
rect 155972 151966 156032 151994
rect 156340 151966 156676 151994
rect 156984 151966 157320 151994
rect 157720 151966 158056 151994
rect 158364 151966 158700 151994
rect 159008 151966 159344 151994
rect 159652 151966 159988 151994
rect 160296 151966 160632 151994
rect 160940 151966 161276 151994
rect 161676 151966 161920 151994
rect 162228 151966 162564 151994
rect 162872 151966 163208 151994
rect 163516 151966 163852 151994
rect 164252 151966 164496 151994
rect 164804 151966 165140 151994
rect 165632 151966 165784 151994
rect 166092 151966 166428 151994
rect 167288 151858 167316 158510
rect 168116 157010 168144 159200
rect 168104 157004 168156 157010
rect 168104 156946 168156 156952
rect 167460 154352 167512 154358
rect 167460 154294 167512 154300
rect 167472 151994 167500 154294
rect 169036 154154 169064 159200
rect 169760 157072 169812 157078
rect 169760 157014 169812 157020
rect 169772 155786 169800 157014
rect 169760 155780 169812 155786
rect 169760 155722 169812 155728
rect 169760 154896 169812 154902
rect 169760 154838 169812 154844
rect 169772 154358 169800 154838
rect 169760 154352 169812 154358
rect 169760 154294 169812 154300
rect 170048 154306 170076 159200
rect 170680 157140 170732 157146
rect 170680 157082 170732 157088
rect 170048 154278 170168 154306
rect 170036 154216 170088 154222
rect 170036 154158 170088 154164
rect 169024 154148 169076 154154
rect 169024 154090 169076 154096
rect 169392 153264 169444 153270
rect 169392 153206 169444 153212
rect 168380 152380 168432 152386
rect 168380 152322 168432 152328
rect 168392 151994 168420 152322
rect 169070 152244 169122 152250
rect 169070 152186 169122 152192
rect 167472 151966 167808 151994
rect 168392 151966 168452 151994
rect 169082 151980 169110 152186
rect 169404 151994 169432 153206
rect 170048 151994 170076 154158
rect 170140 153202 170168 154278
rect 170128 153196 170180 153202
rect 170128 153138 170180 153144
rect 170692 151994 170720 157082
rect 171060 156074 171088 159200
rect 171416 157208 171468 157214
rect 171416 157150 171468 157156
rect 171060 156046 171272 156074
rect 171244 155038 171272 156046
rect 171232 155032 171284 155038
rect 171232 154974 171284 154980
rect 171140 153264 171192 153270
rect 171140 153206 171192 153212
rect 169404 151966 169740 151994
rect 170048 151966 170384 151994
rect 170692 151966 171028 151994
rect 119894 151807 119950 151816
rect 146484 151836 146536 151842
rect 118332 151564 118384 151570
rect 118332 151506 118384 151512
rect 118238 127936 118294 127945
rect 118238 127871 118294 127880
rect 118238 121408 118294 121417
rect 118238 121343 118294 121352
rect 118252 4350 118280 121343
rect 118344 118697 118372 151506
rect 118424 151428 118476 151434
rect 118424 151370 118476 151376
rect 118330 118688 118386 118697
rect 118330 118623 118386 118632
rect 118436 115841 118464 151370
rect 118608 150748 118660 150754
rect 118608 150690 118660 150696
rect 118514 149968 118570 149977
rect 118514 149903 118570 149912
rect 118422 115832 118478 115841
rect 118422 115767 118478 115776
rect 118422 112704 118478 112713
rect 118422 112639 118478 112648
rect 118332 11756 118384 11762
rect 118332 11698 118384 11704
rect 118240 4344 118292 4350
rect 118240 4286 118292 4292
rect 118146 2136 118202 2145
rect 118146 2071 118202 2080
rect 118344 1873 118372 11698
rect 118436 4486 118464 112639
rect 118528 89729 118556 149903
rect 118620 92449 118648 150690
rect 118698 106856 118754 106865
rect 118698 106791 118754 106800
rect 118606 92440 118662 92449
rect 118606 92375 118662 92384
rect 118514 89720 118570 89729
rect 118514 89655 118570 89664
rect 118608 88868 118660 88874
rect 118608 88810 118660 88816
rect 118620 75721 118648 88810
rect 118606 75712 118662 75721
rect 118606 75647 118662 75656
rect 118606 60480 118662 60489
rect 118606 60415 118662 60424
rect 118514 54632 118570 54641
rect 118514 54567 118570 54576
rect 118528 39506 118556 54567
rect 118620 53854 118648 60415
rect 118608 53848 118660 53854
rect 118608 53790 118660 53796
rect 118516 39500 118568 39506
rect 118516 39442 118568 39448
rect 118514 28520 118570 28529
rect 118514 28455 118570 28464
rect 118528 5846 118556 28455
rect 118606 25664 118662 25673
rect 118606 25599 118662 25608
rect 118620 5914 118648 25599
rect 118608 5908 118660 5914
rect 118608 5850 118660 5856
rect 118516 5840 118568 5846
rect 118516 5782 118568 5788
rect 118712 4962 118740 106791
rect 118700 4956 118752 4962
rect 118700 4898 118752 4904
rect 118424 4480 118476 4486
rect 118424 4422 118476 4428
rect 119356 2718 119384 151786
rect 119618 151192 119674 151201
rect 119618 151127 119674 151136
rect 119434 150920 119490 150929
rect 119434 150855 119490 150864
rect 119344 2712 119396 2718
rect 119344 2654 119396 2660
rect 119448 2281 119476 150855
rect 119528 150612 119580 150618
rect 119528 150554 119580 150560
rect 119434 2272 119490 2281
rect 119434 2207 119490 2216
rect 119540 2174 119568 150554
rect 119632 2689 119660 151127
rect 119802 151056 119858 151065
rect 119802 150991 119858 151000
rect 119712 99476 119764 99482
rect 119712 99418 119764 99424
rect 119724 4026 119752 99418
rect 119816 4706 119844 150991
rect 119908 67454 119936 151807
rect 167164 151830 167316 151858
rect 146484 151778 146536 151784
rect 127716 151768 127768 151774
rect 127768 151716 128064 151722
rect 127716 151710 128064 151716
rect 127728 151694 128064 151710
rect 171152 151706 171180 153206
rect 171428 151994 171456 157150
rect 171980 155417 172008 159200
rect 172992 155718 173020 159200
rect 173912 157214 173940 159200
rect 174544 157344 174596 157350
rect 174544 157286 174596 157292
rect 173900 157208 173952 157214
rect 173900 157150 173952 157156
rect 173808 157140 173860 157146
rect 173808 157082 173860 157088
rect 173820 155786 173848 157082
rect 173898 157040 173954 157049
rect 173898 156975 173954 156984
rect 173808 155780 173860 155786
rect 173808 155722 173860 155728
rect 172980 155712 173032 155718
rect 172980 155654 173032 155660
rect 171966 155408 172022 155417
rect 171966 155343 172022 155352
rect 172612 154488 172664 154494
rect 172612 154430 172664 154436
rect 171968 153468 172020 153474
rect 171968 153410 172020 153416
rect 171980 151994 172008 153410
rect 172624 151994 172652 154430
rect 173256 152312 173308 152318
rect 173256 152254 173308 152260
rect 173268 151994 173296 152254
rect 173912 151994 173940 156975
rect 174556 151994 174584 157286
rect 174924 154601 174952 159200
rect 175740 156596 175792 156602
rect 175740 156538 175792 156544
rect 174910 154592 174966 154601
rect 174910 154527 174966 154536
rect 175280 153808 175332 153814
rect 175280 153750 175332 153756
rect 175292 151994 175320 153750
rect 175752 151994 175780 156538
rect 175936 155786 175964 159200
rect 175924 155780 175976 155786
rect 175924 155722 175976 155728
rect 176856 154902 176884 159200
rect 177868 157146 177896 159200
rect 177856 157140 177908 157146
rect 177856 157082 177908 157088
rect 178130 155816 178186 155825
rect 178130 155751 178186 155760
rect 175832 154896 175884 154902
rect 175832 154838 175884 154844
rect 176844 154896 176896 154902
rect 176844 154838 176896 154844
rect 177948 154896 178000 154902
rect 177948 154838 178000 154844
rect 175844 152250 175872 154838
rect 175922 154728 175978 154737
rect 175922 154663 175978 154672
rect 175936 154494 175964 154663
rect 175924 154488 175976 154494
rect 175924 154430 175976 154436
rect 177960 154290 177988 154838
rect 178040 154760 178092 154766
rect 178040 154702 178092 154708
rect 177212 154284 177264 154290
rect 177212 154226 177264 154232
rect 177948 154284 178000 154290
rect 177948 154226 178000 154232
rect 175832 152244 175884 152250
rect 175832 152186 175884 152192
rect 176890 152176 176942 152182
rect 176890 152118 176942 152124
rect 171428 151966 171672 151994
rect 171980 151966 172316 151994
rect 172624 151966 172960 151994
rect 173268 151966 173604 151994
rect 173912 151966 174248 151994
rect 174556 151966 174892 151994
rect 175292 151966 175536 151994
rect 175752 151966 176272 151994
rect 176902 151980 176930 152118
rect 177224 151994 177252 154226
rect 178052 153678 178080 154702
rect 178040 153672 178092 153678
rect 178040 153614 178092 153620
rect 178144 151994 178172 155751
rect 178788 154766 178816 159200
rect 179420 155916 179472 155922
rect 179420 155858 179472 155864
rect 178776 154760 178828 154766
rect 178776 154702 178828 154708
rect 178222 154592 178278 154601
rect 178222 154527 178278 154536
rect 178236 152250 178264 154527
rect 179432 153814 179460 155858
rect 179510 154864 179566 154873
rect 179510 154799 179566 154808
rect 179420 153808 179472 153814
rect 179420 153750 179472 153756
rect 179524 153406 179552 154799
rect 179420 153400 179472 153406
rect 179420 153342 179472 153348
rect 179512 153400 179564 153406
rect 179512 153342 179564 153348
rect 178224 152244 178276 152250
rect 178224 152186 178276 152192
rect 178822 152108 178874 152114
rect 178822 152050 178874 152056
rect 177224 151966 177560 151994
rect 178144 151966 178204 151994
rect 178834 151980 178862 152050
rect 179432 151994 179460 153342
rect 179800 152386 179828 159200
rect 179880 158160 179932 158166
rect 179880 158102 179932 158108
rect 179788 152380 179840 152386
rect 179788 152322 179840 152328
rect 179892 151994 179920 158102
rect 180812 155922 180840 159200
rect 181076 157276 181128 157282
rect 181076 157218 181128 157224
rect 180800 155916 180852 155922
rect 180800 155858 180852 155864
rect 180432 153740 180484 153746
rect 180432 153682 180484 153688
rect 180444 151994 180472 153682
rect 181088 151994 181116 157218
rect 181732 153626 181760 159200
rect 182088 156460 182140 156466
rect 182088 156402 182140 156408
rect 182100 155038 182128 156402
rect 182088 155032 182140 155038
rect 182088 154974 182140 154980
rect 182744 154698 182772 159200
rect 182088 154692 182140 154698
rect 182088 154634 182140 154640
rect 182732 154692 182784 154698
rect 182732 154634 182784 154640
rect 181732 153598 181852 153626
rect 181720 153468 181772 153474
rect 181720 153410 181772 153416
rect 181732 151994 181760 153410
rect 181824 152318 181852 153598
rect 182100 153474 182128 154634
rect 183664 154630 183692 159200
rect 183652 154624 183704 154630
rect 183652 154566 183704 154572
rect 183008 154556 183060 154562
rect 183008 154498 183060 154504
rect 182088 153468 182140 153474
rect 182088 153410 182140 153416
rect 182362 152960 182418 152969
rect 182362 152895 182418 152904
rect 181812 152312 181864 152318
rect 181812 152254 181864 152260
rect 182376 151994 182404 152895
rect 183020 151994 183048 154498
rect 184676 154426 184704 159200
rect 185584 155168 185636 155174
rect 185584 155110 185636 155116
rect 184296 154420 184348 154426
rect 184296 154362 184348 154368
rect 184664 154420 184716 154426
rect 184664 154362 184716 154368
rect 183652 152040 183704 152046
rect 179432 151966 179492 151994
rect 179892 151966 180136 151994
rect 180444 151966 180780 151994
rect 181088 151966 181424 151994
rect 181732 151966 182068 151994
rect 182376 151966 182712 151994
rect 183020 151966 183356 151994
rect 184308 151994 184336 154362
rect 184940 154352 184992 154358
rect 184940 154294 184992 154300
rect 184952 151994 184980 154294
rect 185596 153746 185624 155110
rect 185584 153740 185636 153746
rect 185688 153728 185716 159200
rect 186412 156528 186464 156534
rect 186412 156470 186464 156476
rect 186320 156460 186372 156466
rect 186320 156402 186372 156408
rect 186332 154766 186360 156402
rect 186320 154760 186372 154766
rect 186320 154702 186372 154708
rect 185688 153700 185808 153728
rect 185584 153682 185636 153688
rect 185676 153604 185728 153610
rect 185676 153546 185728 153552
rect 185688 151994 185716 153546
rect 185780 152182 185808 153700
rect 185768 152176 185820 152182
rect 185768 152118 185820 152124
rect 186424 151994 186452 156470
rect 186608 155922 186636 159200
rect 186964 157480 187016 157486
rect 186964 157422 187016 157428
rect 186596 155916 186648 155922
rect 186596 155858 186648 155864
rect 186976 151994 187004 157422
rect 187620 155038 187648 159200
rect 187698 157176 187754 157185
rect 187698 157111 187754 157120
rect 187608 155032 187660 155038
rect 187608 154974 187660 154980
rect 187712 151994 187740 157111
rect 188540 154426 188568 159200
rect 189552 157214 189580 159200
rect 189632 158228 189684 158234
rect 189632 158170 189684 158176
rect 189080 157208 189132 157214
rect 189080 157150 189132 157156
rect 189540 157208 189592 157214
rect 189540 157150 189592 157156
rect 188528 154420 188580 154426
rect 188528 154362 188580 154368
rect 188252 153400 188304 153406
rect 188252 153342 188304 153348
rect 188264 151994 188292 153342
rect 189092 151994 189120 157150
rect 189644 151994 189672 158170
rect 190460 157344 190512 157350
rect 190460 157286 190512 157292
rect 190472 151994 190500 157286
rect 190564 155922 190592 159200
rect 190552 155916 190604 155922
rect 190552 155858 190604 155864
rect 190826 155136 190882 155145
rect 190826 155071 190882 155080
rect 190840 151994 190868 155071
rect 191484 154698 191512 159200
rect 192496 159174 192616 159200
rect 192116 157548 192168 157554
rect 192116 157490 192168 157496
rect 191564 157276 191616 157282
rect 191564 157218 191616 157224
rect 191472 154692 191524 154698
rect 191472 154634 191524 154640
rect 191576 151994 191604 157218
rect 192128 151994 192156 157490
rect 192864 154494 192892 159310
rect 193402 159200 193458 160000
rect 194414 159200 194470 160000
rect 195334 159200 195390 160000
rect 196346 159200 196402 160000
rect 197358 159200 197414 160000
rect 198278 159200 198334 160000
rect 199290 159200 199346 160000
rect 200210 159200 200266 160000
rect 201222 159200 201278 160000
rect 202234 159200 202290 160000
rect 203154 159200 203210 160000
rect 204166 159200 204222 160000
rect 205086 159200 205142 160000
rect 206098 159200 206154 160000
rect 207110 159200 207166 160000
rect 208030 159200 208086 160000
rect 209042 159200 209098 160000
rect 209962 159200 210018 160000
rect 210974 159200 211030 160000
rect 211986 159200 212042 160000
rect 212906 159200 212962 160000
rect 213918 159200 213974 160000
rect 214838 159200 214894 160000
rect 215850 159200 215906 160000
rect 216862 159200 216918 160000
rect 217782 159200 217838 160000
rect 218794 159200 218850 160000
rect 219714 159200 219770 160000
rect 220726 159200 220782 160000
rect 221738 159200 221794 160000
rect 222658 159200 222714 160000
rect 223670 159200 223726 160000
rect 224590 159200 224646 160000
rect 225602 159200 225658 160000
rect 226614 159200 226670 160000
rect 227534 159200 227590 160000
rect 228546 159200 228602 160000
rect 229466 159200 229522 160000
rect 230478 159200 230534 160000
rect 231490 159200 231546 160000
rect 232410 159200 232466 160000
rect 233422 159200 233478 160000
rect 234342 159200 234398 160000
rect 235354 159200 235410 160000
rect 236274 159200 236330 160000
rect 237286 159200 237342 160000
rect 238298 159200 238354 160000
rect 239218 159200 239274 160000
rect 240230 159200 240286 160000
rect 241150 159200 241206 160000
rect 242162 159200 242218 160000
rect 243174 159200 243230 160000
rect 244094 159200 244150 160000
rect 245106 159200 245162 160000
rect 246026 159200 246082 160000
rect 247038 159200 247094 160000
rect 248050 159200 248106 160000
rect 248970 159200 249026 160000
rect 249982 159200 250038 160000
rect 250902 159200 250958 160000
rect 251914 159200 251970 160000
rect 252926 159200 252982 160000
rect 253846 159200 253902 160000
rect 254858 159200 254914 160000
rect 255778 159200 255834 160000
rect 256790 159200 256846 160000
rect 257802 159200 257858 160000
rect 258722 159200 258778 160000
rect 259734 159200 259790 160000
rect 260654 159200 260710 160000
rect 261666 159200 261722 160000
rect 262678 159200 262734 160000
rect 263598 159200 263654 160000
rect 264610 159200 264666 160000
rect 265530 159200 265586 160000
rect 266542 159200 266598 160000
rect 267554 159200 267610 160000
rect 268474 159200 268530 160000
rect 269486 159200 269542 160000
rect 270406 159200 270462 160000
rect 271418 159200 271474 160000
rect 272338 159202 272394 160000
rect 272444 159310 272840 159338
rect 272444 159202 272472 159310
rect 272338 159200 272472 159202
rect 193416 157282 193444 159200
rect 193404 157276 193456 157282
rect 193404 157218 193456 157224
rect 194428 154902 194456 159200
rect 194968 156188 195020 156194
rect 194968 156130 195020 156136
rect 194232 154896 194284 154902
rect 194230 154864 194232 154873
rect 194416 154896 194468 154902
rect 194284 154864 194286 154873
rect 193128 154828 193180 154834
rect 194416 154838 194468 154844
rect 194230 154799 194286 154808
rect 193128 154770 193180 154776
rect 192760 154488 192812 154494
rect 192760 154430 192812 154436
rect 192852 154488 192904 154494
rect 192852 154430 192904 154436
rect 192772 151994 192800 154430
rect 193140 153610 193168 154770
rect 194980 154766 195008 156130
rect 195348 154766 195376 159200
rect 196070 155000 196126 155009
rect 196070 154935 196126 154944
rect 195520 154828 195572 154834
rect 195520 154770 195572 154776
rect 194968 154760 195020 154766
rect 194968 154702 195020 154708
rect 195336 154760 195388 154766
rect 195336 154702 195388 154708
rect 195532 153678 195560 154770
rect 195428 153672 195480 153678
rect 195428 153614 195480 153620
rect 195520 153672 195572 153678
rect 195520 153614 195572 153620
rect 193128 153604 193180 153610
rect 193128 153546 193180 153552
rect 193404 153536 193456 153542
rect 193404 153478 193456 153484
rect 193416 151994 193444 153478
rect 194784 153332 194836 153338
rect 194784 153274 194836 153280
rect 194796 151994 194824 153274
rect 195440 151994 195468 153614
rect 196084 151994 196112 154935
rect 196360 154630 196388 159200
rect 197372 156618 197400 159200
rect 198004 157616 198056 157622
rect 198004 157558 198056 157564
rect 197372 156590 197492 156618
rect 196716 156528 196768 156534
rect 196716 156470 196768 156476
rect 197360 156528 197412 156534
rect 197360 156470 197412 156476
rect 196348 154624 196400 154630
rect 196348 154566 196400 154572
rect 196728 151994 196756 156470
rect 197372 155922 197400 156470
rect 197360 155916 197412 155922
rect 197360 155858 197412 155864
rect 197268 153332 197320 153338
rect 197268 153274 197320 153280
rect 183704 151988 184000 151994
rect 183652 151982 184000 151988
rect 183664 151966 184000 151982
rect 184308 151966 184644 151994
rect 184952 151966 185288 151994
rect 185688 151966 186024 151994
rect 186424 151966 186668 151994
rect 186976 151966 187312 151994
rect 187712 151966 187956 151994
rect 188264 151966 188600 151994
rect 189092 151966 189244 151994
rect 189644 151966 189888 151994
rect 190472 151966 190532 151994
rect 190840 151966 191176 151994
rect 191576 151966 191820 151994
rect 192128 151966 192464 151994
rect 192772 151966 193108 151994
rect 193416 151966 193752 151994
rect 194060 151978 194396 151994
rect 194048 151972 194396 151978
rect 194100 151966 194396 151972
rect 194796 151966 195132 151994
rect 195440 151966 195776 151994
rect 196084 151966 196420 151994
rect 196728 151966 197064 151994
rect 194048 151914 194100 151920
rect 171140 151700 171192 151706
rect 171140 151642 171192 151648
rect 197280 151638 197308 153274
rect 197464 152046 197492 156590
rect 197452 152040 197504 152046
rect 197452 151982 197504 151988
rect 198016 151994 198044 157558
rect 198292 154698 198320 159200
rect 199106 154864 199162 154873
rect 199106 154799 199162 154808
rect 198280 154692 198332 154698
rect 198280 154634 198332 154640
rect 198740 153468 198792 153474
rect 198740 153410 198792 153416
rect 198752 151994 198780 153410
rect 198016 151966 198352 151994
rect 198752 151966 198996 151994
rect 199120 151910 199148 154799
rect 199304 154766 199332 159200
rect 199384 156392 199436 156398
rect 199384 156334 199436 156340
rect 199292 154760 199344 154766
rect 199292 154702 199344 154708
rect 199396 151994 199424 156334
rect 200224 155854 200252 159200
rect 201236 157350 201264 159200
rect 201224 157344 201276 157350
rect 200394 157312 200450 157321
rect 201224 157286 201276 157292
rect 200394 157247 200450 157256
rect 200028 155848 200080 155854
rect 200212 155848 200264 155854
rect 200080 155796 200160 155802
rect 200028 155790 200160 155796
rect 200212 155790 200264 155796
rect 200040 155774 200160 155790
rect 200132 153542 200160 155774
rect 200120 153536 200172 153542
rect 200120 153478 200172 153484
rect 199396 151966 199640 151994
rect 197360 151904 197412 151910
rect 199108 151904 199160 151910
rect 197412 151852 197708 151858
rect 197360 151846 197708 151852
rect 200408 151858 200436 157247
rect 201958 155952 202014 155961
rect 201958 155887 201960 155896
rect 202012 155887 202014 155896
rect 201960 155858 202012 155864
rect 202248 155242 202276 159200
rect 202788 155848 202840 155854
rect 202788 155790 202840 155796
rect 202236 155236 202288 155242
rect 202236 155178 202288 155184
rect 202800 154562 202828 155790
rect 203168 155310 203196 159200
rect 203246 155952 203302 155961
rect 203246 155887 203302 155896
rect 203156 155304 203208 155310
rect 203156 155246 203208 155252
rect 202880 155100 202932 155106
rect 202932 155060 203104 155088
rect 202880 155042 202932 155048
rect 201500 154556 201552 154562
rect 201500 154498 201552 154504
rect 202788 154556 202840 154562
rect 202788 154498 202840 154504
rect 200580 153536 200632 153542
rect 200580 153478 200632 153484
rect 200592 151994 200620 153478
rect 201512 151994 201540 154498
rect 201868 152516 201920 152522
rect 201868 152458 201920 152464
rect 201880 151994 201908 152458
rect 203076 151994 203104 155060
rect 203260 152522 203288 155887
rect 204180 153882 204208 159200
rect 205100 156534 205128 159200
rect 205824 157684 205876 157690
rect 205824 157626 205876 157632
rect 205088 156528 205140 156534
rect 205088 156470 205140 156476
rect 204812 156120 204864 156126
rect 204812 156062 204864 156068
rect 203892 153876 203944 153882
rect 203892 153818 203944 153824
rect 204168 153876 204220 153882
rect 204168 153818 204220 153824
rect 203248 152516 203300 152522
rect 203248 152458 203300 152464
rect 203904 151994 203932 153818
rect 204536 152584 204588 152590
rect 204536 152526 204588 152532
rect 204548 151994 204576 152526
rect 204824 152130 204852 156062
rect 204824 152102 205128 152130
rect 205100 151994 205128 152102
rect 205836 151994 205864 157626
rect 206112 154698 206140 159200
rect 207124 156670 207152 159200
rect 207756 157820 207808 157826
rect 207756 157762 207808 157768
rect 207020 156664 207072 156670
rect 207020 156606 207072 156612
rect 207112 156664 207164 156670
rect 207112 156606 207164 156612
rect 206468 155440 206520 155446
rect 206468 155382 206520 155388
rect 206100 154692 206152 154698
rect 206100 154634 206152 154640
rect 206480 151994 206508 155382
rect 207032 151994 207060 156606
rect 207768 151994 207796 157762
rect 208044 152522 208072 159200
rect 208492 155848 208544 155854
rect 208492 155790 208544 155796
rect 208504 153610 208532 155790
rect 209056 155394 209084 159200
rect 209872 156460 209924 156466
rect 209872 156402 209924 156408
rect 209056 155366 209176 155394
rect 209044 155236 209096 155242
rect 209044 155178 209096 155184
rect 208400 153604 208452 153610
rect 208400 153546 208452 153552
rect 208492 153604 208544 153610
rect 208492 153546 208544 153552
rect 208032 152516 208084 152522
rect 208032 152458 208084 152464
rect 208412 151994 208440 153546
rect 209056 151994 209084 155178
rect 209148 152726 209176 155366
rect 209136 152720 209188 152726
rect 209136 152662 209188 152668
rect 209884 151994 209912 156402
rect 209976 155106 210004 159200
rect 210988 155242 211016 159200
rect 212000 155446 212028 159200
rect 212920 156738 212948 159200
rect 212908 156732 212960 156738
rect 212908 156674 212960 156680
rect 211896 155440 211948 155446
rect 211896 155382 211948 155388
rect 211988 155440 212040 155446
rect 211988 155382 212040 155388
rect 210976 155236 211028 155242
rect 210976 155178 211028 155184
rect 209964 155100 210016 155106
rect 209964 155042 210016 155048
rect 211620 153944 211672 153950
rect 211620 153886 211672 153892
rect 211160 153808 211212 153814
rect 211160 153750 211212 153756
rect 210332 152652 210384 152658
rect 210332 152594 210384 152600
rect 210344 151994 210372 152594
rect 211172 151994 211200 153750
rect 211632 151994 211660 153886
rect 211908 152658 211936 155382
rect 213932 154630 213960 159200
rect 214852 155553 214880 159200
rect 214838 155544 214894 155553
rect 214838 155479 214894 155488
rect 213920 154624 213972 154630
rect 213920 154566 213972 154572
rect 215864 153950 215892 159200
rect 216220 157752 216272 157758
rect 216220 157694 216272 157700
rect 215852 153944 215904 153950
rect 215852 153886 215904 153892
rect 213920 153740 213972 153746
rect 213920 153682 213972 153688
rect 212540 152788 212592 152794
rect 212540 152730 212592 152736
rect 211896 152652 211948 152658
rect 211896 152594 211948 152600
rect 212448 152652 212500 152658
rect 212448 152594 212500 152600
rect 200592 151966 200928 151994
rect 201512 151966 201572 151994
rect 201880 151966 202216 151994
rect 202524 151978 202860 151994
rect 202512 151972 202860 151978
rect 202564 151966 202860 151972
rect 203076 151966 203504 151994
rect 203904 151966 204240 151994
rect 204548 151966 204884 151994
rect 205100 151966 205528 151994
rect 205836 151966 206172 151994
rect 206480 151966 206816 151994
rect 207032 151966 207460 151994
rect 207768 151966 208104 151994
rect 208412 151966 208748 151994
rect 209056 151966 209392 151994
rect 209884 151966 210036 151994
rect 210344 151966 210680 151994
rect 211172 151966 211324 151994
rect 211632 151966 211968 151994
rect 202512 151914 202564 151920
rect 199108 151846 199160 151852
rect 197372 151830 197708 151846
rect 200284 151830 200436 151858
rect 212460 151842 212488 152594
rect 212552 151994 212580 152730
rect 213932 151994 213960 153682
rect 214288 153604 214340 153610
rect 214288 153546 214340 153552
rect 214300 151994 214328 153546
rect 214932 152856 214984 152862
rect 214932 152798 214984 152804
rect 214944 151994 214972 152798
rect 215576 152448 215628 152454
rect 215576 152390 215628 152396
rect 215588 151994 215616 152390
rect 216232 151994 216260 157694
rect 216876 154612 216904 159200
rect 217508 156460 217560 156466
rect 217508 156402 217560 156408
rect 216876 154584 216996 154612
rect 216864 154012 216916 154018
rect 216864 153954 216916 153960
rect 216876 151994 216904 153954
rect 216968 152658 216996 154584
rect 216956 152652 217008 152658
rect 216956 152594 217008 152600
rect 217520 151994 217548 156402
rect 217796 155446 217824 159200
rect 218152 156052 218204 156058
rect 218152 155994 218204 156000
rect 217784 155440 217836 155446
rect 217784 155382 217836 155388
rect 218164 151994 218192 155994
rect 218808 155689 218836 159200
rect 218888 157888 218940 157894
rect 218888 157830 218940 157836
rect 218794 155680 218850 155689
rect 218794 155615 218850 155624
rect 218900 151994 218928 157830
rect 219624 154692 219676 154698
rect 219624 154634 219676 154640
rect 219256 154624 219308 154630
rect 219254 154592 219256 154601
rect 219636 154601 219664 154634
rect 219308 154592 219310 154601
rect 219254 154527 219310 154536
rect 219622 154592 219678 154601
rect 219622 154527 219678 154536
rect 219728 154018 219756 159200
rect 220636 156052 220688 156058
rect 220636 155994 220688 156000
rect 220648 155310 220676 155994
rect 220636 155304 220688 155310
rect 220636 155246 220688 155252
rect 219716 154012 219768 154018
rect 219716 153954 219768 153960
rect 219624 153672 219676 153678
rect 219624 153614 219676 153620
rect 219636 151994 219664 153614
rect 220084 152924 220136 152930
rect 220084 152866 220136 152872
rect 220096 151994 220124 152866
rect 220740 152590 220768 159200
rect 220820 155984 220872 155990
rect 220820 155926 220872 155932
rect 220728 152584 220780 152590
rect 220728 152526 220780 152532
rect 220832 151994 220860 155926
rect 221752 155514 221780 159200
rect 222108 155984 222160 155990
rect 222108 155926 222160 155932
rect 221740 155508 221792 155514
rect 221740 155450 221792 155456
rect 222120 155446 222148 155926
rect 222108 155440 222160 155446
rect 222108 155382 222160 155388
rect 222672 154630 222700 159200
rect 222750 156632 222806 156641
rect 222750 156567 222806 156576
rect 222108 154624 222160 154630
rect 222108 154566 222160 154572
rect 222660 154624 222712 154630
rect 222660 154566 222712 154572
rect 222120 153218 222148 154566
rect 222120 153190 222240 153218
rect 221372 152992 221424 152998
rect 221372 152934 221424 152940
rect 221384 151994 221412 152934
rect 222212 151994 222240 153190
rect 222764 151994 222792 156567
rect 223684 155310 223712 159200
rect 224040 155644 224092 155650
rect 224040 155586 224092 155592
rect 223672 155304 223724 155310
rect 223672 155246 223724 155252
rect 223580 153128 223632 153134
rect 223580 153070 223632 153076
rect 223592 151994 223620 153070
rect 224052 151994 224080 155586
rect 224604 152794 224632 159200
rect 225328 156868 225380 156874
rect 225328 156810 225380 156816
rect 224960 154080 225012 154086
rect 224960 154022 225012 154028
rect 224592 152788 224644 152794
rect 224592 152730 224644 152736
rect 224972 151994 225000 154022
rect 225340 151994 225368 156810
rect 225616 155582 225644 159200
rect 225972 156596 226024 156602
rect 225972 156538 226024 156544
rect 225604 155576 225656 155582
rect 225604 155518 225656 155524
rect 225984 151994 226012 156538
rect 226628 155446 226656 159200
rect 226524 155440 226576 155446
rect 226524 155382 226576 155388
rect 226616 155440 226668 155446
rect 226616 155382 226668 155388
rect 226536 151994 226564 155382
rect 227258 155272 227314 155281
rect 227258 155207 227314 155216
rect 227272 151994 227300 155207
rect 227548 154086 227576 159200
rect 228560 156806 228588 159200
rect 228548 156800 228600 156806
rect 228548 156742 228600 156748
rect 228548 156324 228600 156330
rect 228548 156266 228600 156272
rect 227536 154080 227588 154086
rect 227536 154022 227588 154028
rect 227904 153060 227956 153066
rect 227904 153002 227956 153008
rect 227916 151994 227944 153002
rect 228560 151994 228588 156266
rect 229376 155712 229428 155718
rect 229376 155654 229428 155660
rect 229388 155582 229416 155654
rect 229480 155582 229508 159200
rect 229376 155576 229428 155582
rect 229376 155518 229428 155524
rect 229468 155576 229520 155582
rect 229468 155518 229520 155524
rect 229284 155372 229336 155378
rect 229284 155314 229336 155320
rect 229296 151994 229324 155314
rect 230492 155281 230520 159200
rect 230572 156936 230624 156942
rect 230572 156878 230624 156884
rect 230478 155272 230534 155281
rect 230478 155207 230534 155216
rect 229836 154148 229888 154154
rect 229836 154090 229888 154096
rect 229848 151994 229876 154090
rect 230584 151994 230612 156878
rect 231504 154154 231532 159200
rect 231860 157004 231912 157010
rect 231860 156946 231912 156952
rect 231492 154148 231544 154154
rect 231492 154090 231544 154096
rect 231446 152108 231498 152114
rect 231446 152050 231498 152056
rect 212552 151966 212612 151994
rect 213932 151966 213992 151994
rect 214300 151966 214636 151994
rect 214944 151966 215280 151994
rect 215588 151966 215924 151994
rect 216232 151966 216568 151994
rect 216876 151966 217212 151994
rect 217520 151966 217856 151994
rect 218164 151966 218500 151994
rect 218900 151966 219144 151994
rect 219636 151966 219788 151994
rect 220096 151966 220432 151994
rect 220832 151966 221076 151994
rect 221384 151966 221720 151994
rect 222212 151966 222364 151994
rect 222764 151966 223100 151994
rect 223592 151966 223744 151994
rect 224052 151966 224388 151994
rect 224972 151966 225032 151994
rect 225340 151966 225676 151994
rect 225984 151966 226320 151994
rect 226536 151966 226964 151994
rect 227272 151966 227608 151994
rect 227916 151966 228252 151994
rect 228560 151966 228896 151994
rect 229296 151966 229540 151994
rect 229848 151966 230184 151994
rect 230584 151966 230828 151994
rect 231458 151980 231486 152050
rect 231872 151994 231900 156946
rect 232424 152862 232452 159200
rect 233436 156874 233464 159200
rect 233424 156868 233476 156874
rect 233424 156810 233476 156816
rect 233792 156256 233844 156262
rect 233792 156198 233844 156204
rect 232504 154216 232556 154222
rect 232504 154158 232556 154164
rect 232412 152856 232464 152862
rect 232412 152798 232464 152804
rect 232516 151994 232544 154158
rect 233240 153196 233292 153202
rect 233240 153138 233292 153144
rect 233252 151994 233280 153138
rect 233804 151994 233832 156198
rect 234356 155825 234384 159200
rect 234342 155816 234398 155825
rect 234342 155751 234398 155760
rect 235080 155780 235132 155786
rect 235080 155722 235132 155728
rect 234618 155408 234674 155417
rect 234618 155343 234674 155352
rect 234632 151994 234660 155343
rect 235092 151994 235120 155722
rect 235368 154222 235396 159200
rect 236000 157072 236052 157078
rect 236000 157014 236052 157020
rect 235356 154216 235408 154222
rect 235356 154158 235408 154164
rect 236012 151994 236040 157014
rect 236288 156942 236316 159200
rect 236276 156936 236328 156942
rect 236276 156878 236328 156884
rect 237300 155718 237328 159200
rect 237012 155712 237064 155718
rect 237012 155654 237064 155660
rect 237288 155712 237340 155718
rect 237288 155654 237340 155660
rect 236690 152244 236742 152250
rect 236690 152186 236742 152192
rect 231872 151966 232208 151994
rect 232516 151966 232852 151994
rect 233252 151966 233496 151994
rect 233804 151966 234140 151994
rect 234632 151966 234784 151994
rect 235092 151966 235428 151994
rect 236012 151966 236072 151994
rect 236702 151980 236730 152186
rect 237024 151994 237052 155654
rect 237656 154284 237708 154290
rect 237656 154226 237708 154232
rect 237668 151994 237696 154226
rect 238312 152930 238340 159200
rect 238392 157140 238444 157146
rect 238392 157082 238444 157088
rect 238300 152924 238352 152930
rect 238300 152866 238352 152872
rect 238404 151994 238432 157082
rect 239036 156392 239088 156398
rect 239036 156334 239088 156340
rect 239048 151994 239076 156334
rect 239232 154290 239260 159200
rect 240244 157010 240272 159200
rect 240232 157004 240284 157010
rect 240232 156946 240284 156952
rect 240232 155168 240284 155174
rect 240232 155110 240284 155116
rect 239220 154284 239272 154290
rect 239220 154226 239272 154232
rect 239588 152380 239640 152386
rect 239588 152322 239640 152328
rect 239600 151994 239628 152322
rect 240244 151994 240272 155110
rect 241164 154902 241192 159200
rect 241612 156120 241664 156126
rect 241612 156062 241664 156068
rect 241152 154896 241204 154902
rect 241152 154838 241204 154844
rect 240968 152312 241020 152318
rect 240968 152254 241020 152260
rect 240980 151994 241008 152254
rect 241624 151994 241652 156062
rect 242176 155922 242204 159200
rect 242164 155916 242216 155922
rect 242164 155858 242216 155864
rect 242256 155032 242308 155038
rect 242256 154974 242308 154980
rect 242268 151994 242296 154974
rect 243188 154358 243216 159200
rect 244108 157078 244136 159200
rect 244096 157072 244148 157078
rect 244096 157014 244148 157020
rect 243452 155100 243504 155106
rect 243452 155042 243504 155048
rect 244832 155100 244884 155106
rect 244832 155042 244884 155048
rect 243464 155009 243492 155042
rect 243450 155000 243506 155009
rect 243450 154935 243506 154944
rect 242900 154352 242952 154358
rect 242900 154294 242952 154300
rect 243176 154352 243228 154358
rect 243176 154294 243228 154300
rect 242912 151994 242940 154294
rect 243866 152176 243918 152182
rect 243866 152118 243918 152124
rect 237024 151966 237360 151994
rect 237668 151966 238004 151994
rect 238404 151966 238648 151994
rect 239048 151966 239292 151994
rect 239600 151966 239936 151994
rect 240244 151966 240580 151994
rect 240980 151966 241316 151994
rect 241624 151966 241960 151994
rect 242268 151966 242604 151994
rect 242912 151966 243248 151994
rect 243878 151980 243906 152118
rect 244844 151994 244872 155042
rect 245120 154970 245148 159200
rect 246040 155786 246068 159200
rect 246120 157208 246172 157214
rect 246120 157150 246172 157156
rect 246028 155780 246080 155786
rect 246028 155722 246080 155728
rect 245108 154964 245160 154970
rect 245108 154906 245160 154912
rect 245660 154420 245712 154426
rect 245660 154362 245712 154368
rect 245672 151994 245700 154362
rect 246132 151994 246160 157150
rect 247052 155718 247080 159200
rect 248064 157334 248092 159200
rect 248064 157306 248184 157334
rect 247224 156188 247276 156194
rect 247224 156130 247276 156136
rect 246948 155712 247000 155718
rect 246948 155654 247000 155660
rect 247040 155712 247092 155718
rect 247040 155654 247092 155660
rect 246960 155530 246988 155654
rect 246960 155502 247080 155530
rect 247052 154834 247080 155502
rect 246948 154828 247000 154834
rect 246948 154770 247000 154776
rect 247040 154828 247092 154834
rect 247040 154770 247092 154776
rect 246960 153406 246988 154770
rect 246948 153400 247000 153406
rect 246948 153342 247000 153348
rect 244844 151966 245180 151994
rect 245672 151966 245824 151994
rect 246132 151966 246468 151994
rect 244372 151904 244424 151910
rect 247236 151858 247264 156130
rect 247408 154828 247460 154834
rect 247408 154770 247460 154776
rect 247420 151994 247448 154770
rect 248052 154488 248104 154494
rect 248052 154430 248104 154436
rect 248064 151994 248092 154430
rect 248156 152998 248184 157306
rect 248696 157276 248748 157282
rect 248696 157218 248748 157224
rect 248144 152992 248196 152998
rect 248144 152934 248196 152940
rect 248708 151994 248736 157218
rect 248984 154834 249012 159200
rect 249064 155644 249116 155650
rect 249064 155586 249116 155592
rect 248972 154828 249024 154834
rect 248972 154770 249024 154776
rect 249076 154426 249104 155586
rect 249996 155174 250024 159200
rect 250916 155650 250944 159200
rect 251928 157146 251956 159200
rect 251916 157140 251968 157146
rect 251916 157082 251968 157088
rect 252940 155854 252968 159200
rect 252928 155848 252980 155854
rect 252928 155790 252980 155796
rect 250904 155644 250956 155650
rect 250904 155586 250956 155592
rect 253860 155242 253888 159200
rect 253940 157344 253992 157350
rect 253940 157286 253992 157292
rect 252652 155236 252704 155242
rect 252652 155178 252704 155184
rect 253848 155236 253900 155242
rect 253848 155178 253900 155184
rect 249984 155168 250036 155174
rect 249984 155110 250036 155116
rect 249798 155000 249854 155009
rect 249798 154935 249854 154944
rect 249064 154420 249116 154426
rect 249064 154362 249116 154368
rect 249812 153542 249840 154935
rect 252560 154692 252612 154698
rect 252560 154634 252612 154640
rect 252572 154562 252600 154634
rect 252560 154556 252612 154562
rect 252560 154498 252612 154504
rect 249984 154488 250036 154494
rect 249984 154430 250036 154436
rect 249800 153536 249852 153542
rect 249800 153478 249852 153484
rect 249996 151994 250024 154430
rect 250720 153400 250772 153406
rect 250720 153342 250772 153348
rect 250732 151994 250760 153342
rect 251364 152040 251416 152046
rect 247420 151966 247756 151994
rect 248064 151966 248400 151994
rect 248708 151966 249044 151994
rect 249352 151978 249688 151994
rect 249340 151972 249688 151978
rect 249392 151966 249688 151972
rect 249996 151966 250332 151994
rect 250732 151966 251068 151994
rect 252664 151994 252692 155178
rect 253296 154488 253348 154494
rect 253296 154430 253348 154436
rect 253308 151994 253336 154430
rect 253952 151994 253980 157286
rect 254584 156460 254636 156466
rect 254584 156402 254636 156408
rect 254596 151994 254624 156402
rect 254872 154834 254900 159200
rect 255412 155916 255464 155922
rect 255412 155858 255464 155864
rect 255320 154896 255372 154902
rect 255320 154838 255372 154844
rect 254860 154828 254912 154834
rect 254860 154770 254912 154776
rect 255332 154494 255360 154838
rect 255320 154488 255372 154494
rect 255320 154430 255372 154436
rect 255424 151994 255452 155858
rect 255792 153066 255820 159200
rect 256700 156528 256752 156534
rect 256700 156470 256752 156476
rect 255872 153876 255924 153882
rect 255872 153818 255924 153824
rect 255780 153060 255832 153066
rect 255780 153002 255832 153008
rect 255884 151994 255912 153818
rect 256712 151994 256740 156470
rect 256804 154698 256832 159200
rect 257816 155922 257844 159200
rect 258080 156664 258132 156670
rect 258080 156606 258132 156612
rect 257804 155916 257856 155922
rect 257804 155858 257856 155864
rect 256792 154692 256844 154698
rect 256792 154634 256844 154640
rect 257160 153536 257212 153542
rect 257160 153478 257212 153484
rect 257172 151994 257200 153478
rect 258092 151994 258120 156606
rect 258736 155378 258764 159200
rect 258724 155372 258776 155378
rect 258724 155314 258776 155320
rect 259368 155100 259420 155106
rect 259368 155042 259420 155048
rect 259380 153542 259408 155042
rect 259368 153536 259420 153542
rect 259368 153478 259420 153484
rect 259092 152720 259144 152726
rect 259092 152662 259144 152668
rect 258448 152516 258500 152522
rect 258448 152458 258500 152464
rect 258460 151994 258488 152458
rect 259104 151994 259132 152662
rect 259748 152522 259776 159200
rect 259828 156052 259880 156058
rect 259828 155994 259880 156000
rect 259736 152516 259788 152522
rect 259736 152458 259788 152464
rect 259840 151994 259868 155994
rect 260668 155378 260696 159200
rect 260930 155544 260986 155553
rect 260930 155479 260986 155488
rect 260564 155372 260616 155378
rect 260564 155314 260616 155320
rect 260656 155372 260708 155378
rect 260656 155314 260708 155320
rect 260576 153814 260604 155314
rect 260564 153808 260616 153814
rect 260564 153750 260616 153756
rect 260944 153678 260972 155479
rect 261680 155417 261708 159200
rect 261760 156732 261812 156738
rect 261760 156674 261812 156680
rect 261666 155408 261722 155417
rect 261666 155343 261722 155352
rect 261116 154420 261168 154426
rect 261116 154362 261168 154368
rect 260932 153672 260984 153678
rect 260932 153614 260984 153620
rect 260472 153536 260524 153542
rect 260472 153478 260524 153484
rect 260484 151994 260512 153478
rect 261128 151994 261156 154362
rect 261772 151994 261800 156674
rect 262218 155680 262274 155689
rect 262218 155615 262274 155624
rect 262232 153746 262260 155615
rect 262404 154556 262456 154562
rect 262404 154498 262456 154504
rect 262220 153740 262272 153746
rect 262220 153682 262272 153688
rect 262416 151994 262444 154498
rect 262692 154426 262720 159200
rect 263612 156670 263640 159200
rect 263600 156664 263652 156670
rect 263600 156606 263652 156612
rect 262864 154896 262916 154902
rect 262864 154838 262916 154844
rect 262876 154766 262904 154838
rect 264624 154766 264652 159200
rect 265072 155984 265124 155990
rect 265072 155926 265124 155932
rect 264980 155576 265032 155582
rect 264980 155518 265032 155524
rect 262864 154760 262916 154766
rect 262864 154702 262916 154708
rect 264612 154760 264664 154766
rect 264612 154702 264664 154708
rect 263600 154692 263652 154698
rect 263600 154634 263652 154640
rect 262680 154420 262732 154426
rect 262680 154362 262732 154368
rect 263612 153950 263640 154634
rect 264992 154562 265020 155518
rect 264980 154556 265032 154562
rect 264980 154498 265032 154504
rect 263600 153944 263652 153950
rect 263600 153886 263652 153892
rect 263692 153876 263744 153882
rect 263692 153818 263744 153824
rect 263048 153672 263100 153678
rect 263048 153614 263100 153620
rect 263060 151994 263088 153614
rect 263704 151994 263732 153818
rect 264336 152652 264388 152658
rect 264336 152594 264388 152600
rect 264348 151994 264376 152594
rect 265084 151994 265112 155926
rect 265544 155378 265572 159200
rect 266556 155582 266584 159200
rect 266544 155576 266596 155582
rect 266544 155518 266596 155524
rect 265532 155372 265584 155378
rect 265532 155314 265584 155320
rect 266360 154012 266412 154018
rect 266360 153954 266412 153960
rect 265624 153740 265676 153746
rect 265624 153682 265676 153688
rect 265636 151994 265664 153682
rect 266372 151994 266400 153954
rect 267568 152590 267596 159200
rect 268488 154970 268516 159200
rect 269500 155446 269528 159200
rect 269396 155440 269448 155446
rect 269396 155382 269448 155388
rect 269488 155440 269540 155446
rect 269488 155382 269540 155388
rect 269028 155304 269080 155310
rect 269028 155246 269080 155252
rect 268476 154964 268528 154970
rect 268476 154906 268528 154912
rect 267832 154488 267884 154494
rect 267832 154430 267884 154436
rect 266912 152584 266964 152590
rect 266912 152526 266964 152532
rect 267556 152584 267608 152590
rect 267556 152526 267608 152532
rect 266924 151994 266952 152526
rect 267844 151994 267872 154430
rect 268200 153400 268252 153406
rect 268200 153342 268252 153348
rect 268212 151994 268240 153342
rect 269040 153218 269068 155246
rect 269408 153678 269436 155382
rect 270420 155310 270448 159200
rect 270408 155304 270460 155310
rect 270408 155246 270460 155252
rect 270408 154896 270460 154902
rect 270408 154838 270460 154844
rect 270420 153814 270448 154838
rect 270500 153944 270552 153950
rect 270500 153886 270552 153892
rect 270408 153808 270460 153814
rect 270408 153750 270460 153756
rect 269396 153672 269448 153678
rect 269396 153614 269448 153620
rect 269040 153190 269160 153218
rect 269132 151994 269160 153190
rect 269580 152788 269632 152794
rect 269580 152730 269632 152736
rect 269592 151994 269620 152730
rect 270512 151994 270540 153886
rect 270868 153672 270920 153678
rect 270868 153614 270920 153620
rect 270880 151994 270908 153614
rect 271432 152658 271460 159200
rect 272352 159174 272472 159200
rect 272156 156800 272208 156806
rect 272156 156742 272208 156748
rect 271788 154488 271840 154494
rect 271788 154430 271840 154436
rect 271512 154080 271564 154086
rect 271512 154022 271564 154028
rect 271420 152652 271472 152658
rect 271420 152594 271472 152600
rect 271524 151994 271552 154022
rect 271800 153474 271828 154430
rect 271788 153468 271840 153474
rect 271788 153410 271840 153416
rect 272168 151994 272196 156742
rect 272812 155378 272840 159310
rect 273350 159200 273406 160000
rect 274362 159200 274418 160000
rect 275282 159200 275338 160000
rect 276294 159200 276350 160000
rect 277214 159200 277270 160000
rect 278226 159200 278282 160000
rect 279238 159200 279294 160000
rect 280158 159200 280214 160000
rect 281170 159200 281226 160000
rect 282090 159200 282146 160000
rect 283102 159200 283158 160000
rect 284114 159200 284170 160000
rect 285034 159200 285090 160000
rect 286046 159200 286102 160000
rect 286966 159200 287022 160000
rect 287978 159200 288034 160000
rect 288990 159200 289046 160000
rect 289910 159200 289966 160000
rect 290922 159200 290978 160000
rect 291842 159200 291898 160000
rect 292854 159200 292910 160000
rect 293866 159200 293922 160000
rect 294786 159200 294842 160000
rect 295798 159200 295854 160000
rect 296718 159200 296774 160000
rect 297730 159200 297786 160000
rect 298742 159200 298798 160000
rect 299662 159200 299718 160000
rect 300674 159200 300730 160000
rect 301594 159200 301650 160000
rect 302606 159200 302662 160000
rect 303618 159200 303674 160000
rect 304538 159200 304594 160000
rect 305550 159200 305606 160000
rect 306470 159200 306526 160000
rect 307482 159200 307538 160000
rect 308494 159200 308550 160000
rect 309414 159200 309470 160000
rect 310426 159200 310482 160000
rect 311346 159200 311402 160000
rect 312358 159200 312414 160000
rect 313278 159200 313334 160000
rect 314290 159200 314346 160000
rect 315302 159200 315358 160000
rect 316222 159202 316278 160000
rect 316328 159310 316632 159338
rect 316328 159202 316356 159310
rect 316222 159200 316356 159202
rect 272800 155372 272852 155378
rect 272800 155314 272852 155320
rect 273166 155272 273222 155281
rect 273166 155207 273222 155216
rect 272800 154556 272852 154562
rect 272800 154498 272852 154504
rect 272812 151994 272840 154498
rect 273180 153218 273208 155207
rect 273364 154834 273392 159200
rect 274376 155281 274404 159200
rect 275296 155310 275324 159200
rect 275376 156868 275428 156874
rect 275376 156810 275428 156816
rect 275284 155304 275336 155310
rect 274362 155272 274418 155281
rect 275284 155246 275336 155252
rect 274362 155207 274418 155216
rect 273260 154828 273312 154834
rect 273260 154770 273312 154776
rect 273352 154828 273404 154834
rect 273352 154770 273404 154776
rect 273272 154154 273300 154770
rect 273352 154488 273404 154494
rect 273352 154430 273404 154436
rect 273260 154148 273312 154154
rect 273260 154090 273312 154096
rect 273364 153746 273392 154430
rect 274088 154080 274140 154086
rect 274088 154022 274140 154028
rect 273352 153740 273404 153746
rect 273352 153682 273404 153688
rect 273180 153190 273392 153218
rect 273364 151994 273392 153190
rect 274100 151994 274128 154022
rect 274732 152856 274784 152862
rect 274732 152798 274784 152804
rect 274744 151994 274772 152798
rect 275388 151994 275416 156810
rect 275834 155816 275890 155825
rect 275834 155751 275890 155760
rect 275848 153490 275876 155751
rect 276308 154970 276336 159200
rect 277124 155372 277176 155378
rect 277124 155314 277176 155320
rect 276296 154964 276348 154970
rect 276296 154906 276348 154912
rect 277136 154873 277164 155314
rect 277122 154864 277178 154873
rect 277122 154799 277178 154808
rect 277228 154698 277256 159200
rect 277584 156936 277636 156942
rect 277584 156878 277636 156884
rect 277400 155644 277452 155650
rect 277400 155586 277452 155592
rect 277412 155530 277440 155586
rect 277412 155502 277532 155530
rect 277504 155446 277532 155502
rect 277492 155440 277544 155446
rect 277492 155382 277544 155388
rect 277492 155032 277544 155038
rect 277492 154974 277544 154980
rect 277504 154873 277532 154974
rect 277490 154864 277546 154873
rect 277490 154799 277546 154808
rect 277216 154692 277268 154698
rect 277216 154634 277268 154640
rect 275928 154624 275980 154630
rect 275980 154572 276060 154578
rect 275928 154566 276060 154572
rect 275940 154550 276060 154566
rect 276032 154018 276060 154550
rect 276664 154216 276716 154222
rect 276664 154158 276716 154164
rect 276020 154012 276072 154018
rect 276020 153954 276072 153960
rect 275848 153462 276060 153490
rect 276032 151994 276060 153462
rect 276676 151994 276704 154158
rect 277596 151994 277624 156878
rect 278240 153950 278268 159200
rect 279252 155446 279280 159200
rect 280172 155650 280200 159200
rect 280252 157004 280304 157010
rect 280252 156946 280304 156952
rect 280160 155644 280212 155650
rect 280160 155586 280212 155592
rect 279148 155440 279200 155446
rect 279148 155382 279200 155388
rect 279240 155440 279292 155446
rect 279240 155382 279292 155388
rect 279160 154873 279188 155382
rect 279146 154864 279202 154873
rect 279146 154799 279202 154808
rect 279332 154760 279384 154766
rect 279332 154702 279384 154708
rect 279344 154494 279372 154702
rect 279332 154488 279384 154494
rect 279332 154430 279384 154436
rect 279332 154284 279384 154290
rect 279332 154226 279384 154232
rect 278228 153944 278280 153950
rect 278228 153886 278280 153892
rect 277952 153468 278004 153474
rect 277952 153410 278004 153416
rect 277964 151994 277992 153410
rect 278780 152924 278832 152930
rect 278780 152866 278832 152872
rect 278792 151994 278820 152866
rect 279344 151994 279372 154226
rect 280264 151994 280292 156946
rect 281184 155786 281212 159200
rect 280712 155780 280764 155786
rect 280712 155722 280764 155728
rect 281172 155780 281224 155786
rect 281172 155722 281224 155728
rect 280620 153808 280672 153814
rect 280620 153750 280672 153756
rect 280632 151994 280660 153750
rect 280724 153406 280752 155722
rect 282104 155718 282132 159200
rect 282552 157072 282604 157078
rect 282552 157014 282604 157020
rect 282092 155712 282144 155718
rect 282092 155654 282144 155660
rect 281540 155508 281592 155514
rect 281540 155450 281592 155456
rect 281448 155168 281500 155174
rect 281448 155110 281500 155116
rect 281460 154086 281488 155110
rect 281448 154080 281500 154086
rect 281448 154022 281500 154028
rect 280712 153400 280764 153406
rect 280712 153342 280764 153348
rect 281552 151994 281580 155450
rect 282366 154864 282422 154873
rect 282366 154799 282422 154808
rect 282380 154630 282408 154799
rect 282368 154624 282420 154630
rect 282368 154566 282420 154572
rect 281908 154352 281960 154358
rect 281908 154294 281960 154300
rect 281920 151994 281948 154294
rect 282564 151994 282592 157014
rect 283116 154834 283144 159200
rect 284128 155514 284156 159200
rect 284024 155508 284076 155514
rect 284024 155450 284076 155456
rect 284116 155508 284168 155514
rect 284116 155450 284168 155456
rect 284036 155394 284064 155450
rect 284036 155366 284340 155394
rect 283104 154828 283156 154834
rect 283104 154770 283156 154776
rect 283196 153740 283248 153746
rect 283196 153682 283248 153688
rect 283208 151994 283236 153682
rect 284312 153542 284340 155366
rect 285048 155106 285076 159200
rect 285036 155100 285088 155106
rect 285036 155042 285088 155048
rect 285680 155032 285732 155038
rect 285680 154974 285732 154980
rect 285692 154290 285720 154974
rect 286060 154834 286088 159200
rect 286980 156058 287008 159200
rect 287796 157140 287848 157146
rect 287796 157082 287848 157088
rect 286968 156052 287020 156058
rect 286968 155994 287020 156000
rect 287060 155984 287112 155990
rect 287060 155926 287112 155932
rect 286968 155916 287020 155922
rect 286968 155858 287020 155864
rect 286980 155802 287008 155858
rect 286704 155786 287008 155802
rect 286692 155780 287008 155786
rect 286744 155774 287008 155780
rect 286692 155722 286744 155728
rect 286048 154828 286100 154834
rect 286048 154770 286100 154776
rect 285864 154624 285916 154630
rect 285864 154566 285916 154572
rect 284484 154284 284536 154290
rect 284484 154226 284536 154232
rect 285680 154284 285732 154290
rect 285680 154226 285732 154232
rect 284300 153536 284352 153542
rect 284300 153478 284352 153484
rect 283840 153400 283892 153406
rect 283840 153342 283892 153348
rect 283852 151994 283880 153342
rect 284496 151994 284524 154226
rect 285772 154148 285824 154154
rect 285772 154090 285824 154096
rect 285128 152992 285180 152998
rect 285128 152934 285180 152940
rect 285140 151994 285168 152934
rect 285784 151994 285812 154090
rect 285876 153406 285904 154566
rect 287072 153814 287100 155926
rect 287060 153808 287112 153814
rect 287060 153750 287112 153756
rect 286416 153536 286468 153542
rect 286416 153478 286468 153484
rect 285864 153400 285916 153406
rect 285864 153342 285916 153348
rect 286428 151994 286456 153478
rect 287244 153400 287296 153406
rect 287244 153342 287296 153348
rect 287256 151994 287284 153342
rect 287808 151994 287836 157082
rect 287992 155854 288020 159200
rect 287980 155848 288032 155854
rect 287980 155790 288032 155796
rect 289004 155582 289032 159200
rect 289924 155922 289952 159200
rect 289912 155916 289964 155922
rect 289912 155858 289964 155864
rect 288992 155576 289044 155582
rect 288992 155518 289044 155524
rect 290936 155378 290964 159200
rect 291856 155650 291884 159200
rect 291752 155644 291804 155650
rect 291752 155586 291804 155592
rect 291844 155644 291896 155650
rect 291844 155586 291896 155592
rect 290004 155372 290056 155378
rect 290004 155314 290056 155320
rect 290924 155372 290976 155378
rect 290924 155314 290976 155320
rect 289728 154692 289780 154698
rect 289728 154634 289780 154640
rect 288440 154556 288492 154562
rect 288440 154498 288492 154504
rect 288452 151994 288480 154498
rect 289084 153808 289136 153814
rect 289084 153750 289136 153756
rect 289096 151994 289124 153750
rect 289740 153218 289768 154634
rect 290016 153814 290044 155314
rect 291108 154896 291160 154902
rect 291108 154838 291160 154844
rect 291120 154358 291148 154838
rect 291568 154556 291620 154562
rect 291568 154498 291620 154504
rect 291108 154352 291160 154358
rect 291108 154294 291160 154300
rect 291200 154012 291252 154018
rect 291200 153954 291252 153960
rect 290004 153808 290056 153814
rect 290004 153750 290056 153756
rect 289740 153190 289860 153218
rect 289832 151994 289860 153190
rect 290372 153060 290424 153066
rect 290372 153002 290424 153008
rect 290384 151994 290412 153002
rect 291212 151994 291240 153954
rect 291580 153542 291608 154498
rect 291764 154154 291792 155586
rect 292868 154902 292896 159200
rect 293040 155848 293092 155854
rect 293040 155790 293092 155796
rect 292856 154896 292908 154902
rect 292856 154838 292908 154844
rect 291752 154148 291804 154154
rect 291752 154090 291804 154096
rect 293052 154018 293080 155790
rect 293880 155582 293908 159200
rect 294800 155854 294828 159200
rect 295524 156664 295576 156670
rect 295524 156606 295576 156612
rect 294788 155848 294840 155854
rect 294788 155790 294840 155796
rect 293868 155576 293920 155582
rect 293868 155518 293920 155524
rect 293866 155408 293922 155417
rect 293866 155343 293922 155352
rect 293592 154488 293644 154494
rect 293592 154430 293644 154436
rect 293040 154012 293092 154018
rect 293040 153954 293092 153960
rect 292580 153876 292632 153882
rect 292580 153818 292632 153824
rect 291660 153808 291712 153814
rect 291660 153750 291712 153756
rect 291568 153536 291620 153542
rect 291568 153478 291620 153484
rect 291672 151994 291700 153750
rect 292592 151994 292620 153818
rect 292948 152516 293000 152522
rect 292948 152458 293000 152464
rect 292960 151994 292988 152458
rect 293604 151994 293632 154430
rect 293880 153218 293908 155343
rect 293960 154556 294012 154562
rect 293960 154498 294012 154504
rect 293972 153406 294000 154498
rect 294880 154420 294932 154426
rect 294880 154362 294932 154368
rect 293960 153400 294012 153406
rect 293960 153342 294012 153348
rect 293880 153190 294184 153218
rect 294156 151994 294184 153190
rect 294892 151994 294920 154362
rect 295536 151994 295564 156606
rect 295812 153882 295840 159200
rect 296732 155258 296760 159200
rect 296732 155242 296944 155258
rect 296732 155236 296956 155242
rect 296732 155230 296904 155236
rect 296904 155178 296956 155184
rect 297744 155038 297772 159200
rect 298756 155446 298784 159200
rect 298744 155440 298796 155446
rect 298744 155382 298796 155388
rect 297916 155168 297968 155174
rect 297916 155110 297968 155116
rect 297732 155032 297784 155038
rect 297732 154974 297784 154980
rect 296168 154080 296220 154086
rect 296168 154022 296220 154028
rect 295800 153876 295852 153882
rect 295800 153818 295852 153824
rect 296180 151994 296208 154022
rect 297928 153542 297956 155110
rect 298008 154760 298060 154766
rect 298008 154702 298060 154708
rect 297548 153536 297600 153542
rect 297548 153478 297600 153484
rect 297916 153536 297968 153542
rect 297916 153478 297968 153484
rect 296996 153400 297048 153406
rect 296996 153342 297048 153348
rect 297008 151994 297036 153342
rect 297560 151994 297588 153478
rect 298020 153406 298048 154702
rect 299676 154698 299704 159200
rect 300688 155786 300716 159200
rect 300676 155780 300728 155786
rect 300676 155722 300728 155728
rect 301608 155310 301636 159200
rect 300124 155304 300176 155310
rect 300124 155246 300176 155252
rect 301596 155304 301648 155310
rect 301596 155246 301648 155252
rect 299572 154692 299624 154698
rect 299572 154634 299624 154640
rect 299664 154692 299716 154698
rect 299664 154634 299716 154640
rect 298836 154216 298888 154222
rect 298836 154158 298888 154164
rect 298008 153400 298060 153406
rect 298008 153342 298060 153348
rect 298192 152584 298244 152590
rect 298192 152526 298244 152532
rect 298204 151994 298232 152526
rect 298848 151994 298876 154158
rect 299480 153536 299532 153542
rect 299480 153478 299532 153484
rect 299492 151994 299520 153478
rect 299584 153474 299612 154634
rect 299572 153468 299624 153474
rect 299572 153410 299624 153416
rect 300136 151994 300164 155246
rect 302240 155100 302292 155106
rect 302240 155042 302292 155048
rect 301412 154284 301464 154290
rect 301412 154226 301464 154232
rect 300860 152652 300912 152658
rect 300860 152594 300912 152600
rect 300872 151994 300900 152594
rect 301424 151994 301452 154226
rect 302252 154222 302280 155042
rect 302620 154970 302648 159200
rect 302698 155272 302754 155281
rect 302698 155207 302754 155216
rect 302608 154964 302660 154970
rect 302608 154906 302660 154912
rect 302240 154216 302292 154222
rect 302240 154158 302292 154164
rect 302332 153400 302384 153406
rect 302332 153342 302384 153348
rect 302344 151994 302372 153342
rect 302712 151994 302740 155207
rect 303632 154766 303660 159200
rect 304552 155650 304580 159200
rect 304540 155644 304592 155650
rect 304540 155586 304592 155592
rect 305564 155242 305592 159200
rect 304908 155236 304960 155242
rect 304908 155178 304960 155184
rect 305552 155236 305604 155242
rect 305552 155178 305604 155184
rect 303620 154760 303672 154766
rect 303620 154702 303672 154708
rect 304632 154488 304684 154494
rect 304632 154430 304684 154436
rect 303620 154420 303672 154426
rect 303620 154362 303672 154368
rect 303632 151994 303660 154362
rect 303988 154352 304040 154358
rect 303988 154294 304040 154300
rect 304000 151994 304028 154294
rect 304644 151994 304672 154430
rect 304920 154086 304948 155178
rect 306288 154896 306340 154902
rect 306288 154838 306340 154844
rect 305920 154624 305972 154630
rect 305920 154566 305972 154572
rect 304908 154080 304960 154086
rect 304908 154022 304960 154028
rect 305276 153944 305328 153950
rect 305276 153886 305328 153892
rect 305288 151994 305316 153886
rect 305932 151994 305960 154566
rect 306300 154290 306328 154838
rect 306484 154630 306512 159200
rect 307300 155780 307352 155786
rect 307300 155722 307352 155728
rect 307312 155666 307340 155722
rect 306944 155638 307340 155666
rect 306944 155582 306972 155638
rect 306932 155576 306984 155582
rect 306932 155518 306984 155524
rect 307496 155038 307524 159200
rect 308036 155508 308088 155514
rect 308036 155450 308088 155456
rect 307484 155032 307536 155038
rect 307484 154974 307536 154980
rect 306564 154828 306616 154834
rect 306564 154770 306616 154776
rect 306472 154624 306524 154630
rect 306472 154566 306524 154572
rect 306288 154284 306340 154290
rect 306288 154226 306340 154232
rect 306576 153406 306604 154770
rect 306656 154148 306708 154154
rect 306656 154090 306708 154096
rect 306564 153400 306616 153406
rect 306564 153342 306616 153348
rect 306668 151994 306696 154090
rect 307300 153468 307352 153474
rect 307300 153410 307352 153416
rect 307312 151994 307340 153410
rect 308048 153406 308076 155450
rect 308508 155310 308536 159200
rect 309428 155922 309456 159200
rect 309140 155916 309192 155922
rect 309140 155858 309192 155864
rect 309416 155916 309468 155922
rect 309416 155858 309468 155864
rect 308588 155440 308640 155446
rect 308588 155382 308640 155388
rect 308496 155304 308548 155310
rect 308496 155246 308548 155252
rect 307944 153400 307996 153406
rect 307944 153342 307996 153348
rect 308036 153400 308088 153406
rect 308036 153342 308088 153348
rect 307956 151994 307984 153342
rect 308600 151994 308628 155382
rect 309152 153950 309180 155858
rect 309232 155780 309284 155786
rect 309232 155722 309284 155728
rect 309140 153944 309192 153950
rect 309140 153886 309192 153892
rect 309244 151994 309272 155722
rect 310440 155514 310468 159200
rect 310428 155508 310480 155514
rect 310428 155450 310480 155456
rect 311360 155446 311388 159200
rect 312372 155786 312400 159200
rect 312360 155780 312412 155786
rect 312360 155722 312412 155728
rect 311992 155644 312044 155650
rect 311992 155586 312044 155592
rect 311164 155440 311216 155446
rect 311164 155382 311216 155388
rect 311348 155440 311400 155446
rect 311348 155382 311400 155388
rect 309876 154556 309928 154562
rect 309876 154498 309928 154504
rect 309888 151994 309916 154498
rect 310520 153400 310572 153406
rect 310520 153342 310572 153348
rect 310532 151994 310560 153342
rect 311176 151994 311204 155382
rect 312004 154018 312032 155586
rect 313096 155576 313148 155582
rect 313148 155524 313228 155530
rect 313096 155518 313228 155524
rect 313108 155502 313228 155518
rect 313292 155514 313320 159200
rect 314304 155718 314332 159200
rect 315316 155922 315344 159200
rect 316236 159174 316356 159200
rect 315304 155916 315356 155922
rect 315304 155858 315356 155864
rect 316040 155848 316092 155854
rect 316040 155790 316092 155796
rect 313740 155712 313792 155718
rect 313740 155654 313792 155660
rect 314292 155712 314344 155718
rect 314292 155654 314344 155660
rect 313200 155394 313228 155502
rect 313280 155508 313332 155514
rect 313280 155450 313332 155456
rect 313200 155366 313320 155394
rect 312452 154216 312504 154222
rect 312452 154158 312504 154164
rect 311900 154012 311952 154018
rect 311900 153954 311952 153960
rect 311992 154012 312044 154018
rect 311992 153954 312044 153960
rect 311912 151994 311940 153954
rect 312464 151994 312492 154158
rect 313292 151994 313320 155366
rect 313752 151994 313780 155654
rect 314660 155100 314712 155106
rect 314660 155042 314712 155048
rect 314672 151994 314700 155042
rect 315028 154284 315080 154290
rect 315028 154226 315080 154232
rect 315040 151994 315068 154226
rect 316052 151994 316080 155790
rect 316408 155168 316460 155174
rect 316408 155110 316460 155116
rect 316420 151994 316448 155110
rect 316604 154902 316632 159310
rect 317234 159200 317290 160000
rect 318154 159200 318210 160000
rect 319166 159200 319222 160000
rect 320178 159200 320234 160000
rect 321098 159200 321154 160000
rect 322110 159200 322166 160000
rect 323030 159200 323086 160000
rect 324042 159200 324098 160000
rect 325054 159200 325110 160000
rect 325974 159200 326030 160000
rect 326986 159200 327042 160000
rect 327906 159200 327962 160000
rect 328918 159200 328974 160000
rect 329930 159200 329986 160000
rect 330850 159200 330906 160000
rect 331862 159200 331918 160000
rect 332782 159200 332838 160000
rect 333794 159200 333850 160000
rect 334806 159200 334862 160000
rect 335726 159200 335782 160000
rect 336738 159200 336794 160000
rect 337658 159200 337714 160000
rect 338670 159200 338726 160000
rect 339682 159200 339738 160000
rect 340602 159200 340658 160000
rect 341614 159200 341670 160000
rect 342534 159200 342590 160000
rect 343546 159200 343602 160000
rect 344558 159200 344614 160000
rect 345478 159200 345534 160000
rect 346490 159200 346546 160000
rect 347410 159202 347466 160000
rect 347516 159310 347728 159338
rect 347516 159202 347544 159310
rect 347410 159200 347544 159202
rect 317248 155106 317276 159200
rect 317236 155100 317288 155106
rect 317236 155042 317288 155048
rect 316592 154896 316644 154902
rect 316592 154838 316644 154844
rect 317328 154828 317380 154834
rect 317328 154770 317380 154776
rect 317052 153876 317104 153882
rect 317052 153818 317104 153824
rect 317064 151994 317092 153818
rect 317340 153406 317368 154770
rect 318168 154698 318196 159200
rect 319180 155582 319208 159200
rect 320192 155854 320220 159200
rect 320180 155848 320232 155854
rect 320180 155790 320232 155796
rect 319168 155576 319220 155582
rect 319168 155518 319220 155524
rect 321112 155378 321140 159200
rect 322124 155650 322152 159200
rect 321652 155644 321704 155650
rect 321652 155586 321704 155592
rect 322112 155644 322164 155650
rect 322112 155586 322164 155592
rect 318984 155372 319036 155378
rect 318984 155314 319036 155320
rect 321100 155372 321152 155378
rect 321100 155314 321152 155320
rect 318156 154692 318208 154698
rect 318156 154634 318208 154640
rect 317696 154080 317748 154086
rect 317696 154022 317748 154028
rect 317328 153400 317380 153406
rect 317328 153342 317380 153348
rect 317708 151994 317736 154022
rect 318340 153400 318392 153406
rect 318340 153342 318392 153348
rect 318352 151994 318380 153342
rect 318996 151994 319024 155314
rect 320088 155168 320140 155174
rect 320088 155110 320140 155116
rect 319628 154964 319680 154970
rect 319628 154906 319680 154912
rect 319640 151994 319668 154906
rect 320100 153474 320128 155110
rect 321560 155032 321612 155038
rect 321560 154974 321612 154980
rect 320916 154488 320968 154494
rect 320916 154430 320968 154436
rect 320272 153944 320324 153950
rect 320272 153886 320324 153892
rect 320088 153468 320140 153474
rect 320088 153410 320140 153416
rect 320284 151994 320312 153886
rect 320928 151994 320956 154430
rect 321572 151994 321600 154974
rect 321664 153610 321692 155586
rect 323044 155242 323072 159200
rect 322848 155236 322900 155242
rect 322848 155178 322900 155184
rect 323032 155236 323084 155242
rect 323032 155178 323084 155184
rect 321744 154828 321796 154834
rect 321744 154770 321796 154776
rect 321756 153678 321784 154770
rect 322204 154760 322256 154766
rect 322204 154702 322256 154708
rect 321744 153672 321796 153678
rect 321744 153614 321796 153620
rect 321652 153604 321704 153610
rect 321652 153546 321704 153552
rect 322216 151994 322244 154702
rect 322860 153542 322888 155178
rect 324056 155174 324084 159200
rect 324412 155304 324464 155310
rect 324412 155246 324464 155252
rect 324044 155168 324096 155174
rect 324044 155110 324096 155116
rect 324320 154556 324372 154562
rect 324320 154498 324372 154504
rect 322940 154012 322992 154018
rect 322940 153954 322992 153960
rect 322848 153536 322900 153542
rect 322848 153478 322900 153484
rect 322952 151994 322980 153954
rect 323492 153536 323544 153542
rect 323492 153478 323544 153484
rect 323504 151994 323532 153478
rect 324332 151994 324360 154498
rect 324424 153406 324452 155246
rect 325068 155038 325096 159200
rect 325056 155032 325108 155038
rect 325056 154974 325108 154980
rect 325988 154970 326016 159200
rect 326804 155780 326856 155786
rect 326804 155722 326856 155728
rect 326712 155440 326764 155446
rect 326712 155382 326764 155388
rect 325976 154964 326028 154970
rect 325976 154906 326028 154912
rect 326724 153678 326752 155382
rect 326816 153814 326844 155722
rect 327000 155106 327028 159200
rect 327920 155446 327948 159200
rect 328932 155854 328960 159200
rect 329944 155922 329972 159200
rect 329748 155916 329800 155922
rect 329748 155858 329800 155864
rect 329932 155916 329984 155922
rect 329932 155858 329984 155864
rect 328920 155848 328972 155854
rect 328920 155790 328972 155796
rect 328184 155712 328236 155718
rect 328184 155654 328236 155660
rect 327908 155440 327960 155446
rect 327908 155382 327960 155388
rect 326896 155100 326948 155106
rect 326896 155042 326948 155048
rect 326988 155100 327040 155106
rect 326988 155042 327040 155048
rect 326908 154986 326936 155042
rect 326908 154958 327120 154986
rect 326804 153808 326856 153814
rect 326804 153750 326856 153756
rect 327092 153746 327120 154958
rect 328196 153814 328224 155654
rect 328368 155508 328420 155514
rect 328368 155450 328420 155456
rect 328092 153808 328144 153814
rect 328092 153750 328144 153756
rect 328184 153808 328236 153814
rect 328184 153750 328236 153756
rect 327080 153740 327132 153746
rect 327080 153682 327132 153688
rect 326712 153672 326764 153678
rect 326712 153614 326764 153620
rect 327448 153672 327500 153678
rect 327448 153614 327500 153620
rect 327080 153604 327132 153610
rect 327080 153546 327132 153552
rect 324872 153468 324924 153474
rect 324872 153410 324924 153416
rect 326160 153468 326212 153474
rect 326160 153410 326212 153416
rect 324412 153400 324464 153406
rect 324412 153342 324464 153348
rect 324884 151994 324912 153410
rect 325792 153400 325844 153406
rect 325792 153342 325844 153348
rect 325804 151994 325832 153342
rect 326172 151994 326200 153410
rect 327092 151994 327120 153546
rect 327460 151994 327488 153614
rect 328104 151994 328132 153750
rect 328380 153218 328408 155450
rect 329380 153808 329432 153814
rect 329380 153750 329432 153756
rect 328380 153190 328684 153218
rect 328656 151994 328684 153190
rect 329392 151994 329420 153750
rect 329760 153218 329788 155858
rect 330864 155514 330892 159200
rect 330852 155508 330904 155514
rect 330852 155450 330904 155456
rect 331876 155310 331904 159200
rect 332600 155576 332652 155582
rect 332600 155518 332652 155524
rect 331864 155304 331916 155310
rect 331864 155246 331916 155252
rect 330668 154556 330720 154562
rect 330668 154498 330720 154504
rect 329760 153190 329972 153218
rect 329944 151994 329972 153190
rect 330680 151994 330708 154498
rect 331956 154488 332008 154494
rect 331956 154430 332008 154436
rect 331312 153740 331364 153746
rect 331312 153682 331364 153688
rect 331324 151994 331352 153682
rect 331968 151994 331996 154430
rect 332612 151994 332640 155518
rect 332796 154902 332824 159200
rect 333244 155780 333296 155786
rect 333244 155722 333296 155728
rect 332784 154896 332836 154902
rect 332784 154838 332836 154844
rect 333256 151994 333284 155722
rect 333808 155718 333836 159200
rect 334820 155854 334848 159200
rect 334440 155848 334492 155854
rect 334440 155790 334492 155796
rect 334808 155848 334860 155854
rect 334808 155790 334860 155796
rect 333796 155712 333848 155718
rect 333796 155654 333848 155660
rect 334164 155372 334216 155378
rect 334164 155314 334216 155320
rect 334072 155236 334124 155242
rect 334072 155178 334124 155184
rect 333980 155168 334032 155174
rect 333980 155110 334032 155116
rect 333992 153474 334020 155110
rect 333980 153468 334032 153474
rect 333980 153410 334032 153416
rect 334084 153406 334112 155178
rect 334072 153400 334124 153406
rect 334072 153342 334124 153348
rect 334176 151994 334204 155314
rect 334452 153950 334480 155790
rect 334624 155644 334676 155650
rect 334624 155586 334676 155592
rect 334440 153944 334492 153950
rect 334440 153886 334492 153892
rect 334636 151994 334664 155586
rect 335740 155582 335768 159200
rect 336464 155916 336516 155922
rect 336464 155858 336516 155864
rect 335728 155576 335780 155582
rect 335728 155518 335780 155524
rect 336476 153882 336504 155858
rect 336556 155508 336608 155514
rect 336556 155450 336608 155456
rect 336464 153876 336516 153882
rect 336464 153818 336516 153824
rect 336568 153678 336596 155450
rect 336648 155032 336700 155038
rect 336648 154974 336700 154980
rect 336556 153672 336608 153678
rect 336556 153614 336608 153620
rect 335912 153468 335964 153474
rect 335912 153410 335964 153416
rect 335452 153400 335504 153406
rect 335452 153342 335504 153348
rect 335464 151994 335492 153342
rect 335924 151994 335952 153410
rect 336660 153218 336688 154974
rect 336752 154630 336780 159200
rect 337672 155650 337700 159200
rect 338684 155922 338712 159200
rect 338672 155916 338724 155922
rect 338672 155858 338724 155864
rect 339408 155712 339460 155718
rect 339408 155654 339460 155660
rect 337660 155644 337712 155650
rect 337660 155586 337712 155592
rect 338488 155440 338540 155446
rect 338488 155382 338540 155388
rect 337936 155304 337988 155310
rect 337936 155246 337988 155252
rect 337200 154964 337252 154970
rect 337200 154906 337252 154912
rect 336740 154624 336792 154630
rect 336740 154566 336792 154572
rect 336660 153190 336780 153218
rect 336752 151994 336780 153190
rect 337212 151994 337240 154906
rect 337948 153610 337976 155246
rect 338028 155100 338080 155106
rect 338028 155042 338080 155048
rect 337936 153604 337988 153610
rect 337936 153546 337988 153552
rect 338040 153218 338068 155042
rect 338040 153190 338160 153218
rect 338132 151994 338160 153190
rect 338500 151994 338528 155382
rect 338672 154896 338724 154902
rect 338672 154838 338724 154844
rect 338684 153406 338712 154838
rect 339132 153944 339184 153950
rect 339132 153886 339184 153892
rect 338672 153400 338724 153406
rect 338672 153342 338724 153348
rect 339144 151994 339172 153886
rect 339420 153814 339448 155654
rect 339696 154698 339724 159200
rect 340616 154766 340644 159200
rect 340788 155848 340840 155854
rect 340788 155790 340840 155796
rect 340604 154760 340656 154766
rect 340604 154702 340656 154708
rect 339684 154692 339736 154698
rect 339684 154634 339736 154640
rect 340800 153882 340828 155790
rect 340972 155576 341024 155582
rect 340972 155518 341024 155524
rect 340984 154494 341012 155518
rect 341628 154834 341656 159200
rect 342548 155718 342576 159200
rect 342536 155712 342588 155718
rect 342536 155654 342588 155660
rect 342720 155644 342772 155650
rect 342720 155586 342772 155592
rect 341616 154828 341668 154834
rect 341616 154770 341668 154776
rect 340972 154488 341024 154494
rect 340972 154430 341024 154436
rect 339776 153876 339828 153882
rect 339776 153818 339828 153824
rect 340788 153876 340840 153882
rect 340788 153818 340840 153824
rect 339408 153808 339460 153814
rect 339408 153750 339460 153756
rect 339788 151994 339816 153818
rect 342352 153808 342404 153814
rect 342352 153750 342404 153756
rect 340420 153672 340472 153678
rect 340420 153614 340472 153620
rect 340432 151994 340460 153614
rect 341064 153604 341116 153610
rect 341064 153546 341116 153552
rect 341076 151994 341104 153546
rect 341708 153400 341760 153406
rect 341708 153342 341760 153348
rect 341720 151994 341748 153342
rect 342364 151994 342392 153750
rect 342732 153474 342760 155586
rect 343560 155242 343588 159200
rect 344192 155916 344244 155922
rect 344192 155858 344244 155864
rect 343548 155236 343600 155242
rect 343548 155178 343600 155184
rect 343732 154488 343784 154494
rect 343732 154430 343784 154436
rect 342996 153876 343048 153882
rect 342996 153818 343048 153824
rect 342720 153468 342772 153474
rect 342720 153410 342772 153416
rect 343008 151994 343036 153818
rect 343744 151994 343772 154430
rect 344204 153542 344232 155858
rect 344572 155650 344600 159200
rect 344560 155644 344612 155650
rect 344560 155586 344612 155592
rect 345492 154970 345520 159200
rect 345480 154964 345532 154970
rect 345480 154906 345532 154912
rect 346308 154692 346360 154698
rect 346308 154634 346360 154640
rect 344376 154556 344428 154562
rect 344376 154498 344428 154504
rect 344192 153536 344244 153542
rect 344192 153478 344244 153484
rect 344388 151994 344416 154498
rect 345664 153536 345716 153542
rect 345664 153478 345716 153484
rect 345204 153468 345256 153474
rect 345204 153410 345256 153416
rect 345216 151994 345244 153410
rect 345676 151994 345704 153478
rect 346320 153218 346348 154634
rect 346504 154630 346532 159200
rect 347424 159174 347544 159200
rect 347596 154964 347648 154970
rect 347596 154906 347648 154912
rect 347504 154828 347556 154834
rect 347504 154770 347556 154776
rect 346492 154624 346544 154630
rect 346492 154566 346544 154572
rect 347044 154556 347096 154562
rect 347044 154498 347096 154504
rect 346320 153190 346440 153218
rect 346412 151994 346440 153190
rect 347056 151994 347084 154498
rect 347516 153354 347544 154770
rect 347608 154222 347636 154906
rect 347700 154574 347728 159310
rect 348422 159200 348478 160000
rect 349342 159200 349398 160000
rect 350354 159200 350410 160000
rect 351366 159200 351422 160000
rect 352286 159200 352342 160000
rect 353298 159200 353354 160000
rect 354218 159200 354274 160000
rect 355230 159200 355286 160000
rect 356242 159200 356298 160000
rect 357162 159200 357218 160000
rect 358174 159200 358230 160000
rect 359094 159200 359150 160000
rect 360106 159200 360162 160000
rect 361118 159200 361174 160000
rect 362038 159200 362094 160000
rect 363050 159200 363106 160000
rect 363970 159200 364026 160000
rect 364982 159200 365038 160000
rect 365994 159200 366050 160000
rect 366914 159200 366970 160000
rect 367926 159200 367982 160000
rect 368846 159200 368902 160000
rect 369858 159200 369914 160000
rect 370870 159200 370926 160000
rect 371790 159200 371846 160000
rect 372802 159200 372858 160000
rect 373722 159200 373778 160000
rect 374734 159200 374790 160000
rect 375746 159200 375802 160000
rect 376666 159200 376722 160000
rect 377678 159200 377734 160000
rect 378598 159200 378654 160000
rect 379610 159200 379666 160000
rect 380622 159200 380678 160000
rect 381542 159200 381598 160000
rect 382554 159200 382610 160000
rect 383474 159200 383530 160000
rect 384486 159200 384542 160000
rect 385498 159200 385554 160000
rect 386418 159200 386474 160000
rect 387430 159200 387486 160000
rect 388350 159200 388406 160000
rect 389362 159200 389418 160000
rect 390282 159200 390338 160000
rect 391294 159200 391350 160000
rect 392306 159200 392362 160000
rect 393226 159200 393282 160000
rect 394238 159200 394294 160000
rect 395158 159200 395214 160000
rect 396170 159200 396226 160000
rect 397182 159200 397238 160000
rect 398102 159200 398158 160000
rect 398852 159310 399064 159338
rect 348240 155712 348292 155718
rect 348240 155654 348292 155660
rect 347700 154546 347820 154574
rect 347596 154216 347648 154222
rect 347596 154158 347648 154164
rect 347792 154018 347820 154546
rect 347780 154012 347832 154018
rect 347780 153954 347832 153960
rect 347516 153326 347820 153354
rect 347792 151994 347820 153326
rect 348252 151994 348280 155654
rect 348436 154630 348464 159200
rect 349068 155236 349120 155242
rect 349068 155178 349120 155184
rect 348424 154624 348476 154630
rect 348424 154566 348476 154572
rect 349080 153218 349108 155178
rect 349356 154630 349384 159200
rect 349528 155644 349580 155650
rect 349528 155586 349580 155592
rect 349344 154624 349396 154630
rect 349344 154566 349396 154572
rect 349080 153190 349200 153218
rect 349172 151994 349200 153190
rect 349540 151994 349568 155586
rect 350368 154630 350396 159200
rect 351380 154630 351408 159200
rect 352300 154698 352328 159200
rect 353312 155854 353340 159200
rect 354232 155922 354260 159200
rect 354220 155916 354272 155922
rect 354220 155858 354272 155864
rect 353300 155848 353352 155854
rect 353300 155790 353352 155796
rect 355244 155174 355272 159200
rect 355968 155916 356020 155922
rect 355968 155858 356020 155864
rect 355416 155848 355468 155854
rect 355416 155790 355468 155796
rect 355232 155168 355284 155174
rect 355232 155110 355284 155116
rect 352288 154692 352340 154698
rect 352288 154634 352340 154640
rect 353392 154692 353444 154698
rect 353392 154634 353444 154640
rect 350356 154624 350408 154630
rect 350356 154566 350408 154572
rect 351368 154624 351420 154630
rect 351368 154566 351420 154572
rect 352840 154420 352892 154426
rect 352840 154362 352892 154368
rect 352104 154352 352156 154358
rect 352104 154294 352156 154300
rect 350816 154284 350868 154290
rect 350816 154226 350868 154232
rect 350172 154216 350224 154222
rect 350172 154158 350224 154164
rect 350184 151994 350212 154158
rect 350828 151994 350856 154226
rect 351460 154012 351512 154018
rect 351460 153954 351512 153960
rect 351472 151994 351500 153954
rect 352116 151994 352144 154294
rect 352852 151994 352880 154362
rect 353404 153406 353432 154634
rect 354128 154556 354180 154562
rect 354128 154498 354180 154504
rect 353484 154488 353536 154494
rect 353484 154430 353536 154436
rect 353392 153400 353444 153406
rect 353392 153342 353444 153348
rect 353496 151994 353524 154430
rect 354140 151994 354168 154498
rect 354864 153400 354916 153406
rect 354864 153342 354916 153348
rect 354876 151994 354904 153342
rect 355428 151994 355456 155790
rect 355980 153218 356008 155858
rect 356256 155106 356284 159200
rect 356704 155168 356756 155174
rect 356704 155110 356756 155116
rect 356244 155100 356296 155106
rect 356244 155042 356296 155048
rect 355980 153190 356100 153218
rect 356072 151994 356100 153190
rect 356716 151994 356744 155110
rect 357176 154970 357204 159200
rect 358188 155582 358216 159200
rect 358176 155576 358228 155582
rect 358176 155518 358228 155524
rect 358820 155576 358872 155582
rect 358820 155518 358872 155524
rect 357440 155100 357492 155106
rect 357440 155042 357492 155048
rect 357164 154964 357216 154970
rect 357164 154906 357216 154912
rect 357452 151994 357480 155042
rect 357992 154964 358044 154970
rect 357992 154906 358044 154912
rect 358004 151994 358032 154906
rect 358832 151994 358860 155518
rect 359108 151994 359136 159200
rect 360120 154578 360148 159200
rect 360120 154550 360240 154578
rect 360212 151994 360240 154550
rect 361132 151994 361160 159200
rect 362052 154562 362080 159200
rect 363064 154562 363092 159200
rect 361488 154556 361540 154562
rect 361488 154498 361540 154504
rect 362040 154556 362092 154562
rect 362040 154498 362092 154504
rect 362592 154556 362644 154562
rect 362592 154498 362644 154504
rect 363052 154556 363104 154562
rect 363052 154498 363104 154504
rect 251416 151988 251712 151994
rect 251364 151982 251712 151988
rect 251376 151966 251712 151982
rect 252664 151966 253000 151994
rect 253308 151966 253644 151994
rect 253952 151966 254288 151994
rect 254596 151966 254932 151994
rect 255424 151966 255576 151994
rect 255884 151966 256220 151994
rect 256712 151966 256864 151994
rect 257172 151966 257508 151994
rect 258092 151966 258152 151994
rect 258460 151966 258796 151994
rect 259104 151966 259440 151994
rect 259840 151966 260176 151994
rect 260484 151966 260820 151994
rect 261128 151966 261464 151994
rect 261772 151966 262108 151994
rect 262416 151966 262752 151994
rect 263060 151966 263396 151994
rect 263704 151966 264040 151994
rect 264348 151966 264684 151994
rect 265084 151966 265328 151994
rect 265636 151966 265972 151994
rect 266372 151966 266616 151994
rect 266924 151966 267260 151994
rect 267844 151966 267904 151994
rect 268212 151966 268548 151994
rect 269132 151966 269284 151994
rect 269592 151966 269928 151994
rect 270512 151966 270572 151994
rect 270880 151966 271216 151994
rect 271524 151966 271860 151994
rect 272168 151966 272504 151994
rect 272812 151966 273148 151994
rect 273364 151966 273792 151994
rect 274100 151966 274436 151994
rect 274744 151966 275080 151994
rect 275388 151966 275724 151994
rect 276032 151966 276368 151994
rect 276676 151966 277012 151994
rect 277596 151966 277656 151994
rect 277964 151966 278300 151994
rect 278792 151966 279036 151994
rect 279344 151966 279680 151994
rect 280264 151966 280324 151994
rect 280632 151966 280968 151994
rect 281552 151966 281612 151994
rect 281920 151966 282256 151994
rect 282564 151966 282900 151994
rect 283208 151966 283544 151994
rect 283852 151966 284188 151994
rect 284496 151966 284832 151994
rect 285140 151966 285476 151994
rect 285784 151966 286120 151994
rect 286428 151966 286764 151994
rect 287256 151966 287408 151994
rect 287808 151966 288144 151994
rect 288452 151966 288788 151994
rect 289096 151966 289432 151994
rect 289832 151966 290076 151994
rect 290384 151966 290720 151994
rect 291212 151966 291364 151994
rect 291672 151966 292008 151994
rect 292592 151966 292652 151994
rect 292960 151966 293296 151994
rect 293604 151966 293940 151994
rect 294156 151966 294584 151994
rect 294892 151966 295228 151994
rect 295536 151966 295872 151994
rect 296180 151966 296516 151994
rect 297008 151966 297252 151994
rect 297560 151966 297896 151994
rect 298204 151966 298540 151994
rect 298848 151966 299184 151994
rect 299492 151966 299828 151994
rect 300136 151966 300472 151994
rect 300872 151966 301116 151994
rect 301424 151966 301760 151994
rect 302344 151966 302404 151994
rect 302712 151966 303048 151994
rect 303632 151966 303692 151994
rect 304000 151966 304336 151994
rect 304644 151966 304980 151994
rect 305288 151966 305624 151994
rect 305932 151966 306268 151994
rect 306668 151966 307004 151994
rect 307312 151966 307648 151994
rect 307956 151966 308292 151994
rect 308600 151966 308936 151994
rect 309244 151966 309580 151994
rect 309888 151966 310224 151994
rect 310532 151966 310868 151994
rect 311176 151966 311512 151994
rect 311912 151966 312156 151994
rect 312464 151966 312800 151994
rect 313292 151966 313444 151994
rect 313752 151966 314088 151994
rect 314672 151966 314732 151994
rect 315040 151966 315376 151994
rect 316052 151966 316112 151994
rect 316420 151966 316756 151994
rect 317064 151966 317400 151994
rect 317708 151966 318044 151994
rect 318352 151966 318688 151994
rect 318996 151966 319332 151994
rect 319640 151966 319976 151994
rect 320284 151966 320620 151994
rect 320928 151966 321264 151994
rect 321572 151966 321908 151994
rect 322216 151966 322552 151994
rect 322952 151966 323196 151994
rect 323504 151966 323840 151994
rect 324332 151966 324484 151994
rect 324884 151966 325220 151994
rect 325804 151966 325864 151994
rect 326172 151966 326508 151994
rect 327092 151966 327152 151994
rect 327460 151966 327796 151994
rect 328104 151966 328440 151994
rect 328656 151966 329084 151994
rect 329392 151966 329728 151994
rect 329944 151966 330372 151994
rect 330680 151966 331016 151994
rect 331324 151966 331660 151994
rect 331968 151966 332304 151994
rect 332612 151966 332948 151994
rect 333256 151966 333592 151994
rect 334176 151966 334328 151994
rect 334636 151966 334972 151994
rect 335464 151966 335616 151994
rect 335924 151966 336260 151994
rect 336752 151966 336904 151994
rect 337212 151966 337548 151994
rect 338132 151966 338192 151994
rect 338500 151966 338836 151994
rect 339144 151966 339480 151994
rect 339788 151966 340124 151994
rect 340432 151966 340768 151994
rect 341076 151966 341412 151994
rect 341720 151966 342056 151994
rect 342364 151966 342700 151994
rect 343008 151966 343344 151994
rect 343744 151966 344080 151994
rect 344388 151966 344724 151994
rect 345216 151966 345368 151994
rect 345676 151966 346012 151994
rect 346412 151966 346656 151994
rect 347056 151966 347300 151994
rect 347792 151966 347944 151994
rect 348252 151966 348588 151994
rect 349172 151966 349232 151994
rect 349540 151966 349876 151994
rect 350184 151966 350520 151994
rect 350828 151966 351164 151994
rect 351472 151966 351808 151994
rect 352116 151966 352452 151994
rect 352852 151966 353188 151994
rect 353496 151966 353832 151994
rect 354140 151966 354476 151994
rect 354876 151966 355120 151994
rect 355428 151966 355764 151994
rect 356072 151966 356408 151994
rect 356716 151966 357052 151994
rect 357452 151966 357696 151994
rect 358004 151966 358340 151994
rect 358832 151966 358984 151994
rect 359108 151966 359628 151994
rect 360212 151966 360272 151994
rect 360916 151966 361160 151994
rect 361500 151994 361528 154498
rect 362604 151994 362632 154498
rect 363984 154494 364012 159200
rect 362868 154488 362920 154494
rect 362868 154430 362920 154436
rect 363972 154488 364024 154494
rect 363972 154430 364024 154436
rect 361500 151966 361560 151994
rect 362296 151966 362632 151994
rect 362880 151994 362908 154430
rect 364156 153468 364208 153474
rect 364156 153410 364208 153416
rect 363880 153400 363932 153406
rect 363880 153342 363932 153348
rect 363892 151994 363920 153342
rect 362880 151966 362940 151994
rect 363584 151966 363920 151994
rect 249340 151914 249392 151920
rect 364168 151858 364196 153410
rect 364996 153406 365024 159200
rect 366008 155854 366036 159200
rect 365076 155848 365128 155854
rect 365076 155790 365128 155796
rect 365996 155848 366048 155854
rect 365996 155790 366048 155796
rect 365088 153474 365116 155790
rect 365628 154556 365680 154562
rect 365628 154498 365680 154504
rect 366456 154556 366508 154562
rect 366456 154498 366508 154504
rect 365076 153468 365128 153474
rect 365076 153410 365128 153416
rect 365168 153468 365220 153474
rect 365168 153410 365220 153416
rect 364984 153400 365036 153406
rect 364984 153342 365036 153348
rect 365180 151994 365208 153410
rect 365640 151994 365668 154498
rect 366468 151994 366496 154498
rect 366928 153474 366956 159200
rect 367940 154630 367968 159200
rect 368860 154630 368888 159200
rect 367928 154624 367980 154630
rect 367928 154566 367980 154572
rect 368848 154624 368900 154630
rect 368848 154566 368900 154572
rect 369872 154494 369900 159200
rect 370884 154630 370912 159200
rect 370872 154624 370924 154630
rect 370872 154566 370924 154572
rect 367008 154488 367060 154494
rect 367008 154430 367060 154436
rect 369860 154488 369912 154494
rect 369860 154430 369912 154436
rect 366916 153468 366968 153474
rect 366916 153410 366968 153416
rect 367020 151994 367048 154430
rect 367744 154420 367796 154426
rect 367744 154362 367796 154368
rect 367756 151994 367784 154362
rect 371804 154358 371832 159200
rect 368388 154352 368440 154358
rect 368388 154294 368440 154300
rect 371792 154352 371844 154358
rect 371792 154294 371844 154300
rect 368400 151994 368428 154294
rect 369676 154284 369728 154290
rect 369676 154226 369728 154232
rect 369032 153604 369084 153610
rect 369032 153546 369084 153552
rect 369044 151994 369072 153546
rect 369688 151994 369716 154226
rect 372344 154148 372396 154154
rect 372344 154090 372396 154096
rect 370964 153672 371016 153678
rect 370964 153614 371016 153620
rect 370320 153536 370372 153542
rect 370320 153478 370372 153484
rect 370332 151994 370360 153478
rect 370976 151994 371004 153614
rect 371608 153468 371660 153474
rect 371608 153410 371660 153416
rect 371620 151994 371648 153410
rect 372356 151994 372384 154090
rect 372816 153610 372844 159200
rect 373736 154290 373764 159200
rect 373724 154284 373776 154290
rect 373724 154226 373776 154232
rect 372988 154216 373040 154222
rect 372988 154158 373040 154164
rect 372804 153604 372856 153610
rect 372804 153546 372856 153552
rect 373000 151994 373028 154158
rect 373908 154012 373960 154018
rect 373908 153954 373960 153960
rect 373632 153876 373684 153882
rect 373632 153818 373684 153824
rect 373644 151994 373672 153818
rect 364872 151966 365208 151994
rect 365516 151966 365668 151994
rect 366160 151966 366496 151994
rect 366804 151966 367048 151994
rect 367448 151966 367784 151994
rect 368092 151966 368428 151994
rect 368736 151966 369072 151994
rect 369380 151966 369716 151994
rect 370024 151966 370360 151994
rect 370668 151966 371004 151994
rect 371312 151966 371648 151994
rect 372048 151966 372384 151994
rect 372692 151966 373028 151994
rect 373336 151966 373672 151994
rect 373920 151994 373948 153954
rect 374748 153542 374776 159200
rect 374920 154556 374972 154562
rect 374920 154498 374972 154504
rect 374736 153536 374788 153542
rect 374736 153478 374788 153484
rect 374932 151994 374960 154498
rect 375196 154488 375248 154494
rect 375196 154430 375248 154436
rect 373920 151966 373980 151994
rect 374624 151966 374960 151994
rect 375208 151994 375236 154430
rect 375760 153678 375788 159200
rect 376208 154420 376260 154426
rect 376208 154362 376260 154368
rect 375748 153672 375800 153678
rect 375748 153614 375800 153620
rect 376220 151994 376248 154362
rect 376484 153944 376536 153950
rect 376484 153886 376536 153892
rect 375208 151966 375268 151994
rect 375912 151966 376248 151994
rect 376496 151858 376524 153886
rect 376680 153474 376708 159200
rect 377692 154154 377720 159200
rect 378140 155508 378192 155514
rect 378140 155450 378192 155456
rect 377680 154148 377732 154154
rect 377680 154090 377732 154096
rect 378152 154018 378180 155450
rect 378612 154222 378640 159200
rect 379624 156618 379652 159200
rect 379532 156590 379652 156618
rect 379532 154578 379560 156590
rect 379612 155576 379664 155582
rect 379612 155518 379664 155524
rect 379440 154550 379560 154578
rect 378600 154216 378652 154222
rect 378600 154158 378652 154164
rect 378140 154012 378192 154018
rect 378140 153954 378192 153960
rect 379440 153882 379468 154550
rect 379624 154494 379652 155518
rect 380636 155514 380664 159200
rect 380900 155780 380952 155786
rect 380900 155722 380952 155728
rect 380624 155508 380676 155514
rect 380624 155450 380676 155456
rect 379612 154488 379664 154494
rect 379612 154430 379664 154436
rect 380912 153950 380940 155722
rect 381556 154630 381584 159200
rect 382568 155582 382596 159200
rect 382556 155576 382608 155582
rect 382556 155518 382608 155524
rect 382372 155508 382424 155514
rect 382372 155450 382424 155456
rect 382280 155372 382332 155378
rect 382280 155314 382332 155320
rect 381544 154624 381596 154630
rect 381544 154566 381596 154572
rect 381452 154284 381504 154290
rect 381452 154226 381504 154232
rect 380900 153944 380952 153950
rect 380900 153886 380952 153892
rect 379428 153876 379480 153882
rect 379428 153818 379480 153824
rect 377496 153808 377548 153814
rect 377496 153750 377548 153756
rect 376668 153468 376720 153474
rect 376668 153410 376720 153416
rect 377508 151994 377536 153750
rect 378784 153740 378836 153746
rect 378784 153682 378836 153688
rect 378048 153604 378100 153610
rect 378048 153546 378100 153552
rect 378060 151994 378088 153546
rect 378796 151994 378824 153682
rect 380072 153672 380124 153678
rect 380072 153614 380124 153620
rect 379428 153400 379480 153406
rect 379428 153342 379480 153348
rect 379440 151994 379468 153342
rect 380084 151994 380112 153614
rect 380716 153536 380768 153542
rect 380716 153478 380768 153484
rect 380728 151994 380756 153478
rect 381464 151994 381492 154226
rect 382096 154216 382148 154222
rect 382096 154158 382148 154164
rect 382108 151994 382136 154158
rect 382292 153610 382320 155314
rect 382384 153814 382412 155450
rect 383488 154630 383516 159200
rect 384500 155786 384528 159200
rect 384488 155780 384540 155786
rect 384488 155722 384540 155728
rect 385512 155514 385540 159200
rect 385868 155644 385920 155650
rect 385868 155586 385920 155592
rect 385500 155508 385552 155514
rect 385500 155450 385552 155456
rect 384856 155236 384908 155242
rect 384856 155178 384908 155184
rect 384212 154964 384264 154970
rect 384212 154906 384264 154912
rect 383476 154624 383528 154630
rect 383476 154566 383528 154572
rect 383292 154420 383344 154426
rect 383292 154362 383344 154368
rect 382740 153944 382792 153950
rect 382740 153886 382792 153892
rect 382372 153808 382424 153814
rect 382372 153750 382424 153756
rect 382280 153604 382332 153610
rect 382280 153546 382332 153552
rect 382752 151994 382780 153886
rect 383304 151994 383332 154362
rect 384028 154352 384080 154358
rect 384028 154294 384080 154300
rect 384040 151994 384068 154294
rect 384224 153746 384252 154906
rect 384212 153740 384264 153746
rect 384212 153682 384264 153688
rect 384672 153468 384724 153474
rect 384672 153410 384724 153416
rect 384684 151994 384712 153410
rect 384868 153406 384896 155178
rect 384948 154148 385000 154154
rect 384948 154090 385000 154096
rect 384856 153400 384908 153406
rect 384856 153342 384908 153348
rect 377200 151966 377536 151994
rect 377844 151966 378088 151994
rect 378488 151966 378824 151994
rect 379132 151966 379468 151994
rect 379776 151966 380112 151994
rect 380420 151966 380756 151994
rect 381156 151966 381492 151994
rect 381800 151966 382136 151994
rect 382444 151966 382780 151994
rect 383088 151966 383332 151994
rect 383732 151966 384068 151994
rect 384376 151966 384712 151994
rect 384960 151994 384988 154090
rect 385776 153808 385828 153814
rect 385776 153750 385828 153756
rect 385788 151994 385816 153750
rect 385880 153678 385908 155586
rect 385960 155576 386012 155582
rect 385960 155518 386012 155524
rect 385868 153672 385920 153678
rect 385868 153614 385920 153620
rect 385972 153542 386000 155518
rect 386432 155378 386460 159200
rect 386788 155508 386840 155514
rect 386788 155450 386840 155456
rect 386420 155372 386472 155378
rect 386420 155314 386472 155320
rect 386800 154290 386828 155450
rect 387444 154970 387472 159200
rect 388168 155916 388220 155922
rect 388168 155858 388220 155864
rect 387432 154964 387484 154970
rect 387432 154906 387484 154912
rect 387708 154556 387760 154562
rect 387708 154498 387760 154504
rect 386788 154284 386840 154290
rect 386788 154226 386840 154232
rect 386236 154080 386288 154086
rect 386236 154022 386288 154028
rect 385960 153536 386012 153542
rect 385960 153478 386012 153484
rect 384960 151966 385020 151994
rect 385664 151966 385816 151994
rect 386248 151858 386276 154022
rect 387248 153400 387300 153406
rect 387248 153342 387300 153348
rect 387260 151994 387288 153342
rect 387720 151994 387748 154498
rect 388180 153950 388208 155858
rect 388364 155242 388392 159200
rect 389376 155650 389404 159200
rect 389364 155644 389416 155650
rect 389364 155586 389416 155592
rect 390296 155582 390324 159200
rect 390284 155576 390336 155582
rect 390284 155518 390336 155524
rect 391308 155514 391336 159200
rect 391296 155508 391348 155514
rect 391296 155450 391348 155456
rect 388352 155236 388404 155242
rect 388352 155178 388404 155184
rect 390468 154488 390520 154494
rect 390468 154430 390520 154436
rect 389824 154012 389876 154018
rect 389824 153954 389876 153960
rect 388168 153944 388220 153950
rect 388168 153886 388220 153892
rect 389088 153876 389140 153882
rect 389088 153818 389140 153824
rect 388536 153672 388588 153678
rect 388536 153614 388588 153620
rect 388548 151994 388576 153614
rect 389100 151994 389128 153818
rect 389836 151994 389864 153954
rect 390480 151994 390508 154430
rect 392320 154222 392348 159200
rect 393240 155922 393268 159200
rect 393228 155916 393280 155922
rect 393228 155858 393280 155864
rect 394252 154426 394280 159200
rect 394240 154420 394292 154426
rect 394240 154362 394292 154368
rect 395068 154420 395120 154426
rect 395068 154362 395120 154368
rect 393044 154284 393096 154290
rect 393044 154226 393096 154232
rect 392308 154216 392360 154222
rect 392308 154158 392360 154164
rect 391204 153944 391256 153950
rect 391204 153886 391256 153892
rect 391216 151994 391244 153886
rect 391848 153740 391900 153746
rect 391848 153682 391900 153688
rect 391860 151994 391888 153682
rect 392492 153536 392544 153542
rect 392492 153478 392544 153484
rect 392504 151994 392532 153478
rect 393056 151994 393084 154226
rect 394424 154216 394476 154222
rect 394424 154158 394476 154164
rect 393780 153604 393832 153610
rect 393780 153546 393832 153552
rect 393792 151994 393820 153546
rect 394436 151994 394464 154158
rect 395080 151994 395108 154362
rect 395172 154358 395200 159200
rect 395988 154828 396040 154834
rect 395988 154770 396040 154776
rect 395160 154352 395212 154358
rect 395160 154294 395212 154300
rect 395712 154216 395764 154222
rect 395712 154158 395764 154164
rect 395724 151994 395752 154158
rect 386952 151966 387288 151994
rect 387596 151966 387748 151994
rect 388240 151966 388576 151994
rect 388884 151966 389128 151994
rect 389528 151966 389864 151994
rect 390264 151966 390508 151994
rect 390908 151966 391244 151994
rect 391552 151966 391888 151994
rect 392196 151966 392532 151994
rect 392840 151966 393084 151994
rect 393484 151966 393820 151994
rect 394128 151966 394464 151994
rect 394772 151966 395108 151994
rect 395416 151966 395752 151994
rect 396000 151994 396028 154770
rect 396184 153474 396212 159200
rect 397196 154154 397224 159200
rect 397184 154148 397236 154154
rect 397184 154090 397236 154096
rect 397276 154148 397328 154154
rect 397276 154090 397328 154096
rect 396172 153468 396224 153474
rect 396172 153410 396224 153416
rect 397000 153468 397052 153474
rect 397000 153410 397052 153416
rect 397012 151994 397040 153410
rect 396000 151966 396060 151994
rect 396704 151966 397040 151994
rect 397288 151994 397316 154090
rect 398116 153814 398144 159200
rect 398564 155440 398616 155446
rect 398564 155382 398616 155388
rect 398104 153808 398156 153814
rect 398104 153750 398156 153756
rect 398288 153808 398340 153814
rect 398288 153750 398340 153756
rect 398300 151994 398328 153750
rect 397288 151966 397348 151994
rect 397992 151966 398328 151994
rect 398576 151858 398604 155382
rect 398852 154578 398880 159310
rect 399036 159202 399064 159310
rect 399114 159202 399170 160000
rect 399036 159200 399170 159202
rect 400034 159200 400090 160000
rect 401046 159200 401102 160000
rect 402058 159200 402114 160000
rect 402978 159200 403034 160000
rect 403990 159200 404046 160000
rect 404910 159200 404966 160000
rect 405922 159200 405978 160000
rect 406934 159200 406990 160000
rect 407854 159200 407910 160000
rect 408866 159200 408922 160000
rect 409786 159200 409842 160000
rect 410798 159200 410854 160000
rect 411810 159200 411866 160000
rect 412730 159200 412786 160000
rect 413742 159200 413798 160000
rect 414662 159200 414718 160000
rect 415674 159200 415730 160000
rect 416686 159200 416742 160000
rect 417606 159200 417662 160000
rect 418618 159200 418674 160000
rect 419538 159200 419594 160000
rect 420550 159200 420606 160000
rect 421562 159200 421618 160000
rect 422482 159200 422538 160000
rect 423494 159200 423550 160000
rect 424414 159200 424470 160000
rect 425426 159200 425482 160000
rect 426346 159200 426402 160000
rect 427358 159200 427414 160000
rect 428370 159200 428426 160000
rect 429290 159200 429346 160000
rect 430302 159200 430358 160000
rect 431222 159200 431278 160000
rect 432234 159200 432290 160000
rect 433246 159200 433302 160000
rect 434166 159200 434222 160000
rect 435178 159200 435234 160000
rect 436098 159200 436154 160000
rect 437110 159200 437166 160000
rect 438122 159200 438178 160000
rect 439042 159200 439098 160000
rect 440054 159200 440110 160000
rect 440974 159200 441030 160000
rect 441986 159200 442042 160000
rect 442998 159200 443054 160000
rect 443918 159200 443974 160000
rect 444930 159200 444986 160000
rect 445850 159200 445906 160000
rect 446862 159200 446918 160000
rect 447874 159200 447930 160000
rect 448794 159200 448850 160000
rect 449806 159200 449862 160000
rect 450726 159200 450782 160000
rect 451738 159200 451794 160000
rect 452750 159200 452806 160000
rect 453670 159200 453726 160000
rect 454682 159200 454738 160000
rect 455602 159200 455658 160000
rect 456614 159200 456670 160000
rect 457626 159200 457682 160000
rect 458546 159200 458602 160000
rect 459558 159200 459614 160000
rect 460478 159200 460534 160000
rect 461490 159200 461546 160000
rect 462502 159200 462558 160000
rect 463422 159200 463478 160000
rect 464434 159200 464490 160000
rect 465354 159200 465410 160000
rect 466366 159200 466422 160000
rect 467286 159200 467342 160000
rect 468298 159200 468354 160000
rect 469310 159200 469366 160000
rect 470230 159200 470286 160000
rect 471242 159200 471298 160000
rect 472162 159200 472218 160000
rect 473174 159200 473230 160000
rect 474186 159200 474242 160000
rect 475106 159200 475162 160000
rect 476118 159200 476174 160000
rect 477038 159200 477094 160000
rect 478050 159200 478106 160000
rect 479062 159200 479118 160000
rect 479982 159200 480038 160000
rect 480994 159200 481050 160000
rect 481914 159200 481970 160000
rect 482926 159200 482982 160000
rect 483938 159200 483994 160000
rect 484858 159200 484914 160000
rect 485870 159200 485926 160000
rect 486790 159200 486846 160000
rect 487802 159200 487858 160000
rect 488814 159200 488870 160000
rect 489734 159200 489790 160000
rect 490746 159200 490802 160000
rect 491666 159200 491722 160000
rect 492678 159200 492734 160000
rect 493690 159200 493746 160000
rect 494610 159200 494666 160000
rect 495622 159200 495678 160000
rect 496542 159200 496598 160000
rect 497554 159200 497610 160000
rect 498566 159200 498622 160000
rect 499486 159200 499542 160000
rect 500498 159200 500554 160000
rect 501418 159200 501474 160000
rect 502430 159200 502486 160000
rect 503350 159200 503406 160000
rect 504362 159200 504418 160000
rect 505374 159200 505430 160000
rect 506294 159200 506350 160000
rect 507306 159200 507362 160000
rect 508226 159200 508282 160000
rect 509238 159200 509294 160000
rect 510250 159200 510306 160000
rect 511170 159200 511226 160000
rect 512182 159200 512238 160000
rect 513102 159200 513158 160000
rect 514114 159200 514170 160000
rect 515126 159200 515182 160000
rect 516046 159200 516102 160000
rect 517058 159200 517114 160000
rect 517978 159200 518034 160000
rect 518990 159200 519046 160000
rect 520002 159200 520058 160000
rect 520922 159200 520978 160000
rect 521934 159200 521990 160000
rect 522854 159200 522910 160000
rect 523866 159200 523922 160000
rect 524878 159200 524934 160000
rect 525798 159200 525854 160000
rect 526810 159200 526866 160000
rect 527730 159200 527786 160000
rect 528742 159200 528798 160000
rect 529754 159200 529810 160000
rect 530674 159200 530730 160000
rect 531686 159200 531742 160000
rect 532606 159200 532662 160000
rect 533618 159200 533674 160000
rect 534630 159200 534686 160000
rect 535550 159200 535606 160000
rect 536562 159200 536618 160000
rect 537482 159200 537538 160000
rect 538494 159200 538550 160000
rect 539506 159200 539562 160000
rect 540426 159200 540482 160000
rect 541438 159200 541494 160000
rect 542358 159200 542414 160000
rect 543370 159200 543426 160000
rect 544290 159200 544346 160000
rect 545302 159200 545358 160000
rect 546314 159200 546370 160000
rect 547234 159200 547290 160000
rect 548246 159200 548302 160000
rect 549166 159200 549222 160000
rect 550178 159200 550234 160000
rect 551190 159200 551246 160000
rect 552110 159200 552166 160000
rect 553122 159200 553178 160000
rect 554042 159200 554098 160000
rect 555054 159200 555110 160000
rect 556066 159200 556122 160000
rect 556986 159200 557042 160000
rect 557998 159200 558054 160000
rect 558918 159200 558974 160000
rect 559930 159200 559986 160000
rect 560942 159200 560998 160000
rect 561862 159200 561918 160000
rect 562874 159200 562930 160000
rect 563794 159200 563850 160000
rect 564806 159200 564862 160000
rect 565818 159200 565874 160000
rect 566738 159200 566794 160000
rect 567750 159200 567806 160000
rect 568670 159200 568726 160000
rect 569682 159200 569738 160000
rect 570694 159200 570750 160000
rect 571614 159200 571670 160000
rect 572626 159200 572682 160000
rect 573546 159200 573602 160000
rect 574558 159200 574614 160000
rect 575570 159200 575626 160000
rect 576490 159200 576546 160000
rect 576872 159310 577452 159338
rect 399036 159174 399156 159200
rect 399576 155032 399628 155038
rect 399576 154974 399628 154980
rect 398760 154550 398880 154578
rect 398760 154086 398788 154550
rect 398748 154080 398800 154086
rect 398748 154022 398800 154028
rect 399588 151994 399616 154974
rect 400048 153406 400076 159200
rect 400312 155100 400364 155106
rect 400312 155042 400364 155048
rect 400220 154964 400272 154970
rect 400220 154906 400272 154912
rect 400128 154080 400180 154086
rect 400128 154022 400180 154028
rect 400036 153400 400088 153406
rect 400036 153342 400088 153348
rect 400140 151994 400168 154022
rect 400232 153882 400260 154906
rect 400220 153876 400272 153882
rect 400220 153818 400272 153824
rect 400324 153678 400352 155042
rect 400956 154896 401008 154902
rect 400956 154838 401008 154844
rect 400312 153672 400364 153678
rect 400312 153614 400364 153620
rect 400968 151994 400996 154838
rect 401060 154630 401088 159200
rect 401692 155916 401744 155922
rect 401692 155858 401744 155864
rect 401600 155372 401652 155378
rect 401600 155314 401652 155320
rect 401508 155236 401560 155242
rect 401508 155178 401560 155184
rect 401048 154624 401100 154630
rect 401048 154566 401100 154572
rect 401520 151994 401548 155178
rect 401612 154494 401640 155314
rect 401600 154488 401652 154494
rect 401600 154430 401652 154436
rect 401704 154018 401732 155858
rect 402072 155106 402100 159200
rect 402244 155304 402296 155310
rect 402244 155246 402296 155252
rect 402060 155100 402112 155106
rect 402060 155042 402112 155048
rect 401692 154012 401744 154018
rect 401692 153954 401744 153960
rect 402256 151994 402284 155246
rect 402992 154970 403020 159200
rect 404004 155922 404032 159200
rect 403992 155916 404044 155922
rect 403992 155858 404044 155864
rect 404820 155916 404872 155922
rect 404820 155858 404872 155864
rect 403440 155848 403492 155854
rect 403440 155790 403492 155796
rect 402980 154964 403032 154970
rect 402980 154906 403032 154912
rect 402704 153876 402756 153882
rect 402704 153818 402756 153824
rect 402716 151994 402744 153818
rect 403452 153746 403480 155790
rect 404176 155712 404228 155718
rect 404176 155654 404228 155660
rect 403440 153740 403492 153746
rect 403440 153682 403492 153688
rect 403532 153672 403584 153678
rect 403532 153614 403584 153620
rect 403544 151994 403572 153614
rect 404188 151994 404216 155654
rect 404268 155508 404320 155514
rect 404268 155450 404320 155456
rect 404280 153950 404308 155450
rect 404728 154964 404780 154970
rect 404728 154906 404780 154912
rect 404268 153944 404320 153950
rect 404268 153886 404320 153892
rect 404740 151994 404768 154906
rect 404832 153542 404860 155858
rect 404924 155378 404952 159200
rect 405936 155514 405964 159200
rect 406948 155854 406976 159200
rect 407868 155922 407896 159200
rect 407856 155916 407908 155922
rect 407856 155858 407908 155864
rect 406936 155848 406988 155854
rect 406936 155790 406988 155796
rect 406108 155644 406160 155650
rect 406108 155586 406160 155592
rect 405924 155508 405976 155514
rect 405924 155450 405976 155456
rect 404912 155372 404964 155378
rect 404912 155314 404964 155320
rect 405924 155168 405976 155174
rect 405924 155110 405976 155116
rect 405464 154012 405516 154018
rect 405464 153954 405516 153960
rect 404820 153536 404872 153542
rect 404820 153478 404872 153484
rect 405476 151994 405504 153954
rect 405936 153610 405964 155110
rect 405924 153604 405976 153610
rect 405924 153546 405976 153552
rect 406120 151994 406148 155586
rect 407764 155508 407816 155514
rect 407764 155450 407816 155456
rect 407028 154828 407080 154834
rect 407028 154770 407080 154776
rect 406752 154760 406804 154766
rect 406752 154702 406804 154708
rect 406764 151994 406792 154702
rect 399280 151966 399616 151994
rect 400016 151966 400168 151994
rect 400660 151966 400996 151994
rect 401304 151966 401548 151994
rect 401948 151966 402284 151994
rect 402592 151966 402744 151994
rect 403236 151966 403572 151994
rect 403880 151966 404216 151994
rect 404524 151966 404768 151994
rect 405168 151966 405504 151994
rect 405812 151966 406148 151994
rect 406456 151966 406792 151994
rect 407040 151994 407068 154770
rect 407776 153474 407804 155450
rect 408316 154488 408368 154494
rect 408316 154430 408368 154436
rect 408040 153944 408092 153950
rect 408040 153886 408092 153892
rect 407764 153468 407816 153474
rect 407764 153410 407816 153416
rect 408052 151994 408080 153886
rect 407040 151966 407100 151994
rect 407744 151966 408080 151994
rect 408328 151858 408356 154430
rect 408880 154290 408908 159200
rect 409696 155712 409748 155718
rect 409696 155654 409748 155660
rect 409420 154692 409472 154698
rect 409420 154634 409472 154640
rect 408868 154284 408920 154290
rect 408868 154226 408920 154232
rect 409432 151994 409460 154634
rect 409124 151966 409460 151994
rect 409708 151994 409736 155654
rect 409800 155174 409828 159200
rect 409788 155168 409840 155174
rect 409788 155110 409840 155116
rect 410708 154556 410760 154562
rect 410708 154498 410760 154504
rect 410720 151994 410748 154498
rect 410812 154426 410840 159200
rect 411168 155440 411220 155446
rect 411168 155382 411220 155388
rect 410800 154420 410852 154426
rect 410800 154362 410852 154368
rect 411180 151994 411208 155382
rect 411824 154358 411852 159200
rect 412548 155916 412600 155922
rect 412548 155858 412600 155864
rect 412640 155916 412692 155922
rect 412744 155904 412772 159200
rect 412692 155876 412772 155904
rect 412640 155858 412692 155864
rect 411996 155576 412048 155582
rect 411996 155518 412048 155524
rect 411812 154352 411864 154358
rect 411812 154294 411864 154300
rect 412008 151994 412036 155518
rect 412456 155508 412508 155514
rect 412456 155450 412508 155456
rect 412468 151994 412496 155450
rect 412560 154222 412588 155858
rect 413756 155038 413784 159200
rect 414676 155786 414704 159200
rect 414664 155780 414716 155786
rect 414664 155722 414716 155728
rect 413836 155576 413888 155582
rect 413836 155518 413888 155524
rect 413744 155032 413796 155038
rect 413744 154974 413796 154980
rect 413652 154964 413704 154970
rect 413652 154906 413704 154912
rect 413284 154352 413336 154358
rect 413284 154294 413336 154300
rect 412548 154216 412600 154222
rect 412548 154158 412600 154164
rect 413296 151994 413324 154294
rect 413664 153678 413692 154906
rect 413848 153814 413876 155518
rect 415216 154964 415268 154970
rect 415216 154906 415268 154912
rect 414572 154624 414624 154630
rect 414572 154566 414624 154572
rect 413928 154420 413980 154426
rect 413928 154362 413980 154368
rect 413836 153808 413888 153814
rect 413836 153750 413888 153756
rect 413652 153672 413704 153678
rect 413652 153614 413704 153620
rect 413940 151994 413968 154362
rect 414584 151994 414612 154566
rect 415228 151994 415256 154906
rect 415688 154154 415716 159200
rect 415860 156664 415912 156670
rect 415860 156606 415912 156612
rect 415676 154148 415728 154154
rect 415676 154090 415728 154096
rect 415872 151994 415900 156606
rect 416700 155582 416728 159200
rect 416688 155576 416740 155582
rect 416688 155518 416740 155524
rect 417620 155378 417648 159200
rect 417608 155372 417660 155378
rect 417608 155314 417660 155320
rect 417976 155372 418028 155378
rect 417976 155314 418028 155320
rect 417792 154760 417844 154766
rect 417792 154702 417844 154708
rect 416504 153808 416556 153814
rect 416504 153750 416556 153756
rect 416516 151994 416544 153750
rect 417148 153604 417200 153610
rect 417148 153546 417200 153552
rect 417160 151994 417188 153546
rect 417804 151994 417832 154702
rect 417988 153610 418016 155314
rect 418632 155106 418660 159200
rect 418620 155100 418672 155106
rect 418620 155042 418672 155048
rect 419448 155032 419500 155038
rect 419448 154974 419500 154980
rect 419172 154216 419224 154222
rect 419172 154158 419224 154164
rect 417976 153604 418028 153610
rect 417976 153546 418028 153552
rect 418528 152516 418580 152522
rect 418528 152458 418580 152464
rect 418540 151994 418568 152458
rect 419184 151994 419212 154158
rect 409708 151966 409768 151994
rect 410412 151966 410748 151994
rect 411056 151966 411208 151994
rect 411700 151966 412036 151994
rect 412344 151966 412496 151994
rect 412988 151966 413324 151994
rect 413632 151966 413968 151994
rect 414276 151966 414612 151994
rect 414920 151966 415256 151994
rect 415564 151966 415900 151994
rect 416208 151966 416544 151994
rect 416852 151966 417188 151994
rect 417496 151966 417832 151994
rect 418232 151966 418568 151994
rect 418876 151966 419212 151994
rect 419460 151994 419488 154974
rect 419552 154086 419580 159200
rect 420564 154902 420592 159200
rect 420736 156596 420788 156602
rect 420736 156538 420788 156544
rect 420552 154896 420604 154902
rect 420552 154838 420604 154844
rect 420460 154828 420512 154834
rect 420460 154770 420512 154776
rect 419540 154080 419592 154086
rect 419540 154022 419592 154028
rect 420472 151994 420500 154770
rect 419460 151966 419520 151994
rect 420164 151966 420500 151994
rect 420748 151858 420776 156538
rect 421576 155242 421604 159200
rect 422496 155310 422524 159200
rect 422484 155304 422536 155310
rect 422484 155246 422536 155252
rect 421564 155236 421616 155242
rect 421564 155178 421616 155184
rect 422024 155236 422076 155242
rect 422024 155178 422076 155184
rect 421748 154148 421800 154154
rect 421748 154090 421800 154096
rect 421760 151994 421788 154090
rect 421452 151966 421788 151994
rect 422036 151994 422064 155178
rect 423036 154964 423088 154970
rect 423036 154906 423088 154912
rect 423048 151994 423076 154906
rect 423508 153882 423536 159200
rect 424428 155106 424456 159200
rect 425440 155854 425468 159200
rect 426256 157344 426308 157350
rect 426256 157286 426308 157292
rect 425428 155848 425480 155854
rect 425428 155790 425480 155796
rect 424968 155304 425020 155310
rect 424968 155246 425020 155252
rect 424416 155100 424468 155106
rect 424416 155042 424468 155048
rect 423496 153876 423548 153882
rect 423496 153818 423548 153824
rect 424324 153740 424376 153746
rect 424324 153682 424376 153688
rect 423588 153128 423640 153134
rect 423588 153070 423640 153076
rect 423600 151994 423628 153070
rect 424336 151994 424364 153682
rect 424980 151994 425008 155246
rect 425612 155100 425664 155106
rect 425612 155042 425664 155048
rect 425624 151994 425652 155042
rect 426268 151994 426296 157286
rect 426360 155174 426388 159200
rect 426348 155168 426400 155174
rect 426348 155110 426400 155116
rect 426900 154080 426952 154086
rect 426900 154022 426952 154028
rect 426912 151994 426940 154022
rect 427372 154018 427400 159200
rect 428384 155922 428412 159200
rect 428924 157276 428976 157282
rect 428924 157218 428976 157224
rect 428372 155916 428424 155922
rect 428372 155858 428424 155864
rect 427636 155848 427688 155854
rect 427636 155790 427688 155796
rect 427360 154012 427412 154018
rect 427360 153954 427412 153960
rect 427648 151994 427676 155790
rect 428280 155168 428332 155174
rect 428280 155110 428332 155116
rect 428292 151994 428320 155110
rect 428936 151994 428964 157218
rect 429304 155786 429332 159200
rect 430212 155916 430264 155922
rect 430212 155858 430264 155864
rect 429292 155780 429344 155786
rect 429292 155722 429344 155728
rect 429568 154012 429620 154018
rect 429568 153954 429620 153960
rect 429580 151994 429608 153954
rect 430224 151994 430252 155858
rect 430316 155582 430344 159200
rect 430488 155780 430540 155786
rect 430488 155722 430540 155728
rect 430304 155576 430356 155582
rect 430304 155518 430356 155524
rect 422036 151966 422096 151994
rect 422740 151966 423076 151994
rect 423384 151966 423628 151994
rect 424028 151966 424364 151994
rect 424672 151966 425008 151994
rect 425316 151966 425652 151994
rect 425960 151966 426296 151994
rect 426604 151966 426940 151994
rect 427340 151966 427676 151994
rect 427984 151966 428320 151994
rect 428628 151966 428964 151994
rect 429272 151966 429608 151994
rect 429916 151966 430252 151994
rect 430500 151994 430528 155722
rect 431236 153950 431264 159200
rect 432248 154494 432276 159200
rect 433064 155576 433116 155582
rect 433064 155518 433116 155524
rect 432236 154488 432288 154494
rect 432236 154430 432288 154436
rect 432604 154488 432656 154494
rect 432604 154430 432656 154436
rect 431224 153944 431276 153950
rect 431224 153886 431276 153892
rect 431776 153944 431828 153950
rect 431776 153886 431828 153892
rect 431500 153060 431552 153066
rect 431500 153002 431552 153008
rect 431512 151994 431540 153002
rect 430500 151966 430560 151994
rect 431204 151966 431540 151994
rect 431788 151858 431816 153886
rect 432616 151994 432644 154430
rect 432492 151966 432644 151994
rect 433076 151858 433104 155518
rect 433260 154698 433288 159200
rect 434180 155718 434208 159200
rect 434628 157140 434680 157146
rect 434628 157082 434680 157088
rect 434168 155712 434220 155718
rect 434168 155654 434220 155660
rect 433248 154692 433300 154698
rect 433248 154634 433300 154640
rect 434076 152992 434128 152998
rect 434076 152934 434128 152940
rect 434088 151994 434116 152934
rect 434640 151994 434668 157082
rect 435192 154562 435220 159200
rect 435364 155712 435416 155718
rect 435364 155654 435416 155660
rect 435180 154556 435232 154562
rect 435180 154498 435232 154504
rect 435376 151994 435404 155654
rect 436112 155446 436140 159200
rect 436652 157072 436704 157078
rect 436652 157014 436704 157020
rect 436100 155440 436152 155446
rect 436100 155382 436152 155388
rect 436006 155272 436062 155281
rect 436006 155207 436062 155216
rect 436020 151994 436048 155207
rect 436664 151994 436692 157014
rect 437124 155650 437152 159200
rect 437388 157004 437440 157010
rect 437388 156946 437440 156952
rect 437112 155644 437164 155650
rect 437112 155586 437164 155592
rect 437400 151994 437428 156946
rect 438136 155514 438164 159200
rect 438676 155644 438728 155650
rect 438676 155586 438728 155592
rect 438124 155508 438176 155514
rect 438124 155450 438176 155456
rect 438032 155440 438084 155446
rect 438032 155382 438084 155388
rect 438044 151994 438072 155382
rect 438688 151994 438716 155586
rect 439056 154358 439084 159200
rect 439964 156936 440016 156942
rect 439964 156878 440016 156884
rect 439044 154352 439096 154358
rect 439044 154294 439096 154300
rect 439320 152924 439372 152930
rect 439320 152866 439372 152872
rect 439332 151994 439360 152866
rect 439976 151994 440004 156878
rect 440068 154426 440096 159200
rect 440988 154630 441016 159200
rect 441528 156868 441580 156874
rect 441528 156810 441580 156816
rect 441252 155440 441304 155446
rect 441252 155382 441304 155388
rect 440976 154624 441028 154630
rect 440976 154566 441028 154572
rect 440056 154420 440108 154426
rect 440056 154362 440108 154368
rect 440608 152856 440660 152862
rect 440608 152798 440660 152804
rect 440620 151994 440648 152798
rect 441264 151994 441292 155382
rect 433780 151966 434116 151994
rect 434424 151966 434668 151994
rect 435068 151966 435404 151994
rect 435712 151966 436048 151994
rect 436356 151966 436692 151994
rect 437092 151966 437428 151994
rect 437736 151966 438072 151994
rect 438380 151966 438716 151994
rect 439024 151966 439360 151994
rect 439668 151966 440004 151994
rect 440312 151966 440648 151994
rect 440956 151966 441292 151994
rect 441540 151994 441568 156810
rect 442000 154766 442028 159200
rect 442540 157208 442592 157214
rect 442540 157150 442592 157156
rect 441988 154760 442040 154766
rect 441988 154702 442040 154708
rect 442552 151994 442580 157150
rect 442816 156800 442868 156806
rect 442816 156742 442868 156748
rect 441540 151966 441600 151994
rect 442244 151966 442580 151994
rect 442828 151858 442856 156742
rect 443012 156670 443040 159200
rect 443000 156664 443052 156670
rect 443000 156606 443052 156612
rect 443932 153814 443960 159200
rect 444944 155378 444972 159200
rect 445116 156052 445168 156058
rect 445116 155994 445168 156000
rect 444932 155372 444984 155378
rect 444932 155314 444984 155320
rect 443920 153808 443972 153814
rect 443920 153750 443972 153756
rect 443828 153604 443880 153610
rect 443828 153546 443880 153552
rect 443840 151994 443868 153546
rect 445128 151994 445156 155994
rect 445668 155372 445720 155378
rect 445668 155314 445720 155320
rect 445680 153610 445708 155314
rect 445864 154834 445892 159200
rect 445852 154828 445904 154834
rect 445852 154770 445904 154776
rect 445668 153604 445720 153610
rect 445668 153546 445720 153552
rect 445668 152720 445720 152726
rect 445668 152662 445720 152668
rect 445680 151994 445708 152662
rect 446496 152652 446548 152658
rect 446496 152594 446548 152600
rect 446508 151994 446536 152594
rect 446876 152522 446904 159200
rect 447048 156732 447100 156738
rect 447048 156674 447100 156680
rect 446864 152516 446916 152522
rect 446864 152458 446916 152464
rect 447060 151994 447088 156674
rect 447888 154222 447916 159200
rect 448428 156664 448480 156670
rect 448428 156606 448480 156612
rect 447876 154216 447928 154222
rect 447876 154158 447928 154164
rect 447784 152040 447836 152046
rect 443532 151966 443868 151994
rect 444176 151978 444328 151994
rect 444176 151972 444340 151978
rect 444176 151966 444288 151972
rect 444820 151966 445156 151994
rect 445464 151966 445708 151994
rect 446200 151966 446536 151994
rect 446844 151966 447088 151994
rect 447488 151988 447784 151994
rect 448440 151994 448468 156606
rect 448808 155038 448836 159200
rect 449072 156256 449124 156262
rect 449072 156198 449124 156204
rect 448796 155032 448848 155038
rect 448796 154974 448848 154980
rect 449084 151994 449112 156198
rect 449820 154902 449848 159200
rect 450740 156602 450768 159200
rect 450728 156596 450780 156602
rect 450728 156538 450780 156544
rect 450360 156120 450412 156126
rect 450360 156062 450412 156068
rect 449808 154896 449860 154902
rect 449808 154838 449860 154844
rect 449716 152584 449768 152590
rect 449716 152526 449768 152532
rect 449728 151994 449756 152526
rect 450372 151994 450400 156062
rect 451752 154154 451780 159200
rect 452568 156324 452620 156330
rect 452568 156266 452620 156272
rect 451740 154148 451792 154154
rect 451740 154090 451792 154096
rect 452292 152516 452344 152522
rect 452292 152458 452344 152464
rect 450682 152176 450734 152182
rect 450682 152118 450734 152124
rect 447488 151982 447836 151988
rect 447488 151966 447824 151982
rect 448132 151966 448468 151994
rect 448776 151966 449112 151994
rect 449420 151966 449756 151994
rect 450064 151966 450400 151994
rect 450694 151980 450722 152118
rect 451326 152108 451378 152114
rect 451326 152050 451378 152056
rect 451338 151980 451366 152050
rect 452304 151994 452332 152458
rect 451996 151966 452332 151994
rect 452580 151994 452608 156266
rect 452764 155242 452792 159200
rect 453580 156188 453632 156194
rect 453580 156130 453632 156136
rect 452752 155236 452804 155242
rect 452752 155178 452804 155184
rect 453592 151994 453620 156130
rect 453684 154970 453712 159200
rect 453672 154964 453724 154970
rect 453672 154906 453724 154912
rect 454696 153134 454724 159200
rect 454868 155236 454920 155242
rect 454868 155178 454920 155184
rect 454684 153128 454736 153134
rect 454684 153070 454736 153076
rect 453902 152244 453954 152250
rect 453902 152186 453954 152192
rect 452580 151966 452640 151994
rect 453284 151966 453620 151994
rect 453914 151980 453942 152186
rect 454880 151994 454908 155178
rect 455616 153746 455644 159200
rect 456524 156392 456576 156398
rect 456524 156334 456576 156340
rect 456248 153876 456300 153882
rect 456248 153818 456300 153824
rect 455604 153740 455656 153746
rect 455604 153682 455656 153688
rect 455236 153604 455288 153610
rect 455236 153546 455288 153552
rect 454572 151966 454908 151994
rect 444288 151914 444340 151920
rect 455248 151858 455276 153546
rect 456260 151994 456288 153818
rect 455952 151966 456288 151994
rect 456536 151994 456564 156334
rect 456628 155310 456656 159200
rect 456616 155304 456668 155310
rect 456616 155246 456668 155252
rect 456708 155304 456760 155310
rect 456708 155246 456760 155252
rect 456720 153610 456748 155246
rect 457640 155106 457668 159200
rect 458560 157350 458588 159200
rect 458548 157344 458600 157350
rect 458548 157286 458600 157292
rect 457628 155100 457680 155106
rect 457628 155042 457680 155048
rect 459468 154896 459520 154902
rect 459468 154838 459520 154844
rect 457536 154760 457588 154766
rect 457536 154702 457588 154708
rect 456708 153604 456760 153610
rect 456708 153546 456760 153552
rect 457548 151994 457576 154702
rect 458088 153536 458140 153542
rect 458088 153478 458140 153484
rect 458100 151994 458128 153478
rect 458824 152312 458876 152318
rect 458824 152254 458876 152260
rect 458836 151994 458864 152254
rect 459480 151994 459508 154838
rect 459572 154086 459600 159200
rect 460492 155854 460520 159200
rect 460480 155848 460532 155854
rect 460480 155790 460532 155796
rect 461504 155038 461532 159200
rect 462516 157282 462544 159200
rect 462504 157276 462556 157282
rect 462504 157218 462556 157224
rect 462688 156460 462740 156466
rect 462688 156402 462740 156408
rect 461492 155032 461544 155038
rect 461492 154974 461544 154980
rect 462044 155032 462096 155038
rect 462044 154974 462096 154980
rect 460112 154964 460164 154970
rect 460112 154906 460164 154912
rect 459560 154080 459612 154086
rect 459560 154022 459612 154028
rect 460124 151994 460152 154906
rect 460664 154828 460716 154834
rect 460664 154770 460716 154776
rect 460676 151994 460704 154770
rect 461400 154556 461452 154562
rect 461400 154498 461452 154504
rect 461412 151994 461440 154498
rect 462056 151994 462084 154974
rect 462700 151994 462728 156402
rect 463332 155100 463384 155106
rect 463332 155042 463384 155048
rect 463344 151994 463372 155042
rect 463436 154018 463464 159200
rect 464448 155922 464476 159200
rect 464436 155916 464488 155922
rect 464436 155858 464488 155864
rect 464988 155916 465040 155922
rect 464988 155858 465040 155864
rect 464620 155168 464672 155174
rect 464620 155110 464672 155116
rect 463424 154012 463476 154018
rect 463424 153954 463476 153960
rect 463608 153604 463660 153610
rect 463608 153546 463660 153552
rect 456536 151966 456596 151994
rect 457240 151966 457576 151994
rect 457884 151966 458128 151994
rect 458528 151966 458864 151994
rect 459172 151966 459508 151994
rect 459816 151966 460152 151994
rect 460460 151966 460704 151994
rect 461104 151966 461440 151994
rect 461748 151966 462084 151994
rect 462392 151966 462728 151994
rect 463036 151966 463372 151994
rect 463620 151994 463648 153546
rect 464632 151994 464660 155110
rect 463620 151966 463680 151994
rect 464324 151966 464660 151994
rect 465000 151994 465028 155858
rect 465368 155786 465396 159200
rect 465356 155780 465408 155786
rect 465356 155722 465408 155728
rect 466380 153762 466408 159200
rect 467196 156528 467248 156534
rect 467196 156470 467248 156476
rect 466288 153734 466408 153762
rect 466184 153672 466236 153678
rect 466184 153614 466236 153620
rect 466000 152380 466052 152386
rect 466000 152322 466052 152328
rect 466012 151994 466040 152322
rect 465000 151966 465060 151994
rect 465704 151966 466040 151994
rect 466196 151858 466224 153614
rect 466288 153066 466316 153734
rect 466276 153060 466328 153066
rect 466276 153002 466328 153008
rect 467208 151994 467236 156470
rect 467300 153950 467328 159200
rect 467748 155848 467800 155854
rect 467748 155790 467800 155796
rect 467288 153944 467340 153950
rect 467288 153886 467340 153892
rect 467760 151994 467788 155790
rect 468312 154698 468340 159200
rect 469324 155582 469352 159200
rect 469864 156596 469916 156602
rect 469864 156538 469916 156544
rect 469312 155576 469364 155582
rect 469312 155518 469364 155524
rect 468300 154692 468352 154698
rect 468300 154634 468352 154640
rect 469128 153740 469180 153746
rect 469128 153682 469180 153688
rect 468576 152448 468628 152454
rect 468576 152390 468628 152396
rect 468588 151994 468616 152390
rect 469140 151994 469168 153682
rect 469876 151994 469904 156538
rect 470244 152998 470272 159200
rect 471256 157146 471284 159200
rect 471244 157140 471296 157146
rect 471244 157082 471296 157088
rect 472176 155718 472204 159200
rect 472440 157344 472492 157350
rect 472440 157286 472492 157292
rect 472164 155712 472216 155718
rect 472164 155654 472216 155660
rect 471796 154556 471848 154562
rect 471796 154498 471848 154504
rect 470324 153808 470376 153814
rect 470324 153750 470376 153756
rect 470232 152992 470284 152998
rect 470232 152934 470284 152940
rect 470336 151994 470364 153750
rect 471152 153196 471204 153202
rect 471152 153138 471204 153144
rect 471164 151994 471192 153138
rect 471808 151994 471836 154498
rect 472452 151994 472480 157286
rect 473084 155780 473136 155786
rect 473084 155722 473136 155728
rect 473096 151994 473124 155722
rect 473188 155281 473216 159200
rect 473728 157276 473780 157282
rect 473728 157218 473780 157224
rect 473174 155272 473230 155281
rect 473174 155207 473230 155216
rect 473740 151994 473768 157218
rect 474200 157078 474228 159200
rect 474464 157140 474516 157146
rect 474464 157082 474516 157088
rect 474188 157072 474240 157078
rect 474188 157014 474240 157020
rect 474476 151994 474504 157082
rect 475120 157010 475148 159200
rect 476028 157072 476080 157078
rect 476028 157014 476080 157020
rect 475108 157004 475160 157010
rect 475108 156946 475160 156952
rect 475752 153128 475804 153134
rect 475752 153070 475804 153076
rect 475108 153060 475160 153066
rect 475108 153002 475160 153008
rect 475120 151994 475148 153002
rect 475764 151994 475792 153070
rect 466992 151966 467236 151994
rect 467636 151966 467788 151994
rect 468280 151966 468616 151994
rect 468924 151966 469168 151994
rect 469568 151966 469904 151994
rect 470212 151966 470364 151994
rect 470856 151966 471192 151994
rect 471500 151966 471836 151994
rect 472144 151966 472480 151994
rect 472788 151966 473124 151994
rect 473432 151966 473768 151994
rect 474168 151966 474504 151994
rect 474812 151966 475148 151994
rect 475456 151966 475792 151994
rect 476040 151994 476068 157014
rect 476132 155514 476160 159200
rect 476948 157004 477000 157010
rect 476948 156946 477000 156952
rect 476120 155508 476172 155514
rect 476120 155450 476172 155456
rect 476960 151994 476988 156946
rect 477052 155650 477080 159200
rect 477314 156768 477370 156777
rect 477314 156703 477370 156712
rect 477040 155644 477092 155650
rect 477040 155586 477092 155592
rect 476040 151966 476100 151994
rect 476744 151966 476988 151994
rect 477328 151994 477356 156703
rect 478064 152930 478092 159200
rect 479076 156942 479104 159200
rect 479064 156936 479116 156942
rect 479064 156878 479116 156884
rect 478328 155712 478380 155718
rect 478328 155654 478380 155660
rect 478052 152924 478104 152930
rect 478052 152866 478104 152872
rect 478340 151994 478368 155654
rect 479616 155644 479668 155650
rect 479616 155586 479668 155592
rect 478788 152992 478840 152998
rect 478788 152934 478840 152940
rect 478800 151994 478828 152934
rect 479628 151994 479656 155586
rect 479996 152862 480024 159200
rect 480076 156936 480128 156942
rect 480076 156878 480128 156884
rect 479984 152856 480036 152862
rect 479984 152798 480036 152804
rect 480088 151994 480116 156878
rect 481008 155446 481036 159200
rect 481928 156874 481956 159200
rect 482940 157214 482968 159200
rect 482928 157208 482980 157214
rect 482928 157150 482980 157156
rect 481916 156868 481968 156874
rect 481916 156810 481968 156816
rect 483952 156806 483980 159200
rect 484216 156868 484268 156874
rect 484216 156810 484268 156816
rect 483940 156800 483992 156806
rect 483940 156742 483992 156748
rect 481546 156632 481602 156641
rect 481546 156567 481602 156576
rect 480996 155440 481048 155446
rect 480996 155382 481048 155388
rect 480904 154488 480956 154494
rect 480904 154430 480956 154436
rect 480916 151994 480944 154430
rect 481560 151994 481588 156567
rect 482192 155576 482244 155582
rect 482192 155518 482244 155524
rect 482204 151994 482232 155518
rect 483572 155440 483624 155446
rect 483572 155382 483624 155388
rect 482836 152924 482888 152930
rect 482836 152866 482888 152872
rect 482848 151994 482876 152866
rect 483584 151994 483612 155382
rect 484228 151994 484256 156810
rect 484768 155508 484820 155514
rect 484768 155450 484820 155456
rect 484780 151994 484808 155450
rect 484872 155378 484900 159200
rect 484952 157208 485004 157214
rect 484952 157150 485004 157156
rect 484860 155372 484912 155378
rect 484860 155314 484912 155320
rect 484964 154494 484992 157150
rect 484952 154488 485004 154494
rect 484952 154430 485004 154436
rect 485504 152856 485556 152862
rect 485504 152798 485556 152804
rect 485516 151994 485544 152798
rect 485884 152130 485912 159200
rect 486700 156800 486752 156806
rect 486700 156742 486752 156748
rect 486148 152788 486200 152794
rect 486148 152730 486200 152736
rect 477328 151966 477388 151994
rect 478032 151966 478368 151994
rect 478676 151966 478828 151994
rect 479320 151966 479656 151994
rect 479964 151966 480116 151994
rect 480608 151966 480944 151994
rect 481252 151966 481588 151994
rect 481896 151966 482232 151994
rect 482540 151966 482876 151994
rect 483276 151966 483612 151994
rect 483920 151966 484256 151994
rect 484564 151966 484808 151994
rect 485208 151966 485544 151994
rect 485700 152102 485912 152130
rect 485700 151978 485728 152102
rect 486160 151994 486188 152730
rect 486712 151994 486740 156742
rect 486804 156058 486832 159200
rect 486792 156052 486844 156058
rect 486792 155994 486844 156000
rect 487068 154488 487120 154494
rect 487068 154430 487120 154436
rect 485688 151972 485740 151978
rect 485852 151966 486188 151994
rect 486496 151966 486740 151994
rect 487080 151994 487108 154430
rect 487816 152726 487844 159200
rect 488356 155372 488408 155378
rect 488356 155314 488408 155320
rect 487804 152720 487856 152726
rect 487804 152662 487856 152668
rect 488080 152720 488132 152726
rect 488080 152662 488132 152668
rect 488092 151994 488120 152662
rect 487080 151966 487140 151994
rect 487784 151966 488120 151994
rect 488368 151994 488396 155314
rect 488828 152658 488856 159200
rect 489748 156738 489776 159200
rect 489736 156732 489788 156738
rect 489736 156674 489788 156680
rect 490656 156732 490708 156738
rect 490656 156674 490708 156680
rect 489642 155952 489698 155961
rect 489642 155887 489698 155896
rect 488816 152652 488868 152658
rect 488816 152594 488868 152600
rect 489368 152652 489420 152658
rect 489368 152594 489420 152600
rect 489380 151994 489408 152594
rect 488368 151966 488428 151994
rect 489072 151966 489408 151994
rect 489656 151994 489684 155887
rect 490668 151994 490696 156674
rect 490760 152046 490788 159200
rect 491680 156670 491708 159200
rect 491668 156664 491720 156670
rect 491668 156606 491720 156612
rect 491944 156664 491996 156670
rect 491944 156606 491996 156612
rect 491208 154420 491260 154426
rect 491208 154362 491260 154368
rect 489656 151966 489716 151994
rect 490360 151966 490696 151994
rect 490748 152040 490800 152046
rect 491220 151994 491248 154362
rect 491956 151994 491984 156606
rect 492692 156262 492720 159200
rect 492680 156256 492732 156262
rect 492680 156198 492732 156204
rect 492586 155680 492642 155689
rect 492586 155615 492642 155624
rect 492600 151994 492628 155615
rect 493324 152584 493376 152590
rect 493324 152526 493376 152532
rect 493336 151994 493364 152526
rect 493704 152522 493732 159200
rect 494624 156126 494652 159200
rect 494612 156120 494664 156126
rect 494612 156062 494664 156068
rect 495254 155544 495310 155553
rect 495254 155479 495310 155488
rect 493968 154352 494020 154358
rect 493968 154294 494020 154300
rect 493692 152516 493744 152522
rect 493692 152458 493744 152464
rect 493980 151994 494008 154294
rect 494612 154284 494664 154290
rect 494612 154226 494664 154232
rect 494624 151994 494652 154226
rect 495268 151994 495296 155479
rect 495636 152114 495664 159200
rect 495898 155816 495954 155825
rect 495898 155751 495954 155760
rect 495624 152108 495676 152114
rect 495624 152050 495676 152056
rect 495912 151994 495940 155751
rect 496556 154306 496584 159200
rect 497186 155408 497242 155417
rect 497186 155343 497242 155352
rect 496464 154278 496584 154306
rect 496464 152114 496492 154278
rect 496544 154216 496596 154222
rect 496544 154158 496596 154164
rect 496452 152108 496504 152114
rect 496452 152050 496504 152056
rect 496556 151994 496584 154158
rect 497200 151994 497228 155343
rect 497568 152182 497596 159200
rect 498580 156330 498608 159200
rect 498568 156324 498620 156330
rect 498568 156266 498620 156272
rect 499500 156194 499528 159200
rect 499488 156188 499540 156194
rect 499488 156130 499540 156136
rect 499394 155272 499450 155281
rect 499394 155207 499450 155216
rect 497832 154148 497884 154154
rect 497832 154090 497884 154096
rect 497556 152176 497608 152182
rect 497556 152118 497608 152124
rect 497844 151994 497872 154090
rect 499120 154080 499172 154086
rect 499120 154022 499172 154028
rect 498108 152516 498160 152522
rect 498108 152458 498160 152464
rect 490748 151982 490800 151988
rect 491004 151966 491248 151994
rect 491648 151966 491984 151994
rect 492292 151966 492628 151994
rect 493028 151966 493364 151994
rect 493672 151966 494008 151994
rect 494316 151966 494652 151994
rect 494960 151966 495296 151994
rect 495604 151966 495940 151994
rect 496248 151966 496584 151994
rect 496892 151966 497228 151994
rect 497536 151966 497872 151994
rect 498120 151994 498148 152458
rect 499132 151994 499160 154022
rect 498120 151966 498180 151994
rect 498824 151966 499160 151994
rect 499408 151994 499436 155207
rect 500132 154624 500184 154630
rect 500132 154566 500184 154572
rect 500144 153882 500172 154566
rect 500132 153876 500184 153882
rect 500132 153818 500184 153824
rect 500408 153536 500460 153542
rect 500408 153478 500460 153484
rect 500420 151994 500448 153478
rect 500512 152250 500540 159200
rect 501432 155242 501460 159200
rect 502444 155310 502472 159200
rect 502432 155304 502484 155310
rect 502432 155246 502484 155252
rect 502984 155304 503036 155310
rect 502984 155246 503036 155252
rect 501420 155236 501472 155242
rect 501420 155178 501472 155184
rect 502248 155236 502300 155242
rect 502248 155178 502300 155184
rect 500868 154012 500920 154018
rect 500868 153954 500920 153960
rect 500500 152244 500552 152250
rect 500500 152186 500552 152192
rect 500880 151994 500908 153954
rect 501696 153876 501748 153882
rect 501696 153818 501748 153824
rect 501708 151994 501736 153818
rect 502260 151994 502288 155178
rect 502996 153542 503024 155246
rect 503364 154630 503392 159200
rect 504376 156398 504404 159200
rect 504364 156392 504416 156398
rect 504364 156334 504416 156340
rect 505388 154766 505416 159200
rect 505376 154760 505428 154766
rect 505376 154702 505428 154708
rect 503352 154624 503404 154630
rect 503352 154566 503404 154572
rect 503076 153944 503128 153950
rect 503076 153886 503128 153892
rect 502984 153536 503036 153542
rect 502984 153478 503036 153484
rect 503088 151994 503116 153886
rect 506308 153474 506336 159200
rect 506940 155984 506992 155990
rect 506940 155926 506992 155932
rect 506296 153468 506348 153474
rect 506296 153410 506348 153416
rect 505650 153232 505706 153241
rect 505650 153167 505706 153176
rect 499408 151966 499468 151994
rect 500112 151966 500448 151994
rect 500756 151966 500908 151994
rect 501400 151966 501736 151994
rect 502136 151966 502288 151994
rect 502780 151966 503116 151994
rect 505664 151994 505692 153167
rect 506952 151994 506980 155926
rect 507320 152318 507348 159200
rect 508240 154902 508268 159200
rect 509252 154970 509280 159200
rect 510160 157412 510212 157418
rect 510160 157354 510212 157360
rect 509240 154964 509292 154970
rect 509240 154906 509292 154912
rect 508228 154896 508280 154902
rect 508228 154838 508280 154844
rect 509514 153368 509570 153377
rect 509514 153303 509570 153312
rect 507308 152312 507360 152318
rect 507308 152254 507360 152260
rect 505664 151966 506000 151994
rect 506644 151966 506980 151994
rect 509528 151994 509556 153303
rect 510172 151994 510200 157354
rect 510264 154834 510292 159200
rect 510252 154828 510304 154834
rect 510252 154770 510304 154776
rect 511184 154698 511212 159200
rect 512196 155038 512224 159200
rect 513116 156466 513144 159200
rect 513104 156460 513156 156466
rect 513104 156402 513156 156408
rect 514128 155106 514156 159200
rect 514116 155100 514168 155106
rect 514116 155042 514168 155048
rect 512184 155032 512236 155038
rect 512184 154974 512236 154980
rect 511172 154692 511224 154698
rect 511172 154634 511224 154640
rect 513470 153640 513526 153649
rect 515140 153610 515168 159200
rect 516060 155174 516088 159200
rect 517072 155922 517100 159200
rect 517060 155916 517112 155922
rect 517060 155858 517112 155864
rect 516048 155168 516100 155174
rect 516048 155110 516100 155116
rect 517518 154048 517574 154057
rect 517518 153983 517574 153992
rect 516690 153912 516746 153921
rect 516690 153847 516746 153856
rect 516138 153776 516194 153785
rect 516138 153711 516194 153720
rect 513470 153575 513526 153584
rect 515128 153604 515180 153610
rect 510894 153504 510950 153513
rect 510894 153439 510950 153448
rect 511816 153468 511868 153474
rect 510908 151994 510936 153439
rect 511816 153410 511868 153416
rect 511828 151994 511856 153410
rect 512736 153400 512788 153406
rect 512736 153342 512788 153348
rect 512748 151994 512776 153342
rect 512828 153332 512880 153338
rect 512828 153274 512880 153280
rect 509528 151966 509864 151994
rect 510172 151966 510508 151994
rect 510908 151966 511244 151994
rect 511828 151966 511888 151994
rect 512532 151966 512776 151994
rect 512840 151994 512868 153274
rect 513484 151994 513512 153575
rect 515128 153546 515180 153552
rect 514116 153264 514168 153270
rect 514116 153206 514168 153212
rect 515404 153264 515456 153270
rect 515404 153206 515456 153212
rect 514128 151994 514156 153206
rect 515416 151994 515444 153206
rect 512840 151966 513176 151994
rect 513484 151966 513820 151994
rect 514128 151966 514464 151994
rect 515108 151966 515444 151994
rect 516152 151994 516180 153711
rect 516704 151994 516732 153847
rect 517532 151994 517560 153983
rect 517992 152386 518020 159200
rect 519004 153678 519032 159200
rect 520016 156534 520044 159200
rect 520004 156528 520056 156534
rect 520004 156470 520056 156476
rect 520936 155854 520964 159200
rect 520924 155848 520976 155854
rect 520924 155790 520976 155796
rect 519266 154184 519322 154193
rect 519266 154119 519322 154128
rect 518992 153672 519044 153678
rect 518992 153614 519044 153620
rect 517980 152380 518032 152386
rect 517980 152322 518032 152328
rect 519280 151994 519308 154119
rect 520280 153332 520332 153338
rect 520280 153274 520332 153280
rect 516152 151966 516396 151994
rect 516704 151966 517040 151994
rect 517532 151966 517684 151994
rect 519280 151966 519616 151994
rect 485688 151914 485740 151920
rect 508226 151872 508282 151881
rect 244424 151852 244536 151858
rect 244372 151846 244536 151852
rect 212448 151836 212500 151842
rect 244384 151830 244536 151846
rect 247112 151830 247264 151858
rect 252020 151842 252356 151858
rect 252008 151836 252356 151842
rect 212448 151778 212500 151784
rect 252060 151830 252356 151836
rect 364168 151830 364228 151858
rect 376496 151830 376556 151858
rect 386248 151830 386308 151858
rect 398576 151830 398636 151858
rect 408328 151830 408388 151858
rect 420748 151830 420808 151858
rect 431788 151830 431848 151858
rect 433076 151830 433136 151858
rect 442828 151830 442888 151858
rect 455248 151830 455308 151858
rect 466196 151830 466348 151858
rect 503424 151842 503668 151858
rect 503424 151836 503680 151842
rect 503424 151830 503628 151836
rect 252008 151778 252060 151784
rect 508282 151830 508576 151858
rect 508226 151807 508282 151816
rect 503628 151778 503680 151784
rect 212908 151768 212960 151774
rect 212960 151716 213256 151722
rect 212908 151710 213256 151716
rect 212920 151694 213256 151710
rect 504712 151706 505048 151722
rect 504712 151700 505060 151706
rect 504712 151694 505008 151700
rect 505008 151642 505060 151648
rect 197268 151632 197320 151638
rect 506940 151632 506992 151638
rect 197268 151574 197320 151580
rect 503732 151570 504068 151586
rect 503720 151564 504068 151570
rect 503772 151558 504068 151564
rect 505356 151570 505692 151586
rect 506992 151580 507288 151586
rect 506940 151574 507288 151580
rect 505356 151564 505704 151570
rect 505356 151558 505652 151564
rect 503720 151506 503772 151512
rect 506952 151558 507288 151574
rect 505652 151506 505704 151512
rect 507768 151360 507820 151366
rect 508872 151360 508924 151366
rect 507820 151308 507932 151314
rect 507768 151302 507932 151308
rect 515404 151360 515456 151366
rect 508924 151308 509220 151314
rect 508872 151302 509220 151308
rect 518624 151360 518676 151366
rect 515456 151308 515752 151314
rect 515404 151302 515752 151308
rect 507780 151286 507932 151302
rect 508884 151286 509220 151302
rect 515416 151286 515752 151302
rect 518328 151308 518624 151314
rect 519268 151360 519320 151366
rect 518328 151302 518676 151308
rect 518972 151308 519268 151314
rect 518972 151302 519320 151308
rect 518328 151286 518664 151302
rect 518972 151286 519308 151302
rect 119896 67448 119948 67454
rect 119896 67390 119948 67396
rect 119896 20868 119948 20874
rect 119896 20810 119948 20816
rect 119908 5166 119936 20810
rect 119896 5160 119948 5166
rect 119896 5102 119948 5108
rect 119816 4678 120028 4706
rect 444392 4690 444544 4706
rect 119724 3998 119936 4026
rect 119712 3392 119764 3398
rect 119712 3334 119764 3340
rect 119618 2680 119674 2689
rect 119618 2615 119674 2624
rect 119528 2168 119580 2174
rect 119528 2110 119580 2116
rect 118330 1864 118386 1873
rect 118330 1799 118386 1808
rect 119724 1714 119752 3334
rect 119632 1686 119752 1714
rect 116860 1216 116912 1222
rect 116860 1158 116912 1164
rect 119632 800 119660 1686
rect 119908 1154 119936 3998
rect 120000 2553 120028 4678
rect 444380 4684 444544 4690
rect 444432 4678 444544 4684
rect 463036 4690 463372 4706
rect 463036 4684 463384 4690
rect 463036 4678 463332 4684
rect 444380 4626 444432 4632
rect 463332 4626 463384 4632
rect 121472 4134 121532 4162
rect 124232 4134 124568 4162
rect 127268 4134 127604 4162
rect 130396 4134 130732 4162
rect 133432 4134 133768 4162
rect 136652 4134 136896 4162
rect 139596 4134 139932 4162
rect 142724 4134 143060 4162
rect 145760 4134 146096 4162
rect 149072 4134 149224 4162
rect 152016 4134 152260 4162
rect 154960 4134 155296 4162
rect 158088 4134 158424 4162
rect 161124 4134 161460 4162
rect 164252 4134 164588 4162
rect 167288 4134 167624 4162
rect 170416 4134 170752 4162
rect 173452 4134 173788 4162
rect 176672 4134 176916 4162
rect 179616 4134 179952 4162
rect 182652 4134 182988 4162
rect 185780 4134 186116 4162
rect 189092 4134 189152 4162
rect 191944 4134 192280 4162
rect 194980 4134 195316 4162
rect 198108 4134 198444 4162
rect 201144 4134 201480 4162
rect 204272 4134 204608 4162
rect 207308 4134 207644 4162
rect 210344 4134 210680 4162
rect 213472 4134 213808 4162
rect 121472 2990 121500 4134
rect 124232 3058 124260 4134
rect 127268 3126 127296 4134
rect 130396 3194 130424 4134
rect 133432 3262 133460 4134
rect 136652 3330 136680 4134
rect 136640 3324 136692 3330
rect 136640 3266 136692 3272
rect 133420 3256 133472 3262
rect 133420 3198 133472 3204
rect 135536 3256 135588 3262
rect 135536 3198 135588 3204
rect 130384 3188 130436 3194
rect 130384 3130 130436 3136
rect 127256 3120 127308 3126
rect 127256 3062 127308 3068
rect 130292 3120 130344 3126
rect 130292 3062 130344 3068
rect 124220 3052 124272 3058
rect 124220 2994 124272 3000
rect 121460 2984 121512 2990
rect 121460 2926 121512 2932
rect 124956 2984 125008 2990
rect 124956 2926 125008 2932
rect 119986 2544 120042 2553
rect 119986 2479 120042 2488
rect 119896 1148 119948 1154
rect 119896 1090 119948 1096
rect 124968 800 124996 2926
rect 130304 800 130332 3062
rect 135548 800 135576 3198
rect 139596 1766 139624 4134
rect 140872 3324 140924 3330
rect 140872 3266 140924 3272
rect 139584 1760 139636 1766
rect 139584 1702 139636 1708
rect 140884 800 140912 3266
rect 142724 1698 142752 4134
rect 142712 1692 142764 1698
rect 142712 1634 142764 1640
rect 145760 1630 145788 4134
rect 146116 3596 146168 3602
rect 146116 3538 146168 3544
rect 146128 1698 146156 3538
rect 146208 3392 146260 3398
rect 146208 3334 146260 3340
rect 146116 1692 146168 1698
rect 146116 1634 146168 1640
rect 145748 1624 145800 1630
rect 145748 1566 145800 1572
rect 146220 800 146248 3334
rect 149072 1562 149100 4134
rect 149152 3664 149204 3670
rect 149152 3606 149204 3612
rect 149164 1766 149192 3606
rect 151544 3528 151596 3534
rect 151544 3470 151596 3476
rect 149152 1760 149204 1766
rect 149152 1702 149204 1708
rect 149060 1556 149112 1562
rect 149060 1498 149112 1504
rect 151556 800 151584 3470
rect 152016 2786 152044 4134
rect 153108 3732 153160 3738
rect 153108 3674 153160 3680
rect 153120 2786 153148 3674
rect 152004 2780 152056 2786
rect 152004 2722 152056 2728
rect 153108 2780 153160 2786
rect 153108 2722 153160 2728
rect 154960 1698 154988 4134
rect 156512 3868 156564 3874
rect 156512 3810 156564 3816
rect 156524 2718 156552 3810
rect 156880 2984 156932 2990
rect 156880 2926 156932 2932
rect 156512 2712 156564 2718
rect 156512 2654 156564 2660
rect 154948 1692 155000 1698
rect 154948 1634 155000 1640
rect 156892 800 156920 2926
rect 158088 1766 158116 4134
rect 161124 2786 161152 4134
rect 162768 3800 162820 3806
rect 162768 3742 162820 3748
rect 162216 3596 162268 3602
rect 162216 3538 162268 3544
rect 161112 2780 161164 2786
rect 161112 2722 161164 2728
rect 158076 1760 158128 1766
rect 158076 1702 158128 1708
rect 162228 800 162256 3538
rect 162780 2718 162808 3742
rect 164252 2786 164280 4134
rect 165528 3936 165580 3942
rect 165528 3878 165580 3884
rect 165540 2786 165568 3878
rect 164240 2780 164292 2786
rect 164240 2722 164292 2728
rect 165528 2780 165580 2786
rect 165528 2722 165580 2728
rect 167288 2718 167316 4134
rect 167368 4004 167420 4010
rect 167368 3946 167420 3952
rect 167380 2718 167408 3946
rect 167460 3664 167512 3670
rect 167460 3606 167512 3612
rect 162768 2712 162820 2718
rect 162768 2654 162820 2660
rect 167276 2712 167328 2718
rect 167276 2654 167328 2660
rect 167368 2712 167420 2718
rect 167368 2654 167420 2660
rect 167472 800 167500 3606
rect 170416 2786 170444 4134
rect 172796 3936 172848 3942
rect 172796 3878 172848 3884
rect 170404 2780 170456 2786
rect 170404 2722 170456 2728
rect 172808 800 172836 3878
rect 173452 3466 173480 4134
rect 173440 3460 173492 3466
rect 173440 3402 173492 3408
rect 176672 2718 176700 4134
rect 176752 4072 176804 4078
rect 176752 4014 176804 4020
rect 176764 2786 176792 4014
rect 178132 3732 178184 3738
rect 178132 3674 178184 3680
rect 176752 2780 176804 2786
rect 176752 2722 176804 2728
rect 176660 2712 176712 2718
rect 176660 2654 176712 2660
rect 178144 800 178172 3674
rect 179616 2854 179644 4134
rect 179604 2848 179656 2854
rect 179604 2790 179656 2796
rect 182652 2786 182680 4134
rect 183468 3800 183520 3806
rect 183468 3742 183520 3748
rect 182640 2780 182692 2786
rect 182640 2722 182692 2728
rect 183480 800 183508 3742
rect 185780 3058 185808 4134
rect 188804 3868 188856 3874
rect 188804 3810 188856 3816
rect 185768 3052 185820 3058
rect 185768 2994 185820 3000
rect 188816 800 188844 3810
rect 189092 3126 189120 4134
rect 191944 3194 191972 4134
rect 194980 3262 195008 4134
rect 198108 3330 198136 4134
rect 201144 3398 201172 4134
rect 204272 3534 204300 4134
rect 204260 3528 204312 3534
rect 204260 3470 204312 3476
rect 201132 3392 201184 3398
rect 201132 3334 201184 3340
rect 204720 3392 204772 3398
rect 204720 3334 204772 3340
rect 198096 3324 198148 3330
rect 198096 3266 198148 3272
rect 199384 3324 199436 3330
rect 199384 3266 199436 3272
rect 194968 3256 195020 3262
rect 194968 3198 195020 3204
rect 191932 3188 191984 3194
rect 191932 3130 191984 3136
rect 189080 3120 189132 3126
rect 189080 3062 189132 3068
rect 194140 2848 194192 2854
rect 194140 2790 194192 2796
rect 194152 800 194180 2790
rect 199396 800 199424 3266
rect 204732 800 204760 3334
rect 207308 2990 207336 4134
rect 210344 3602 210372 4134
rect 213472 3670 213500 4134
rect 216830 3942 216858 4148
rect 219636 4134 219972 4162
rect 222672 4134 223008 4162
rect 225800 4134 226136 4162
rect 229112 4134 229172 4162
rect 231964 4134 232300 4162
rect 235000 4134 235336 4162
rect 238036 4134 238372 4162
rect 241164 4134 241500 4162
rect 244292 4134 244536 4162
rect 247328 4134 247664 4162
rect 250364 4134 250700 4162
rect 253492 4134 253828 4162
rect 256620 4134 256864 4162
rect 259656 4134 259992 4162
rect 262692 4134 263028 4162
rect 265728 4134 266064 4162
rect 269132 4134 269192 4162
rect 216818 3936 216870 3942
rect 216818 3878 216870 3884
rect 219636 3738 219664 4134
rect 222672 3806 222700 4134
rect 225800 3874 225828 4134
rect 225788 3868 225840 3874
rect 225788 3810 225840 3816
rect 222660 3800 222712 3806
rect 222660 3742 222712 3748
rect 219624 3732 219676 3738
rect 219624 3674 219676 3680
rect 213460 3664 213512 3670
rect 213460 3606 213512 3612
rect 210332 3596 210384 3602
rect 210332 3538 210384 3544
rect 226064 3256 226116 3262
rect 226064 3198 226116 3204
rect 215392 3188 215444 3194
rect 215392 3130 215444 3136
rect 210056 3120 210108 3126
rect 210056 3062 210108 3068
rect 207296 2984 207348 2990
rect 207296 2926 207348 2932
rect 210068 800 210096 3062
rect 215404 800 215432 3130
rect 220728 2984 220780 2990
rect 220728 2926 220780 2932
rect 220740 800 220768 2926
rect 226076 800 226104 3198
rect 229112 2854 229140 4134
rect 231964 3330 231992 4134
rect 235000 3398 235028 4134
rect 234988 3392 235040 3398
rect 234988 3334 235040 3340
rect 231952 3324 232004 3330
rect 231952 3266 232004 3272
rect 238036 3126 238064 4134
rect 241164 3194 241192 4134
rect 241152 3188 241204 3194
rect 241152 3130 241204 3136
rect 238024 3120 238076 3126
rect 238024 3062 238076 3068
rect 241980 3120 242032 3126
rect 241980 3062 242032 3068
rect 231308 3052 231360 3058
rect 231308 2994 231360 3000
rect 229100 2848 229152 2854
rect 229100 2790 229152 2796
rect 231320 800 231348 2994
rect 236644 2848 236696 2854
rect 236644 2790 236696 2796
rect 236656 800 236684 2790
rect 241992 800 242020 3062
rect 244292 2990 244320 4134
rect 247328 3262 247356 4134
rect 247408 3392 247460 3398
rect 247408 3334 247460 3340
rect 247316 3256 247368 3262
rect 247316 3198 247368 3204
rect 244280 2984 244332 2990
rect 244280 2926 244332 2932
rect 247420 1714 247448 3334
rect 250364 3058 250392 4134
rect 250352 3052 250404 3058
rect 250352 2994 250404 3000
rect 252652 2984 252704 2990
rect 252652 2926 252704 2932
rect 247328 1686 247448 1714
rect 247328 800 247356 1686
rect 252664 800 252692 2926
rect 253492 2786 253520 4134
rect 256620 3126 256648 4134
rect 259656 3398 259684 4134
rect 259644 3392 259696 3398
rect 259644 3334 259696 3340
rect 256608 3120 256660 3126
rect 256608 3062 256660 3068
rect 257988 3052 258040 3058
rect 257988 2994 258040 3000
rect 253480 2780 253532 2786
rect 253480 2722 253532 2728
rect 258000 800 258028 2994
rect 262692 2990 262720 4134
rect 265728 3058 265756 4134
rect 268568 3936 268620 3942
rect 268568 3878 268620 3884
rect 265716 3052 265768 3058
rect 265716 2994 265768 3000
rect 262680 2984 262732 2990
rect 262680 2926 262732 2932
rect 263232 2848 263284 2854
rect 263232 2790 263284 2796
rect 263244 800 263272 2790
rect 268580 800 268608 3878
rect 269132 2786 269160 4134
rect 272214 3942 272242 4148
rect 275342 3942 275370 4148
rect 278392 4134 278728 4162
rect 272202 3936 272254 3942
rect 272202 3878 272254 3884
rect 273904 3936 273956 3942
rect 273904 3878 273956 3884
rect 275330 3936 275382 3942
rect 275330 3878 275382 3884
rect 269120 2780 269172 2786
rect 269120 2722 269172 2728
rect 273916 800 273944 3878
rect 278700 1766 278728 4134
rect 281506 3942 281534 4148
rect 284556 4134 284892 4162
rect 287684 4134 288020 4162
rect 290720 4134 291056 4162
rect 293756 4134 293908 4162
rect 296884 4134 297220 4162
rect 299920 4134 300256 4162
rect 303048 4134 303384 4162
rect 306084 4134 306236 4162
rect 309212 4134 309548 4162
rect 312248 4134 312584 4162
rect 315376 4134 315712 4162
rect 318412 4134 318748 4162
rect 281494 3936 281546 3942
rect 281494 3878 281546 3884
rect 284576 3936 284628 3942
rect 284576 3878 284628 3884
rect 278688 1760 278740 1766
rect 278688 1702 278740 1708
rect 279240 1760 279292 1766
rect 279240 1702 279292 1708
rect 279252 800 279280 1702
rect 284588 800 284616 3878
rect 284864 2786 284892 4134
rect 287992 2786 288020 4134
rect 289636 2848 289688 2854
rect 289688 2796 289952 2802
rect 289636 2790 289952 2796
rect 284852 2780 284904 2786
rect 284852 2722 284904 2728
rect 287980 2780 288032 2786
rect 289648 2774 289952 2790
rect 287980 2722 288032 2728
rect 289924 800 289952 2774
rect 291028 1766 291056 4134
rect 291016 1760 291068 1766
rect 291016 1702 291068 1708
rect 293880 1630 293908 4134
rect 295156 2848 295208 2854
rect 295156 2790 295208 2796
rect 293868 1624 293920 1630
rect 293868 1566 293920 1572
rect 295168 800 295196 2790
rect 297192 1562 297220 4134
rect 300228 1698 300256 4134
rect 303356 2854 303384 4134
rect 306208 3262 306236 4134
rect 309520 3398 309548 4134
rect 309508 3392 309560 3398
rect 309508 3334 309560 3340
rect 306196 3256 306248 3262
rect 306196 3198 306248 3204
rect 312556 3058 312584 4134
rect 312544 3052 312596 3058
rect 312544 2994 312596 3000
rect 315684 2990 315712 4134
rect 318720 3602 318748 4134
rect 321480 4134 321540 4162
rect 324576 4134 324912 4162
rect 327612 4134 327948 4162
rect 330740 4134 331076 4162
rect 333776 4134 333928 4162
rect 336904 4134 337240 4162
rect 339940 4134 340276 4162
rect 343068 4134 343404 4162
rect 346104 4134 346348 4162
rect 349232 4134 349568 4162
rect 352268 4134 352604 4162
rect 355304 4134 355640 4162
rect 358432 4134 358768 4162
rect 318708 3596 318760 3602
rect 318708 3538 318760 3544
rect 321480 3126 321508 4134
rect 324884 3670 324912 4134
rect 324872 3664 324924 3670
rect 324872 3606 324924 3612
rect 327080 3256 327132 3262
rect 327080 3198 327132 3204
rect 321468 3120 321520 3126
rect 321468 3062 321520 3068
rect 315672 2984 315724 2990
rect 315672 2926 315724 2932
rect 303344 2848 303396 2854
rect 303344 2790 303396 2796
rect 321836 2848 321888 2854
rect 321836 2790 321888 2796
rect 300492 1760 300544 1766
rect 300492 1702 300544 1708
rect 316500 1760 316552 1766
rect 316500 1702 316552 1708
rect 300216 1692 300268 1698
rect 300216 1634 300268 1640
rect 297180 1556 297232 1562
rect 297180 1498 297232 1504
rect 300504 800 300532 1702
rect 311164 1692 311216 1698
rect 311164 1634 311216 1640
rect 305828 1624 305880 1630
rect 305828 1566 305880 1572
rect 305840 800 305868 1566
rect 311176 800 311204 1634
rect 316512 800 316540 1702
rect 321848 800 321876 2790
rect 327092 800 327120 3198
rect 327920 2854 327948 4134
rect 331048 3262 331076 4134
rect 332416 3392 332468 3398
rect 332416 3334 332468 3340
rect 331036 3256 331088 3262
rect 331036 3198 331088 3204
rect 327908 2848 327960 2854
rect 327908 2790 327960 2796
rect 332428 800 332456 3334
rect 333900 3194 333928 4134
rect 337212 3466 337240 4134
rect 337200 3460 337252 3466
rect 337200 3402 337252 3408
rect 333888 3188 333940 3194
rect 333888 3130 333940 3136
rect 340248 3058 340276 4134
rect 343376 3534 343404 4134
rect 343364 3528 343416 3534
rect 343364 3470 343416 3476
rect 337752 3052 337804 3058
rect 337752 2994 337804 3000
rect 340236 3052 340288 3058
rect 340236 2994 340288 3000
rect 337764 800 337792 2994
rect 346320 2990 346348 4134
rect 348424 3596 348476 3602
rect 348424 3538 348476 3544
rect 343088 2984 343140 2990
rect 343088 2926 343140 2932
rect 346308 2984 346360 2990
rect 346308 2926 346360 2932
rect 343100 800 343128 2926
rect 348436 800 348464 3538
rect 349540 1766 349568 4134
rect 352576 3398 352604 4134
rect 352564 3392 352616 3398
rect 352564 3334 352616 3340
rect 353760 3120 353812 3126
rect 353760 3062 353812 3068
rect 349528 1760 349580 1766
rect 349528 1702 349580 1708
rect 353772 800 353800 3062
rect 355612 1698 355640 4134
rect 358740 3330 358768 4134
rect 361408 4134 361468 4162
rect 364596 4134 364932 4162
rect 367632 4134 367968 4162
rect 370760 4134 371096 4162
rect 373796 4134 373948 4162
rect 376924 4134 377260 4162
rect 361408 3874 361436 4134
rect 361396 3868 361448 3874
rect 361396 3810 361448 3816
rect 359004 3664 359056 3670
rect 359004 3606 359056 3612
rect 358728 3324 358780 3330
rect 358728 3266 358780 3272
rect 355600 1692 355652 1698
rect 355600 1634 355652 1640
rect 359016 800 359044 3606
rect 364904 3126 364932 4134
rect 367940 4010 367968 4134
rect 367928 4004 367980 4010
rect 367928 3946 367980 3952
rect 371068 3806 371096 4134
rect 371056 3800 371108 3806
rect 371056 3742 371108 3748
rect 373920 3738 373948 4134
rect 373908 3732 373960 3738
rect 373908 3674 373960 3680
rect 369676 3256 369728 3262
rect 369676 3198 369728 3204
rect 364892 3120 364944 3126
rect 364892 3062 364944 3068
rect 364340 2848 364392 2854
rect 364340 2790 364392 2796
rect 364352 800 364380 2790
rect 369688 800 369716 3198
rect 375012 3188 375064 3194
rect 375012 3130 375064 3136
rect 375024 800 375052 3130
rect 377232 2854 377260 4134
rect 379946 3942 379974 4148
rect 382996 4134 383332 4162
rect 386124 4134 386368 4162
rect 383304 4078 383332 4134
rect 383292 4072 383344 4078
rect 383292 4014 383344 4020
rect 379934 3936 379986 3942
rect 379934 3878 379986 3884
rect 386340 3670 386368 4134
rect 389100 4134 389160 4162
rect 392288 4134 392624 4162
rect 395324 4134 395660 4162
rect 398452 4134 398788 4162
rect 386328 3664 386380 3670
rect 386328 3606 386380 3612
rect 389100 3602 389128 4134
rect 389088 3596 389140 3602
rect 389088 3538 389140 3544
rect 392596 3534 392624 4134
rect 390928 3528 390980 3534
rect 390928 3470 390980 3476
rect 392584 3528 392636 3534
rect 392584 3470 392636 3476
rect 380348 3460 380400 3466
rect 380348 3402 380400 3408
rect 377220 2848 377272 2854
rect 377220 2790 377272 2796
rect 380360 800 380388 3402
rect 385684 3052 385736 3058
rect 385684 2994 385736 3000
rect 385696 800 385724 2994
rect 390940 800 390968 3470
rect 395632 3466 395660 4134
rect 395620 3460 395672 3466
rect 395620 3402 395672 3408
rect 398760 3262 398788 4134
rect 401428 4134 401488 4162
rect 404616 4134 404952 4162
rect 407652 4134 407988 4162
rect 410688 4134 411024 4162
rect 413816 4134 413968 4162
rect 416852 4134 417188 4162
rect 419980 4134 420316 4162
rect 423016 4134 423352 4162
rect 426144 4134 426388 4162
rect 398748 3256 398800 3262
rect 398748 3198 398800 3204
rect 401428 3058 401456 4134
rect 404924 3398 404952 4134
rect 404912 3392 404964 3398
rect 404912 3334 404964 3340
rect 407764 3392 407816 3398
rect 407764 3334 407816 3340
rect 407776 3262 407804 3334
rect 407764 3256 407816 3262
rect 407764 3198 407816 3204
rect 406936 3188 406988 3194
rect 406936 3130 406988 3136
rect 401416 3052 401468 3058
rect 401416 2994 401468 3000
rect 396264 2984 396316 2990
rect 396264 2926 396316 2932
rect 396276 800 396304 2926
rect 401600 1760 401652 1766
rect 401600 1702 401652 1708
rect 401612 800 401640 1702
rect 406948 800 406976 3130
rect 407960 3058 407988 4134
rect 407948 3052 408000 3058
rect 407948 2994 408000 3000
rect 410996 1766 411024 4134
rect 410984 1760 411036 1766
rect 410984 1702 411036 1708
rect 412272 1692 412324 1698
rect 412272 1634 412324 1640
rect 412284 800 412312 1634
rect 413940 1630 413968 4134
rect 417160 2786 417188 4134
rect 417332 3324 417384 3330
rect 417332 3266 417384 3272
rect 417148 2780 417200 2786
rect 417148 2722 417200 2728
rect 413928 1624 413980 1630
rect 413928 1566 413980 1572
rect 2594 0 2650 800
rect 7838 0 7894 800
rect 13174 0 13230 800
rect 18510 0 18566 800
rect 23846 0 23902 800
rect 29182 0 29238 800
rect 34518 0 34574 800
rect 39762 0 39818 800
rect 45098 0 45154 800
rect 50434 0 50490 800
rect 55770 0 55826 800
rect 61106 0 61162 800
rect 66442 0 66498 800
rect 71686 0 71742 800
rect 77022 0 77078 800
rect 82358 0 82414 800
rect 87694 0 87750 800
rect 93030 0 93086 800
rect 98366 0 98422 800
rect 103610 0 103666 800
rect 108946 0 109002 800
rect 114282 0 114338 800
rect 119618 0 119674 800
rect 124954 0 125010 800
rect 130290 0 130346 800
rect 135534 0 135590 800
rect 140870 0 140926 800
rect 146206 0 146262 800
rect 151542 0 151598 800
rect 156878 0 156934 800
rect 162214 0 162270 800
rect 167458 0 167514 800
rect 172794 0 172850 800
rect 178130 0 178186 800
rect 183466 0 183522 800
rect 188802 0 188858 800
rect 194138 0 194194 800
rect 199382 0 199438 800
rect 204718 0 204774 800
rect 210054 0 210110 800
rect 215390 0 215446 800
rect 220726 0 220782 800
rect 226062 0 226118 800
rect 231306 0 231362 800
rect 236642 0 236698 800
rect 241978 0 242034 800
rect 247314 0 247370 800
rect 252650 0 252706 800
rect 257986 0 258042 800
rect 263230 0 263286 800
rect 268566 0 268622 800
rect 273902 0 273958 800
rect 279238 0 279294 800
rect 284574 0 284630 800
rect 289910 0 289966 800
rect 295154 0 295210 800
rect 300490 0 300546 800
rect 305826 0 305882 800
rect 311162 0 311218 800
rect 316498 0 316554 800
rect 321834 0 321890 800
rect 327078 0 327134 800
rect 332414 0 332470 800
rect 337750 0 337806 800
rect 343086 0 343142 800
rect 348422 0 348478 800
rect 353758 0 353814 800
rect 359002 0 359058 800
rect 364338 0 364394 800
rect 369674 0 369730 800
rect 375010 0 375066 800
rect 380346 0 380402 800
rect 385682 0 385738 800
rect 390926 0 390982 800
rect 396262 0 396318 800
rect 401598 0 401654 800
rect 406934 0 406990 800
rect 412270 0 412326 800
rect 417344 762 417372 3266
rect 420288 2718 420316 4134
rect 422852 3868 422904 3874
rect 422852 3810 422904 3816
rect 420276 2712 420328 2718
rect 420276 2654 420328 2660
rect 417528 870 417648 898
rect 417528 762 417556 870
rect 417620 800 417648 870
rect 422864 800 422892 3810
rect 423324 3058 423352 4134
rect 423312 3052 423364 3058
rect 423312 2994 423364 3000
rect 426360 2990 426388 4134
rect 429120 4134 429180 4162
rect 432156 4134 432308 4162
rect 435344 4134 435680 4162
rect 438380 4134 438716 4162
rect 427820 3868 427872 3874
rect 427820 3810 427872 3816
rect 426348 2984 426400 2990
rect 426348 2926 426400 2932
rect 427832 2718 427860 3810
rect 428188 3120 428240 3126
rect 428188 3062 428240 3068
rect 427820 2712 427872 2718
rect 427820 2654 427872 2660
rect 428200 800 428228 3062
rect 429120 1698 429148 4134
rect 432156 2038 432184 4134
rect 433524 4004 433576 4010
rect 433524 3946 433576 3952
rect 432144 2032 432196 2038
rect 432144 1974 432196 1980
rect 429108 1692 429160 1698
rect 429108 1634 429160 1640
rect 433536 800 433564 3946
rect 435652 2718 435680 4134
rect 438688 3126 438716 4134
rect 441172 4134 441508 4162
rect 447336 4134 447672 4162
rect 450372 4134 450708 4162
rect 453500 4134 453836 4162
rect 456812 4134 456872 4162
rect 459664 4134 460000 4162
rect 465736 4134 466072 4162
rect 468864 4134 469200 4162
rect 471992 4134 472236 4162
rect 475028 4134 475364 4162
rect 478064 4134 478400 4162
rect 481192 4134 481528 4162
rect 484412 4134 484564 4162
rect 487356 4134 487692 4162
rect 490392 4134 490728 4162
rect 493428 4134 493764 4162
rect 496832 4134 496892 4162
rect 499684 4134 499928 4162
rect 502720 4134 503056 4162
rect 505756 4134 506092 4162
rect 508884 4134 509220 4162
rect 512012 4134 512256 4162
rect 515048 4134 515384 4162
rect 518084 4134 518420 4162
rect 438860 3800 438912 3806
rect 438860 3742 438912 3748
rect 438676 3120 438728 3126
rect 438676 3062 438728 3068
rect 435640 2712 435692 2718
rect 435640 2654 435692 2660
rect 438872 800 438900 3742
rect 441172 1154 441200 4134
rect 444196 3800 444248 3806
rect 444196 3742 444248 3748
rect 443736 3732 443788 3738
rect 443736 3674 443788 3680
rect 443748 2718 443776 3674
rect 443736 2712 443788 2718
rect 443736 2654 443788 2660
rect 441160 1148 441212 1154
rect 441160 1090 441212 1096
rect 444208 800 444236 3742
rect 447336 1873 447364 4134
rect 449532 2848 449584 2854
rect 449532 2790 449584 2796
rect 447322 1864 447378 1873
rect 447322 1799 447378 1808
rect 449544 800 449572 2790
rect 450372 2009 450400 4134
rect 450358 2000 450414 2009
rect 450358 1935 450414 1944
rect 453500 1222 453528 4134
rect 454776 3936 454828 3942
rect 454776 3878 454828 3884
rect 454684 3800 454736 3806
rect 454684 3742 454736 3748
rect 454696 2786 454724 3742
rect 454684 2780 454736 2786
rect 454684 2722 454736 2728
rect 453488 1216 453540 1222
rect 453488 1158 453540 1164
rect 454788 800 454816 3878
rect 456812 2145 456840 4134
rect 456798 2136 456854 2145
rect 456798 2071 456854 2080
rect 459664 1290 459692 4134
rect 460112 4072 460164 4078
rect 460112 4014 460164 4020
rect 459652 1284 459704 1290
rect 459652 1226 459704 1232
rect 460124 800 460152 4014
rect 465448 3664 465500 3670
rect 465448 3606 465500 3612
rect 465460 800 465488 3606
rect 465736 2281 465764 4134
rect 465722 2272 465778 2281
rect 465722 2207 465778 2216
rect 468864 1426 468892 4134
rect 470784 3596 470836 3602
rect 470784 3538 470836 3544
rect 468852 1420 468904 1426
rect 468852 1362 468904 1368
rect 470796 800 470824 3538
rect 471992 2417 472020 4134
rect 475028 3097 475056 4134
rect 476120 3528 476172 3534
rect 476120 3470 476172 3476
rect 475014 3088 475070 3097
rect 475014 3023 475070 3032
rect 471978 2408 472034 2417
rect 471978 2343 472034 2352
rect 476132 800 476160 3470
rect 478064 1358 478092 4134
rect 481192 2553 481220 4134
rect 481456 3460 481508 3466
rect 481456 3402 481508 3408
rect 481178 2544 481234 2553
rect 481178 2479 481234 2488
rect 478052 1352 478104 1358
rect 478052 1294 478104 1300
rect 481468 800 481496 3402
rect 484308 2848 484360 2854
rect 484308 2790 484360 2796
rect 484320 1630 484348 2790
rect 484412 2689 484440 4134
rect 486700 3392 486752 3398
rect 486700 3334 486752 3340
rect 484398 2680 484454 2689
rect 484398 2615 484454 2624
rect 484308 1624 484360 1630
rect 484308 1566 484360 1572
rect 486712 800 486740 3334
rect 487356 1834 487384 4134
rect 490392 2582 490420 4134
rect 492036 3324 492088 3330
rect 492036 3266 492088 3272
rect 490380 2576 490432 2582
rect 490380 2518 490432 2524
rect 487344 1828 487396 1834
rect 487344 1770 487396 1776
rect 492048 800 492076 3266
rect 493428 1902 493456 4134
rect 496832 1970 496860 4134
rect 497372 3256 497424 3262
rect 497372 3198 497424 3204
rect 496820 1964 496872 1970
rect 496820 1906 496872 1912
rect 493416 1896 493468 1902
rect 493416 1838 493468 1844
rect 497384 800 497412 3198
rect 499684 2650 499712 4134
rect 502616 3188 502668 3194
rect 502616 3130 502668 3136
rect 499672 2644 499724 2650
rect 499672 2586 499724 2592
rect 502628 1578 502656 3130
rect 502720 2514 502748 4134
rect 502708 2508 502760 2514
rect 502708 2450 502760 2456
rect 505756 2446 505784 4134
rect 505744 2440 505796 2446
rect 505744 2382 505796 2388
rect 508884 2106 508912 4134
rect 512012 2242 512040 4134
rect 512000 2236 512052 2242
rect 512000 2178 512052 2184
rect 515048 2174 515076 4134
rect 518084 2961 518112 4134
rect 518624 3324 518676 3330
rect 518624 3266 518676 3272
rect 518070 2952 518126 2961
rect 518070 2887 518126 2896
rect 515036 2168 515088 2174
rect 515036 2110 515088 2116
rect 508872 2100 508924 2106
rect 508872 2042 508924 2048
rect 513380 1760 513432 1766
rect 513380 1702 513432 1708
rect 508044 1692 508096 1698
rect 508044 1634 508096 1640
rect 502628 1550 502748 1578
rect 502720 800 502748 1550
rect 508056 800 508084 1634
rect 513392 800 513420 1702
rect 518636 800 518664 3266
rect 520292 2825 520320 153274
rect 520464 153264 520516 153270
rect 520464 153206 520516 153212
rect 520372 151360 520424 151366
rect 520372 151302 520424 151308
rect 520278 2816 520334 2825
rect 520278 2751 520334 2760
rect 520384 2310 520412 151302
rect 520476 5137 520504 153206
rect 521948 152454 521976 159200
rect 522868 153746 522896 159200
rect 523880 156602 523908 159200
rect 523868 156596 523920 156602
rect 523868 156538 523920 156544
rect 524892 153814 524920 159200
rect 524880 153808 524932 153814
rect 524880 153750 524932 153756
rect 522856 153740 522908 153746
rect 522856 153682 522908 153688
rect 523040 153468 523092 153474
rect 523040 153410 523092 153416
rect 521936 152448 521988 152454
rect 521936 152390 521988 152396
rect 520556 151836 520608 151842
rect 520556 151778 520608 151784
rect 520462 5128 520518 5137
rect 520462 5063 520518 5072
rect 520568 3330 520596 151778
rect 520648 151292 520700 151298
rect 520648 151234 520700 151240
rect 520556 3324 520608 3330
rect 520556 3266 520608 3272
rect 520660 2378 520688 151234
rect 521752 151156 521804 151162
rect 521752 151098 521804 151104
rect 521658 148200 521714 148209
rect 521658 148135 521714 148144
rect 520738 133376 520794 133385
rect 520738 133311 520794 133320
rect 520752 5098 520780 133311
rect 520830 37224 520886 37233
rect 520830 37159 520886 37168
rect 520740 5092 520792 5098
rect 520740 5034 520792 5040
rect 520648 2372 520700 2378
rect 520648 2314 520700 2320
rect 520372 2304 520424 2310
rect 520372 2246 520424 2252
rect 520844 1494 520872 37159
rect 520922 15056 520978 15065
rect 520922 14991 520978 15000
rect 520936 5302 520964 14991
rect 520924 5296 520976 5302
rect 520924 5238 520976 5244
rect 521672 4729 521700 148135
rect 521764 140865 521792 151098
rect 521844 151020 521896 151026
rect 521844 150962 521896 150968
rect 521750 140856 521806 140865
rect 521750 140791 521806 140800
rect 521750 126032 521806 126041
rect 521750 125967 521806 125976
rect 521764 5273 521792 125967
rect 521856 118697 521884 150962
rect 522304 150952 522356 150958
rect 522304 150894 522356 150900
rect 521842 118688 521898 118697
rect 521842 118623 521898 118632
rect 521842 111208 521898 111217
rect 521842 111143 521898 111152
rect 521750 5264 521806 5273
rect 521750 5199 521806 5208
rect 521856 5030 521884 111143
rect 521934 103864 521990 103873
rect 521934 103799 521990 103808
rect 521844 5024 521896 5030
rect 521948 5001 521976 103799
rect 522026 96384 522082 96393
rect 522026 96319 522082 96328
rect 521844 4966 521896 4972
rect 521934 4992 521990 5001
rect 521934 4927 521990 4936
rect 522040 4894 522068 96319
rect 522118 89040 522174 89049
rect 522118 88975 522174 88984
rect 522028 4888 522080 4894
rect 522028 4830 522080 4836
rect 521658 4720 521714 4729
rect 521658 4655 521714 4664
rect 522132 2922 522160 88975
rect 522210 81696 522266 81705
rect 522210 81631 522266 81640
rect 522224 4146 522252 81631
rect 522316 74225 522344 150894
rect 522302 74216 522358 74225
rect 522302 74151 522358 74160
rect 522580 52420 522632 52426
rect 522580 52362 522632 52368
rect 522592 52057 522620 52362
rect 522578 52048 522634 52057
rect 522578 51983 522634 51992
rect 522394 22400 522450 22409
rect 522394 22335 522450 22344
rect 522408 4826 522436 22335
rect 522946 7712 523002 7721
rect 522946 7647 523002 7656
rect 522396 4820 522448 4826
rect 522396 4762 522448 4768
rect 522212 4140 522264 4146
rect 522212 4082 522264 4088
rect 522960 3466 522988 7647
rect 523052 4865 523080 153410
rect 525812 153202 525840 159200
rect 526824 154562 526852 159200
rect 527744 157350 527772 159200
rect 527732 157344 527784 157350
rect 527732 157286 527784 157292
rect 528756 155786 528784 159200
rect 529768 157282 529796 159200
rect 529756 157276 529808 157282
rect 529756 157218 529808 157224
rect 530688 157146 530716 159200
rect 530676 157140 530728 157146
rect 530676 157082 530728 157088
rect 528744 155780 528796 155786
rect 528744 155722 528796 155728
rect 526812 154556 526864 154562
rect 526812 154498 526864 154504
rect 525800 153196 525852 153202
rect 525800 153138 525852 153144
rect 531700 153066 531728 159200
rect 532620 153134 532648 159200
rect 533632 157078 533660 159200
rect 533620 157072 533672 157078
rect 533620 157014 533672 157020
rect 534644 157010 534672 159200
rect 534632 157004 534684 157010
rect 534632 156946 534684 156952
rect 535564 156777 535592 159200
rect 535550 156768 535606 156777
rect 535550 156703 535606 156712
rect 536576 155718 536604 159200
rect 536564 155712 536616 155718
rect 536564 155654 536616 155660
rect 532608 153128 532660 153134
rect 532608 153070 532660 153076
rect 531688 153060 531740 153066
rect 531688 153002 531740 153008
rect 537496 152998 537524 159200
rect 538508 155650 538536 159200
rect 539520 156942 539548 159200
rect 540440 157214 540468 159200
rect 540428 157208 540480 157214
rect 540428 157150 540480 157156
rect 539508 156936 539560 156942
rect 539508 156878 539560 156884
rect 541452 156641 541480 159200
rect 541438 156632 541494 156641
rect 541438 156567 541494 156576
rect 538496 155644 538548 155650
rect 538496 155586 538548 155592
rect 542372 155582 542400 159200
rect 542360 155576 542412 155582
rect 542360 155518 542412 155524
rect 537484 152992 537536 152998
rect 537484 152934 537536 152940
rect 543384 152930 543412 159200
rect 544304 155446 544332 159200
rect 545316 156874 545344 159200
rect 545304 156868 545356 156874
rect 545304 156810 545356 156816
rect 546328 155514 546356 159200
rect 546316 155508 546368 155514
rect 546316 155450 546368 155456
rect 544292 155440 544344 155446
rect 544292 155382 544344 155388
rect 543372 152924 543424 152930
rect 543372 152866 543424 152872
rect 547248 152862 547276 159200
rect 547236 152856 547288 152862
rect 547236 152798 547288 152804
rect 548260 152794 548288 159200
rect 549180 156806 549208 159200
rect 549168 156800 549220 156806
rect 549168 156742 549220 156748
rect 550192 154494 550220 159200
rect 550180 154488 550232 154494
rect 550180 154430 550232 154436
rect 548248 152788 548300 152794
rect 548248 152730 548300 152736
rect 551204 152726 551232 159200
rect 552124 155378 552152 159200
rect 552112 155372 552164 155378
rect 552112 155314 552164 155320
rect 551192 152720 551244 152726
rect 551192 152662 551244 152668
rect 553136 152658 553164 159200
rect 554056 155961 554084 159200
rect 555068 156738 555096 159200
rect 555056 156732 555108 156738
rect 555056 156674 555108 156680
rect 554042 155952 554098 155961
rect 554042 155887 554098 155896
rect 556080 154426 556108 159200
rect 557000 156670 557028 159200
rect 556988 156664 557040 156670
rect 556988 156606 557040 156612
rect 558012 155689 558040 159200
rect 557998 155680 558054 155689
rect 557998 155615 558054 155624
rect 558932 154578 558960 159200
rect 558840 154550 558960 154578
rect 556068 154420 556120 154426
rect 556068 154362 556120 154368
rect 553124 152652 553176 152658
rect 553124 152594 553176 152600
rect 558840 152590 558868 154550
rect 559944 154358 559972 159200
rect 559932 154352 559984 154358
rect 559932 154294 559984 154300
rect 560956 154290 560984 159200
rect 561876 155553 561904 159200
rect 562888 155825 562916 159200
rect 562874 155816 562930 155825
rect 562874 155751 562930 155760
rect 561862 155544 561918 155553
rect 561862 155479 561918 155488
rect 563808 154970 563836 159200
rect 564820 155417 564848 159200
rect 564806 155408 564862 155417
rect 564806 155343 564862 155352
rect 561680 154964 561732 154970
rect 561680 154906 561732 154912
rect 563796 154964 563848 154970
rect 563796 154906 563848 154912
rect 560944 154284 560996 154290
rect 560944 154226 560996 154232
rect 561692 154222 561720 154906
rect 565832 154578 565860 159200
rect 565740 154550 565860 154578
rect 561680 154216 561732 154222
rect 561680 154158 561732 154164
rect 565740 154154 565768 154550
rect 565728 154148 565780 154154
rect 565728 154090 565780 154096
rect 558828 152584 558880 152590
rect 558828 152526 558880 152532
rect 566752 152522 566780 159200
rect 567764 154086 567792 159200
rect 568684 155281 568712 159200
rect 569696 155310 569724 159200
rect 569684 155304 569736 155310
rect 568670 155272 568726 155281
rect 569684 155246 569736 155252
rect 568670 155207 568726 155216
rect 567752 154080 567804 154086
rect 567752 154022 567804 154028
rect 570708 154018 570736 159200
rect 570696 154012 570748 154018
rect 570696 153954 570748 153960
rect 571628 153882 571656 159200
rect 572640 155242 572668 159200
rect 572628 155236 572680 155242
rect 572628 155178 572680 155184
rect 573560 153950 573588 159200
rect 574572 155922 574600 159200
rect 574560 155916 574612 155922
rect 574560 155858 574612 155864
rect 575480 155576 575532 155582
rect 575480 155518 575532 155524
rect 573548 153944 573600 153950
rect 573548 153886 573600 153892
rect 571616 153876 571668 153882
rect 571616 153818 571668 153824
rect 566740 152516 566792 152522
rect 566740 152458 566792 152464
rect 528560 151700 528612 151706
rect 528560 151642 528612 151648
rect 528572 16574 528600 151642
rect 545120 151564 545172 151570
rect 545120 151506 545172 151512
rect 545132 16574 545160 151506
rect 575492 151502 575520 155518
rect 575480 151496 575532 151502
rect 575480 151438 575532 151444
rect 575584 151434 575612 159200
rect 576504 155582 576532 159200
rect 576492 155576 576544 155582
rect 576492 155518 576544 155524
rect 575572 151428 575624 151434
rect 575572 151370 575624 151376
rect 528572 16546 528968 16574
rect 545132 16546 545344 16574
rect 523038 4856 523094 4865
rect 523038 4791 523094 4800
rect 522948 3460 523000 3466
rect 522948 3402 523000 3408
rect 522120 2916 522172 2922
rect 522120 2858 522172 2864
rect 523960 2848 524012 2854
rect 523960 2790 524012 2796
rect 520832 1488 520884 1494
rect 520832 1430 520884 1436
rect 523972 800 524000 2790
rect 417344 734 417556 762
rect 417606 0 417662 800
rect 422850 0 422906 800
rect 428186 0 428242 800
rect 433522 0 433578 800
rect 438858 0 438914 800
rect 444194 0 444250 800
rect 449530 0 449586 800
rect 454774 0 454830 800
rect 460110 0 460166 800
rect 465446 0 465502 800
rect 470782 0 470838 800
rect 476118 0 476174 800
rect 481454 0 481510 800
rect 486698 0 486754 800
rect 492034 0 492090 800
rect 497370 0 497426 800
rect 502706 0 502762 800
rect 508042 0 508098 800
rect 513378 0 513434 800
rect 518622 0 518678 800
rect 523958 0 524014 800
rect 528940 762 528968 16546
rect 534632 3800 534684 3806
rect 534632 3742 534684 3748
rect 529216 870 529336 898
rect 529216 762 529244 870
rect 529308 800 529336 870
rect 534644 800 534672 3742
rect 539968 3732 540020 3738
rect 539968 3674 540020 3680
rect 539980 800 540008 3674
rect 545316 800 545344 16546
rect 576872 5166 576900 159310
rect 577424 159202 577452 159310
rect 577502 159202 577558 160000
rect 577424 159200 577558 159202
rect 578422 159200 578478 160000
rect 579434 159200 579490 160000
rect 577424 159174 577544 159200
rect 578436 155582 578464 159200
rect 578424 155576 578476 155582
rect 578424 155518 578476 155524
rect 579448 152425 579476 159200
rect 579434 152416 579490 152425
rect 579434 152351 579490 152360
rect 576860 5160 576912 5166
rect 576860 5102 576912 5108
rect 577228 4956 577280 4962
rect 577228 4898 577280 4904
rect 555884 3868 555936 3874
rect 555884 3810 555936 3816
rect 550548 3120 550600 3126
rect 550548 3062 550600 3068
rect 550560 800 550588 3062
rect 555896 800 555924 3810
rect 566556 3460 566608 3466
rect 566556 3402 566608 3408
rect 561220 3052 561272 3058
rect 561220 2994 561272 3000
rect 561232 800 561260 2994
rect 566568 800 566596 3402
rect 571892 2984 571944 2990
rect 571892 2926 571944 2932
rect 571904 800 571932 2926
rect 577240 800 577268 4898
rect 528940 734 529244 762
rect 529294 0 529350 800
rect 534630 0 534686 800
rect 539966 0 540022 800
rect 545302 0 545358 800
rect 550546 0 550602 800
rect 555882 0 555938 800
rect 561218 0 561274 800
rect 566554 0 566610 800
rect 571890 0 571946 800
rect 577226 0 577282 800
<< via2 >>
rect 3422 157528 3478 157584
rect 3330 156576 3386 156632
rect 3054 148416 3110 148472
rect 5998 153176 6054 153232
rect 3514 152904 3570 152960
rect 3514 152224 3570 152280
rect 8206 155216 8262 155272
rect 13082 154264 13138 154320
rect 19890 155352 19946 155408
rect 25778 156712 25834 156768
rect 28722 154400 28778 154456
rect 30010 153448 30066 153504
rect 26606 153312 26662 153368
rect 33506 151952 33562 152008
rect 57518 153584 57574 153640
rect 50158 152632 50214 152688
rect 37462 152496 37518 152552
rect 61842 156848 61898 156904
rect 63774 155488 63830 155544
rect 67730 155624 67786 155680
rect 65706 152768 65762 152824
rect 79414 155896 79470 155952
rect 67500 152088 67556 152144
rect 81346 156984 81402 157040
rect 85026 153856 85082 153912
rect 81162 153720 81218 153776
rect 87142 155760 87198 155816
rect 94042 152904 94098 152960
rect 98826 153992 98882 154048
rect 101770 157120 101826 157176
rect 106646 155080 106702 155136
rect 102782 154808 102838 154864
rect 109590 154672 109646 154728
rect 114466 154944 114522 155000
rect 112534 154128 112590 154184
rect 113822 152088 113878 152144
rect 102046 151816 102102 151872
rect 71318 151408 71374 151464
rect 9402 151272 9458 151328
rect 12806 151272 12862 151328
rect 16302 151272 16358 151328
rect 19706 151272 19762 151328
rect 47030 151272 47086 151328
rect 53930 151272 53986 151328
rect 60830 151272 60886 151328
rect 3330 149912 3386 149968
rect 3238 139304 3294 139360
rect 3422 143792 3478 143848
rect 3330 134680 3386 134736
rect 4066 130056 4122 130112
rect 3974 125568 4030 125624
rect 3882 120944 3938 121000
rect 3790 116456 3846 116512
rect 3698 111832 3754 111888
rect 3606 107208 3662 107264
rect 3514 102720 3570 102776
rect 3422 98096 3478 98152
rect 3698 93608 3754 93664
rect 3422 84360 3478 84416
rect 3330 57024 3386 57080
rect 3238 52400 3294 52456
rect 3146 47912 3202 47968
rect 3054 43288 3110 43344
rect 2962 38664 3018 38720
rect 2870 34176 2926 34232
rect 3514 70760 3570 70816
rect 3422 15816 3478 15872
rect 3238 6704 3294 6760
rect 3606 66136 3662 66192
rect 3790 88984 3846 89040
rect 4066 79872 4122 79928
rect 3974 75248 4030 75304
rect 3882 61512 3938 61568
rect 3698 29552 3754 29608
rect 3790 25064 3846 25120
rect 4066 20440 4122 20496
rect 3974 11328 4030 11384
rect 4986 6024 5042 6080
rect 5446 5888 5502 5944
rect 35806 4528 35862 4584
rect 65982 4528 66038 4584
rect 71962 4528 72018 4584
rect 72422 4528 72478 4584
rect 74906 4528 74962 4584
rect 81990 4528 82046 4584
rect 82174 4528 82230 4584
rect 82634 4528 82690 4584
rect 82818 4528 82874 4584
rect 86406 4528 86462 4584
rect 102690 4528 102746 4584
rect 2962 2216 3018 2272
rect 49330 2760 49386 2816
rect 112534 5888 112590 5944
rect 114926 152224 114982 152280
rect 114098 151272 114154 151328
rect 113914 2896 113970 2952
rect 115018 6024 115074 6080
rect 115478 151952 115534 152008
rect 115294 151816 115350 151872
rect 115202 3032 115258 3088
rect 118238 152360 118294 152416
rect 116582 151408 116638 151464
rect 115662 150592 115718 150648
rect 115478 2352 115534 2408
rect 116306 100544 116362 100600
rect 116306 66408 116362 66464
rect 116490 20868 116546 20904
rect 116490 20848 116492 20868
rect 116492 20848 116544 20868
rect 116544 20848 116546 20868
rect 115662 1944 115718 2000
rect 116674 141616 116730 141672
rect 116766 134680 116822 134736
rect 116858 123256 116914 123312
rect 116950 111968 117006 112024
rect 116950 109792 117006 109848
rect 118146 150728 118202 150784
rect 117962 150456 118018 150512
rect 117134 146104 117190 146160
rect 117870 150320 117926 150376
rect 117318 147464 117374 147520
rect 117226 144744 117282 144800
rect 117686 136448 117742 136504
rect 117594 132912 117650 132968
rect 117318 130056 117374 130112
rect 117318 124228 117374 124264
rect 117318 124208 117320 124228
rect 117320 124208 117372 124228
rect 117372 124208 117374 124228
rect 117502 104624 117558 104680
rect 117042 98776 117098 98832
rect 117502 95920 117558 95976
rect 117318 86808 117374 86864
rect 117318 83816 117374 83872
rect 117318 72664 117374 72720
rect 117318 66952 117374 67008
rect 117318 57568 117374 57624
rect 117318 51720 117374 51776
rect 117410 48864 117466 48920
rect 117318 45872 117374 45928
rect 117318 43016 117374 43072
rect 117226 37168 117282 37224
rect 117134 34312 117190 34368
rect 117042 32272 117098 32328
rect 116950 9560 117006 9616
rect 117318 31456 117374 31512
rect 117502 16904 117558 16960
rect 117318 14048 117374 14104
rect 117318 11076 117374 11112
rect 117318 11056 117320 11076
rect 117320 11056 117372 11076
rect 117372 11056 117374 11076
rect 117318 8200 117374 8256
rect 117318 5344 117374 5400
rect 117870 101768 117926 101824
rect 117686 81368 117742 81424
rect 117686 78512 117742 78568
rect 117870 69808 117926 69864
rect 117870 63280 117926 63336
rect 117870 40160 117926 40216
rect 117870 22752 117926 22808
rect 117778 19760 117834 19816
rect 118054 138760 118110 138816
rect 120354 157256 120410 157312
rect 121918 156576 121974 156632
rect 125138 155216 125194 155272
rect 126150 154536 126206 154592
rect 128358 154264 128414 154320
rect 131210 155352 131266 155408
rect 131302 154536 131358 154592
rect 132774 155352 132830 155408
rect 136822 156712 136878 156768
rect 138202 155352 138258 155408
rect 138846 154400 138902 154456
rect 144918 152496 144974 152552
rect 119894 151816 119950 151872
rect 153198 152632 153254 152688
rect 154486 156576 154542 156632
rect 158810 155488 158866 155544
rect 160098 155624 160154 155680
rect 160926 156848 160982 156904
rect 161294 155216 161350 155272
rect 164054 155896 164110 155952
rect 163502 152768 163558 152824
rect 118238 127880 118294 127936
rect 118238 121352 118294 121408
rect 118330 118632 118386 118688
rect 118514 149912 118570 149968
rect 118422 115776 118478 115832
rect 118422 112648 118478 112704
rect 118146 2080 118202 2136
rect 118698 106800 118754 106856
rect 118606 92384 118662 92440
rect 118514 89664 118570 89720
rect 118606 75656 118662 75712
rect 118606 60424 118662 60480
rect 118514 54576 118570 54632
rect 118514 28464 118570 28520
rect 118606 25608 118662 25664
rect 119618 151136 119674 151192
rect 119434 150864 119490 150920
rect 119434 2216 119490 2272
rect 119802 151000 119858 151056
rect 173898 156984 173954 157040
rect 171966 155352 172022 155408
rect 174910 154536 174966 154592
rect 178130 155760 178186 155816
rect 175922 154672 175978 154728
rect 178222 154536 178278 154592
rect 179510 154808 179566 154864
rect 182362 152904 182418 152960
rect 187698 157120 187754 157176
rect 190826 155080 190882 155136
rect 194230 154844 194232 154864
rect 194232 154844 194284 154864
rect 194284 154844 194286 154864
rect 194230 154808 194286 154844
rect 196070 154944 196126 155000
rect 199106 154808 199162 154864
rect 200394 157256 200450 157312
rect 201958 155916 202014 155952
rect 201958 155896 201960 155916
rect 201960 155896 202012 155916
rect 202012 155896 202014 155916
rect 203246 155896 203302 155952
rect 214838 155488 214894 155544
rect 218794 155624 218850 155680
rect 219254 154572 219256 154592
rect 219256 154572 219308 154592
rect 219308 154572 219310 154592
rect 219254 154536 219310 154572
rect 219622 154536 219678 154592
rect 222750 156576 222806 156632
rect 227258 155216 227314 155272
rect 230478 155216 230534 155272
rect 234342 155760 234398 155816
rect 234618 155352 234674 155408
rect 243450 154944 243506 155000
rect 249798 154944 249854 155000
rect 260930 155488 260986 155544
rect 261666 155352 261722 155408
rect 262218 155624 262274 155680
rect 273166 155216 273222 155272
rect 274362 155216 274418 155272
rect 275834 155760 275890 155816
rect 277122 154808 277178 154864
rect 277490 154808 277546 154864
rect 279146 154808 279202 154864
rect 282366 154808 282422 154864
rect 293866 155352 293922 155408
rect 302698 155216 302754 155272
rect 436006 155216 436062 155272
rect 473174 155216 473230 155272
rect 477314 156712 477370 156768
rect 481546 156576 481602 156632
rect 489642 155896 489698 155952
rect 492586 155624 492642 155680
rect 495254 155488 495310 155544
rect 495898 155760 495954 155816
rect 497186 155352 497242 155408
rect 499394 155216 499450 155272
rect 505650 153176 505706 153232
rect 509514 153312 509570 153368
rect 513470 153584 513526 153640
rect 517518 153992 517574 154048
rect 516690 153856 516746 153912
rect 516138 153720 516194 153776
rect 510894 153448 510950 153504
rect 519266 154128 519322 154184
rect 508226 151816 508282 151872
rect 119618 2624 119674 2680
rect 118330 1808 118386 1864
rect 119986 2488 120042 2544
rect 447322 1808 447378 1864
rect 450358 1944 450414 2000
rect 456798 2080 456854 2136
rect 465722 2216 465778 2272
rect 475014 3032 475070 3088
rect 471978 2352 472034 2408
rect 481178 2488 481234 2544
rect 484398 2624 484454 2680
rect 518070 2896 518126 2952
rect 520278 2760 520334 2816
rect 520462 5072 520518 5128
rect 521658 148144 521714 148200
rect 520738 133320 520794 133376
rect 520830 37168 520886 37224
rect 520922 15000 520978 15056
rect 521750 140800 521806 140856
rect 521750 125976 521806 126032
rect 521842 118632 521898 118688
rect 521842 111152 521898 111208
rect 521750 5208 521806 5264
rect 521934 103808 521990 103864
rect 522026 96328 522082 96384
rect 521934 4936 521990 4992
rect 522118 88984 522174 89040
rect 521658 4664 521714 4720
rect 522210 81640 522266 81696
rect 522302 74160 522358 74216
rect 522578 51992 522634 52048
rect 522394 22344 522450 22400
rect 522946 7656 523002 7712
rect 535550 156712 535606 156768
rect 541438 156576 541494 156632
rect 554042 155896 554098 155952
rect 557998 155624 558054 155680
rect 562874 155760 562930 155816
rect 561862 155488 561918 155544
rect 564806 155352 564862 155408
rect 568670 155216 568726 155272
rect 523038 4800 523094 4856
rect 579434 152360 579490 152416
<< metal3 >>
rect 0 157586 800 157616
rect 3417 157586 3483 157589
rect 0 157584 3483 157586
rect 0 157528 3422 157584
rect 3478 157528 3483 157584
rect 0 157526 3483 157528
rect 0 157496 800 157526
rect 3417 157523 3483 157526
rect 120349 157314 120415 157317
rect 200389 157314 200455 157317
rect 120349 157312 200455 157314
rect 120349 157256 120354 157312
rect 120410 157256 200394 157312
rect 200450 157256 200455 157312
rect 120349 157254 200455 157256
rect 120349 157251 120415 157254
rect 200389 157251 200455 157254
rect 101765 157178 101831 157181
rect 187693 157178 187759 157181
rect 101765 157176 187759 157178
rect 101765 157120 101770 157176
rect 101826 157120 187698 157176
rect 187754 157120 187759 157176
rect 101765 157118 187759 157120
rect 101765 157115 101831 157118
rect 187693 157115 187759 157118
rect 81341 157042 81407 157045
rect 173893 157042 173959 157045
rect 81341 157040 173959 157042
rect 81341 156984 81346 157040
rect 81402 156984 173898 157040
rect 173954 156984 173959 157040
rect 81341 156982 173959 156984
rect 81341 156979 81407 156982
rect 173893 156979 173959 156982
rect 61837 156906 61903 156909
rect 160921 156906 160987 156909
rect 61837 156904 160987 156906
rect 61837 156848 61842 156904
rect 61898 156848 160926 156904
rect 160982 156848 160987 156904
rect 61837 156846 160987 156848
rect 61837 156843 61903 156846
rect 160921 156843 160987 156846
rect 25773 156770 25839 156773
rect 136817 156770 136883 156773
rect 25773 156768 136883 156770
rect 25773 156712 25778 156768
rect 25834 156712 136822 156768
rect 136878 156712 136883 156768
rect 25773 156710 136883 156712
rect 25773 156707 25839 156710
rect 136817 156707 136883 156710
rect 477309 156770 477375 156773
rect 535545 156770 535611 156773
rect 477309 156768 535611 156770
rect 477309 156712 477314 156768
rect 477370 156712 535550 156768
rect 535606 156712 535611 156768
rect 477309 156710 535611 156712
rect 477309 156707 477375 156710
rect 535545 156707 535611 156710
rect 3325 156634 3391 156637
rect 121913 156634 121979 156637
rect 3325 156632 121979 156634
rect 3325 156576 3330 156632
rect 3386 156576 121918 156632
rect 121974 156576 121979 156632
rect 3325 156574 121979 156576
rect 3325 156571 3391 156574
rect 121913 156571 121979 156574
rect 154481 156634 154547 156637
rect 222745 156634 222811 156637
rect 154481 156632 222811 156634
rect 154481 156576 154486 156632
rect 154542 156576 222750 156632
rect 222806 156576 222811 156632
rect 154481 156574 222811 156576
rect 154481 156571 154547 156574
rect 222745 156571 222811 156574
rect 481541 156634 481607 156637
rect 541433 156634 541499 156637
rect 481541 156632 541499 156634
rect 481541 156576 481546 156632
rect 481602 156576 541438 156632
rect 541494 156576 541499 156632
rect 481541 156574 541499 156576
rect 481541 156571 481607 156574
rect 541433 156571 541499 156574
rect 79409 155954 79475 155957
rect 164049 155954 164115 155957
rect 79409 155952 164115 155954
rect 79409 155896 79414 155952
rect 79470 155896 164054 155952
rect 164110 155896 164115 155952
rect 79409 155894 164115 155896
rect 79409 155891 79475 155894
rect 164049 155891 164115 155894
rect 201953 155954 202019 155957
rect 203241 155954 203307 155957
rect 201953 155952 203307 155954
rect 201953 155896 201958 155952
rect 202014 155896 203246 155952
rect 203302 155896 203307 155952
rect 201953 155894 203307 155896
rect 201953 155891 202019 155894
rect 203241 155891 203307 155894
rect 489637 155954 489703 155957
rect 554037 155954 554103 155957
rect 489637 155952 554103 155954
rect 489637 155896 489642 155952
rect 489698 155896 554042 155952
rect 554098 155896 554103 155952
rect 489637 155894 554103 155896
rect 489637 155891 489703 155894
rect 554037 155891 554103 155894
rect 87137 155818 87203 155821
rect 178125 155818 178191 155821
rect 87137 155816 178191 155818
rect 87137 155760 87142 155816
rect 87198 155760 178130 155816
rect 178186 155760 178191 155816
rect 87137 155758 178191 155760
rect 87137 155755 87203 155758
rect 178125 155755 178191 155758
rect 234337 155818 234403 155821
rect 275829 155818 275895 155821
rect 234337 155816 275895 155818
rect 234337 155760 234342 155816
rect 234398 155760 275834 155816
rect 275890 155760 275895 155816
rect 234337 155758 275895 155760
rect 234337 155755 234403 155758
rect 275829 155755 275895 155758
rect 495893 155818 495959 155821
rect 562869 155818 562935 155821
rect 495893 155816 562935 155818
rect 495893 155760 495898 155816
rect 495954 155760 562874 155816
rect 562930 155760 562935 155816
rect 495893 155758 562935 155760
rect 495893 155755 495959 155758
rect 562869 155755 562935 155758
rect 67725 155682 67791 155685
rect 160093 155682 160159 155685
rect 67725 155680 160159 155682
rect 67725 155624 67730 155680
rect 67786 155624 160098 155680
rect 160154 155624 160159 155680
rect 67725 155622 160159 155624
rect 67725 155619 67791 155622
rect 160093 155619 160159 155622
rect 218789 155682 218855 155685
rect 262213 155682 262279 155685
rect 218789 155680 262279 155682
rect 218789 155624 218794 155680
rect 218850 155624 262218 155680
rect 262274 155624 262279 155680
rect 218789 155622 262279 155624
rect 218789 155619 218855 155622
rect 262213 155619 262279 155622
rect 492581 155682 492647 155685
rect 557993 155682 558059 155685
rect 492581 155680 558059 155682
rect 492581 155624 492586 155680
rect 492642 155624 557998 155680
rect 558054 155624 558059 155680
rect 492581 155622 558059 155624
rect 492581 155619 492647 155622
rect 557993 155619 558059 155622
rect 63769 155546 63835 155549
rect 158805 155546 158871 155549
rect 63769 155544 158871 155546
rect 63769 155488 63774 155544
rect 63830 155488 158810 155544
rect 158866 155488 158871 155544
rect 63769 155486 158871 155488
rect 63769 155483 63835 155486
rect 158805 155483 158871 155486
rect 214833 155546 214899 155549
rect 260925 155546 260991 155549
rect 214833 155544 260991 155546
rect 214833 155488 214838 155544
rect 214894 155488 260930 155544
rect 260986 155488 260991 155544
rect 214833 155486 260991 155488
rect 214833 155483 214899 155486
rect 260925 155483 260991 155486
rect 495249 155546 495315 155549
rect 561857 155546 561923 155549
rect 495249 155544 561923 155546
rect 495249 155488 495254 155544
rect 495310 155488 561862 155544
rect 561918 155488 561923 155544
rect 495249 155486 561923 155488
rect 495249 155483 495315 155486
rect 561857 155483 561923 155486
rect 19885 155410 19951 155413
rect 131205 155410 131271 155413
rect 19885 155408 131271 155410
rect 19885 155352 19890 155408
rect 19946 155352 131210 155408
rect 131266 155352 131271 155408
rect 19885 155350 131271 155352
rect 19885 155347 19951 155350
rect 131205 155347 131271 155350
rect 132769 155410 132835 155413
rect 138197 155410 138263 155413
rect 132769 155408 138263 155410
rect 132769 155352 132774 155408
rect 132830 155352 138202 155408
rect 138258 155352 138263 155408
rect 132769 155350 138263 155352
rect 132769 155347 132835 155350
rect 138197 155347 138263 155350
rect 171961 155410 172027 155413
rect 234613 155410 234679 155413
rect 171961 155408 234679 155410
rect 171961 155352 171966 155408
rect 172022 155352 234618 155408
rect 234674 155352 234679 155408
rect 171961 155350 234679 155352
rect 171961 155347 172027 155350
rect 234613 155347 234679 155350
rect 261661 155410 261727 155413
rect 293861 155410 293927 155413
rect 261661 155408 293927 155410
rect 261661 155352 261666 155408
rect 261722 155352 293866 155408
rect 293922 155352 293927 155408
rect 261661 155350 293927 155352
rect 261661 155347 261727 155350
rect 293861 155347 293927 155350
rect 497181 155410 497247 155413
rect 564801 155410 564867 155413
rect 497181 155408 564867 155410
rect 497181 155352 497186 155408
rect 497242 155352 564806 155408
rect 564862 155352 564867 155408
rect 497181 155350 564867 155352
rect 497181 155347 497247 155350
rect 564801 155347 564867 155350
rect 8201 155274 8267 155277
rect 125133 155274 125199 155277
rect 8201 155272 125199 155274
rect 8201 155216 8206 155272
rect 8262 155216 125138 155272
rect 125194 155216 125199 155272
rect 8201 155214 125199 155216
rect 8201 155211 8267 155214
rect 125133 155211 125199 155214
rect 161289 155274 161355 155277
rect 227253 155274 227319 155277
rect 161289 155272 227319 155274
rect 161289 155216 161294 155272
rect 161350 155216 227258 155272
rect 227314 155216 227319 155272
rect 161289 155214 227319 155216
rect 161289 155211 161355 155214
rect 227253 155211 227319 155214
rect 230473 155274 230539 155277
rect 273161 155274 273227 155277
rect 230473 155272 273227 155274
rect 230473 155216 230478 155272
rect 230534 155216 273166 155272
rect 273222 155216 273227 155272
rect 230473 155214 273227 155216
rect 230473 155211 230539 155214
rect 273161 155211 273227 155214
rect 274357 155274 274423 155277
rect 302693 155274 302759 155277
rect 274357 155272 302759 155274
rect 274357 155216 274362 155272
rect 274418 155216 302698 155272
rect 302754 155216 302759 155272
rect 274357 155214 302759 155216
rect 274357 155211 274423 155214
rect 302693 155211 302759 155214
rect 436001 155274 436067 155277
rect 473169 155274 473235 155277
rect 436001 155272 473235 155274
rect 436001 155216 436006 155272
rect 436062 155216 473174 155272
rect 473230 155216 473235 155272
rect 436001 155214 473235 155216
rect 436001 155211 436067 155214
rect 473169 155211 473235 155214
rect 499389 155274 499455 155277
rect 568665 155274 568731 155277
rect 499389 155272 568731 155274
rect 499389 155216 499394 155272
rect 499450 155216 568670 155272
rect 568726 155216 568731 155272
rect 499389 155214 568731 155216
rect 499389 155211 499455 155214
rect 568665 155211 568731 155214
rect 106641 155138 106707 155141
rect 190821 155138 190887 155141
rect 106641 155136 190887 155138
rect 106641 155080 106646 155136
rect 106702 155080 190826 155136
rect 190882 155080 190887 155136
rect 106641 155078 190887 155080
rect 106641 155075 106707 155078
rect 190821 155075 190887 155078
rect 114461 155002 114527 155005
rect 196065 155002 196131 155005
rect 114461 155000 196131 155002
rect 114461 154944 114466 155000
rect 114522 154944 196070 155000
rect 196126 154944 196131 155000
rect 114461 154942 196131 154944
rect 114461 154939 114527 154942
rect 196065 154939 196131 154942
rect 243445 155002 243511 155005
rect 249793 155002 249859 155005
rect 243445 155000 249859 155002
rect 243445 154944 243450 155000
rect 243506 154944 249798 155000
rect 249854 154944 249859 155000
rect 243445 154942 249859 154944
rect 243445 154939 243511 154942
rect 249793 154939 249859 154942
rect 102777 154866 102843 154869
rect 179505 154866 179571 154869
rect 102777 154864 179571 154866
rect 102777 154808 102782 154864
rect 102838 154808 179510 154864
rect 179566 154808 179571 154864
rect 102777 154806 179571 154808
rect 102777 154803 102843 154806
rect 179505 154803 179571 154806
rect 194225 154866 194291 154869
rect 199101 154866 199167 154869
rect 194225 154864 199167 154866
rect 194225 154808 194230 154864
rect 194286 154808 199106 154864
rect 199162 154808 199167 154864
rect 194225 154806 199167 154808
rect 194225 154803 194291 154806
rect 199101 154803 199167 154806
rect 277117 154866 277183 154869
rect 277485 154866 277551 154869
rect 277117 154864 277551 154866
rect 277117 154808 277122 154864
rect 277178 154808 277490 154864
rect 277546 154808 277551 154864
rect 277117 154806 277551 154808
rect 277117 154803 277183 154806
rect 277485 154803 277551 154806
rect 279141 154866 279207 154869
rect 282361 154866 282427 154869
rect 279141 154864 282427 154866
rect 279141 154808 279146 154864
rect 279202 154808 282366 154864
rect 282422 154808 282427 154864
rect 279141 154806 282427 154808
rect 279141 154803 279207 154806
rect 282361 154803 282427 154806
rect 109585 154730 109651 154733
rect 175917 154730 175983 154733
rect 109585 154728 175983 154730
rect 109585 154672 109590 154728
rect 109646 154672 175922 154728
rect 175978 154672 175983 154728
rect 109585 154670 175983 154672
rect 109585 154667 109651 154670
rect 175917 154667 175983 154670
rect 126145 154594 126211 154597
rect 131297 154594 131363 154597
rect 126145 154592 131363 154594
rect 126145 154536 126150 154592
rect 126206 154536 131302 154592
rect 131358 154536 131363 154592
rect 126145 154534 131363 154536
rect 126145 154531 126211 154534
rect 131297 154531 131363 154534
rect 174905 154594 174971 154597
rect 178217 154594 178283 154597
rect 174905 154592 178283 154594
rect 174905 154536 174910 154592
rect 174966 154536 178222 154592
rect 178278 154536 178283 154592
rect 174905 154534 178283 154536
rect 174905 154531 174971 154534
rect 178217 154531 178283 154534
rect 219249 154594 219315 154597
rect 219617 154594 219683 154597
rect 219249 154592 219683 154594
rect 219249 154536 219254 154592
rect 219310 154536 219622 154592
rect 219678 154536 219683 154592
rect 219249 154534 219683 154536
rect 219249 154531 219315 154534
rect 219617 154531 219683 154534
rect 28717 154458 28783 154461
rect 138841 154458 138907 154461
rect 28717 154456 138907 154458
rect 28717 154400 28722 154456
rect 28778 154400 138846 154456
rect 138902 154400 138907 154456
rect 28717 154398 138907 154400
rect 28717 154395 28783 154398
rect 138841 154395 138907 154398
rect 13077 154322 13143 154325
rect 128353 154322 128419 154325
rect 13077 154320 128419 154322
rect 13077 154264 13082 154320
rect 13138 154264 128358 154320
rect 128414 154264 128419 154320
rect 13077 154262 128419 154264
rect 13077 154259 13143 154262
rect 128353 154259 128419 154262
rect 112529 154186 112595 154189
rect 519261 154186 519327 154189
rect 112529 154184 519327 154186
rect 112529 154128 112534 154184
rect 112590 154128 519266 154184
rect 519322 154128 519327 154184
rect 112529 154126 519327 154128
rect 112529 154123 112595 154126
rect 519261 154123 519327 154126
rect 98821 154050 98887 154053
rect 517513 154050 517579 154053
rect 98821 154048 517579 154050
rect 98821 153992 98826 154048
rect 98882 153992 517518 154048
rect 517574 153992 517579 154048
rect 98821 153990 517579 153992
rect 98821 153987 98887 153990
rect 517513 153987 517579 153990
rect 85021 153914 85087 153917
rect 516685 153914 516751 153917
rect 85021 153912 516751 153914
rect 85021 153856 85026 153912
rect 85082 153856 516690 153912
rect 516746 153856 516751 153912
rect 85021 153854 516751 153856
rect 85021 153851 85087 153854
rect 516685 153851 516751 153854
rect 81157 153778 81223 153781
rect 516133 153778 516199 153781
rect 81157 153776 516199 153778
rect 81157 153720 81162 153776
rect 81218 153720 516138 153776
rect 516194 153720 516199 153776
rect 81157 153718 516199 153720
rect 81157 153715 81223 153718
rect 516133 153715 516199 153718
rect 57513 153642 57579 153645
rect 513465 153642 513531 153645
rect 57513 153640 513531 153642
rect 57513 153584 57518 153640
rect 57574 153584 513470 153640
rect 513526 153584 513531 153640
rect 57513 153582 513531 153584
rect 57513 153579 57579 153582
rect 513465 153579 513531 153582
rect 30005 153506 30071 153509
rect 510889 153506 510955 153509
rect 30005 153504 510955 153506
rect 30005 153448 30010 153504
rect 30066 153448 510894 153504
rect 510950 153448 510955 153504
rect 30005 153446 510955 153448
rect 30005 153443 30071 153446
rect 510889 153443 510955 153446
rect 26601 153370 26667 153373
rect 509509 153370 509575 153373
rect 26601 153368 509575 153370
rect 26601 153312 26606 153368
rect 26662 153312 509514 153368
rect 509570 153312 509575 153368
rect 26601 153310 509575 153312
rect 26601 153307 26667 153310
rect 509509 153307 509575 153310
rect 5993 153234 6059 153237
rect 505645 153234 505711 153237
rect 5993 153232 505711 153234
rect 5993 153176 5998 153232
rect 6054 153176 505650 153232
rect 505706 153176 505711 153232
rect 5993 153174 505711 153176
rect 5993 153171 6059 153174
rect 505645 153171 505711 153174
rect 0 152962 800 152992
rect 3509 152962 3575 152965
rect 0 152960 3575 152962
rect 0 152904 3514 152960
rect 3570 152904 3575 152960
rect 0 152902 3575 152904
rect 0 152872 800 152902
rect 3509 152899 3575 152902
rect 94037 152962 94103 152965
rect 182357 152962 182423 152965
rect 94037 152960 182423 152962
rect 94037 152904 94042 152960
rect 94098 152904 182362 152960
rect 182418 152904 182423 152960
rect 94037 152902 182423 152904
rect 94037 152899 94103 152902
rect 182357 152899 182423 152902
rect 65701 152826 65767 152829
rect 163497 152826 163563 152829
rect 65701 152824 163563 152826
rect 65701 152768 65706 152824
rect 65762 152768 163502 152824
rect 163558 152768 163563 152824
rect 65701 152766 163563 152768
rect 65701 152763 65767 152766
rect 163497 152763 163563 152766
rect 50153 152690 50219 152693
rect 153193 152690 153259 152693
rect 50153 152688 153259 152690
rect 50153 152632 50158 152688
rect 50214 152632 153198 152688
rect 153254 152632 153259 152688
rect 50153 152630 153259 152632
rect 50153 152627 50219 152630
rect 153193 152627 153259 152630
rect 37457 152554 37523 152557
rect 144913 152554 144979 152557
rect 37457 152552 144979 152554
rect 37457 152496 37462 152552
rect 37518 152496 144918 152552
rect 144974 152496 144979 152552
rect 37457 152494 144979 152496
rect 37457 152491 37523 152494
rect 144913 152491 144979 152494
rect 118233 152418 118299 152421
rect 579429 152418 579495 152421
rect 118233 152416 579495 152418
rect 118233 152360 118238 152416
rect 118294 152360 579434 152416
rect 579490 152360 579495 152416
rect 118233 152358 579495 152360
rect 118233 152355 118299 152358
rect 579429 152355 579495 152358
rect 3509 152282 3575 152285
rect 114921 152282 114987 152285
rect 3509 152280 114987 152282
rect 3509 152224 3514 152280
rect 3570 152224 114926 152280
rect 114982 152224 114987 152280
rect 3509 152222 114987 152224
rect 3509 152219 3575 152222
rect 114921 152219 114987 152222
rect 67495 152146 67561 152149
rect 113817 152146 113883 152149
rect 67495 152144 113883 152146
rect 67495 152088 67500 152144
rect 67556 152088 113822 152144
rect 113878 152088 113883 152144
rect 67495 152086 113883 152088
rect 67495 152083 67561 152086
rect 113817 152083 113883 152086
rect 33501 152010 33567 152013
rect 115473 152010 115539 152013
rect 33501 152008 115539 152010
rect 33501 151952 33506 152008
rect 33562 151952 115478 152008
rect 115534 151952 115539 152008
rect 33501 151950 115539 151952
rect 33501 151947 33567 151950
rect 115473 151947 115539 151950
rect 102041 151874 102107 151877
rect 115289 151874 115355 151877
rect 102041 151872 115355 151874
rect 102041 151816 102046 151872
rect 102102 151816 115294 151872
rect 115350 151816 115355 151872
rect 102041 151814 115355 151816
rect 102041 151811 102107 151814
rect 115289 151811 115355 151814
rect 119889 151874 119955 151877
rect 508221 151874 508287 151877
rect 119889 151872 508287 151874
rect 119889 151816 119894 151872
rect 119950 151816 508226 151872
rect 508282 151816 508287 151872
rect 119889 151814 508287 151816
rect 119889 151811 119955 151814
rect 508221 151811 508287 151814
rect 71313 151466 71379 151469
rect 116577 151466 116643 151469
rect 71313 151464 116643 151466
rect 71313 151408 71318 151464
rect 71374 151408 116582 151464
rect 116638 151408 116643 151464
rect 71313 151406 116643 151408
rect 71313 151403 71379 151406
rect 116577 151403 116643 151406
rect 9397 151330 9463 151333
rect 12801 151330 12867 151333
rect 16297 151330 16363 151333
rect 19701 151330 19767 151333
rect 47025 151330 47091 151333
rect 53925 151330 53991 151333
rect 60825 151330 60891 151333
rect 114093 151330 114159 151333
rect 9397 151328 12634 151330
rect 9397 151272 9402 151328
rect 9458 151272 12634 151328
rect 9397 151270 12634 151272
rect 9397 151267 9463 151270
rect 12574 150514 12634 151270
rect 12801 151328 14658 151330
rect 12801 151272 12806 151328
rect 12862 151272 14658 151328
rect 12801 151270 14658 151272
rect 12801 151267 12867 151270
rect 14598 150650 14658 151270
rect 16297 151328 16590 151330
rect 16297 151272 16302 151328
rect 16358 151272 16590 151328
rect 16297 151270 16590 151272
rect 16297 151267 16363 151270
rect 16530 150786 16590 151270
rect 19701 151328 26250 151330
rect 19701 151272 19706 151328
rect 19762 151272 26250 151328
rect 19701 151270 26250 151272
rect 19701 151267 19767 151270
rect 26190 150922 26250 151270
rect 47025 151328 51090 151330
rect 47025 151272 47030 151328
rect 47086 151272 51090 151328
rect 47025 151270 51090 151272
rect 47025 151267 47091 151270
rect 51030 151058 51090 151270
rect 53925 151328 55230 151330
rect 53925 151272 53930 151328
rect 53986 151272 55230 151328
rect 53925 151270 55230 151272
rect 53925 151267 53991 151270
rect 55170 151194 55230 151270
rect 60825 151328 114159 151330
rect 60825 151272 60830 151328
rect 60886 151272 114098 151328
rect 114154 151272 114159 151328
rect 60825 151270 114159 151272
rect 60825 151267 60891 151270
rect 114093 151267 114159 151270
rect 119613 151194 119679 151197
rect 55170 151192 119679 151194
rect 55170 151136 119618 151192
rect 119674 151136 119679 151192
rect 55170 151134 119679 151136
rect 119613 151131 119679 151134
rect 119797 151058 119863 151061
rect 51030 151056 119863 151058
rect 51030 151000 119802 151056
rect 119858 151000 119863 151056
rect 51030 150998 119863 151000
rect 119797 150995 119863 150998
rect 119429 150922 119495 150925
rect 26190 150920 119495 150922
rect 26190 150864 119434 150920
rect 119490 150864 119495 150920
rect 26190 150862 119495 150864
rect 119429 150859 119495 150862
rect 118141 150786 118207 150789
rect 16530 150784 118207 150786
rect 16530 150728 118146 150784
rect 118202 150728 118207 150784
rect 16530 150726 118207 150728
rect 118141 150723 118207 150726
rect 115657 150650 115723 150653
rect 14598 150648 115723 150650
rect 14598 150592 115662 150648
rect 115718 150592 115723 150648
rect 14598 150590 115723 150592
rect 115657 150587 115723 150590
rect 117957 150514 118023 150517
rect 12574 150512 118023 150514
rect 12574 150456 117962 150512
rect 118018 150456 118023 150512
rect 12574 150454 118023 150456
rect 117957 150451 118023 150454
rect 117865 150378 117931 150381
rect 117865 150376 120060 150378
rect 117865 150320 117870 150376
rect 117926 150320 120060 150376
rect 117865 150318 120060 150320
rect 117865 150315 117931 150318
rect 3325 149970 3391 149973
rect 118509 149970 118575 149973
rect 3325 149968 118575 149970
rect 3325 149912 3330 149968
rect 3386 149912 118514 149968
rect 118570 149912 118575 149968
rect 3325 149910 118575 149912
rect 3325 149907 3391 149910
rect 118509 149907 118575 149910
rect 0 148474 800 148504
rect 3049 148474 3115 148477
rect 0 148472 3115 148474
rect 0 148416 3054 148472
rect 3110 148416 3115 148472
rect 0 148414 3115 148416
rect 0 148384 800 148414
rect 3049 148411 3115 148414
rect 521653 148202 521719 148205
rect 519892 148200 521719 148202
rect 519892 148144 521658 148200
rect 521714 148144 521719 148200
rect 519892 148142 521719 148144
rect 521653 148139 521719 148142
rect 117313 147522 117379 147525
rect 117313 147520 120060 147522
rect 117313 147464 117318 147520
rect 117374 147464 120060 147520
rect 117313 147462 120060 147464
rect 117313 147459 117379 147462
rect 117129 146162 117195 146165
rect 113804 146160 117195 146162
rect 113804 146104 117134 146160
rect 117190 146104 117195 146160
rect 113804 146102 117195 146104
rect 117129 146099 117195 146102
rect 117221 144802 117287 144805
rect 117221 144800 120090 144802
rect 117221 144744 117226 144800
rect 117282 144744 120090 144800
rect 117221 144742 120090 144744
rect 117221 144739 117287 144742
rect 120030 144704 120090 144742
rect 0 143850 800 143880
rect 3417 143850 3483 143853
rect 0 143848 3483 143850
rect 0 143792 3422 143848
rect 3478 143792 3483 143848
rect 0 143790 3483 143792
rect 0 143760 800 143790
rect 3417 143787 3483 143790
rect 116669 141674 116735 141677
rect 116669 141672 120060 141674
rect 116669 141616 116674 141672
rect 116730 141616 120060 141672
rect 116669 141614 120060 141616
rect 116669 141611 116735 141614
rect 521745 140858 521811 140861
rect 519892 140856 521811 140858
rect 519892 140800 521750 140856
rect 521806 140800 521811 140856
rect 519892 140798 521811 140800
rect 521745 140795 521811 140798
rect 0 139362 800 139392
rect 3233 139362 3299 139365
rect 0 139360 3299 139362
rect 0 139304 3238 139360
rect 3294 139304 3299 139360
rect 0 139302 3299 139304
rect 0 139272 800 139302
rect 3233 139299 3299 139302
rect 118049 138818 118115 138821
rect 118049 138816 120060 138818
rect 118049 138760 118054 138816
rect 118110 138760 120060 138816
rect 118049 138758 120060 138760
rect 118049 138755 118115 138758
rect 117681 136506 117747 136509
rect 117681 136504 120090 136506
rect 117681 136448 117686 136504
rect 117742 136448 120090 136504
rect 117681 136446 120090 136448
rect 117681 136443 117747 136446
rect 120030 136000 120090 136446
rect 0 134738 800 134768
rect 3325 134738 3391 134741
rect 116761 134738 116827 134741
rect 0 134736 3391 134738
rect 0 134680 3330 134736
rect 3386 134680 3391 134736
rect 0 134678 3391 134680
rect 113804 134736 116827 134738
rect 113804 134680 116766 134736
rect 116822 134680 116827 134736
rect 113804 134678 116827 134680
rect 0 134648 800 134678
rect 3325 134675 3391 134678
rect 116761 134675 116827 134678
rect 520733 133378 520799 133381
rect 519892 133376 520799 133378
rect 519892 133320 520738 133376
rect 520794 133320 520799 133376
rect 519892 133318 520799 133320
rect 520733 133315 520799 133318
rect 117589 132970 117655 132973
rect 117589 132968 120060 132970
rect 117589 132912 117594 132968
rect 117650 132912 120060 132968
rect 117589 132910 120060 132912
rect 117589 132907 117655 132910
rect 0 130114 800 130144
rect 4061 130114 4127 130117
rect 0 130112 4127 130114
rect 0 130056 4066 130112
rect 4122 130056 4127 130112
rect 0 130054 4127 130056
rect 0 130024 800 130054
rect 4061 130051 4127 130054
rect 117313 130114 117379 130117
rect 117313 130112 120060 130114
rect 117313 130056 117318 130112
rect 117374 130056 120060 130112
rect 117313 130054 120060 130056
rect 117313 130051 117379 130054
rect 118233 127938 118299 127941
rect 118233 127936 120090 127938
rect 118233 127880 118238 127936
rect 118294 127880 120090 127936
rect 118233 127878 120090 127880
rect 118233 127875 118299 127878
rect 120030 127296 120090 127878
rect 521745 126034 521811 126037
rect 519892 126032 521811 126034
rect 519892 125976 521750 126032
rect 521806 125976 521811 126032
rect 519892 125974 521811 125976
rect 521745 125971 521811 125974
rect 0 125626 800 125656
rect 3969 125626 4035 125629
rect 0 125624 4035 125626
rect 0 125568 3974 125624
rect 4030 125568 4035 125624
rect 0 125566 4035 125568
rect 0 125536 800 125566
rect 3969 125563 4035 125566
rect 117313 124266 117379 124269
rect 117313 124264 120060 124266
rect 117313 124208 117318 124264
rect 117374 124208 120060 124264
rect 117313 124206 120060 124208
rect 117313 124203 117379 124206
rect 116853 123314 116919 123317
rect 113804 123312 116919 123314
rect 113804 123256 116858 123312
rect 116914 123256 116919 123312
rect 113804 123254 116919 123256
rect 116853 123251 116919 123254
rect 118233 121410 118299 121413
rect 118233 121408 120060 121410
rect 118233 121352 118238 121408
rect 118294 121352 120060 121408
rect 118233 121350 120060 121352
rect 118233 121347 118299 121350
rect 0 121002 800 121032
rect 3877 121002 3943 121005
rect 0 121000 3943 121002
rect 0 120944 3882 121000
rect 3938 120944 3943 121000
rect 0 120942 3943 120944
rect 0 120912 800 120942
rect 3877 120939 3943 120942
rect 118325 118690 118391 118693
rect 521837 118690 521903 118693
rect 118325 118688 120090 118690
rect 118325 118632 118330 118688
rect 118386 118632 120090 118688
rect 118325 118630 120090 118632
rect 519892 118688 521903 118690
rect 519892 118632 521842 118688
rect 521898 118632 521903 118688
rect 519892 118630 521903 118632
rect 118325 118627 118391 118630
rect 120030 118592 120090 118630
rect 521837 118627 521903 118630
rect 0 116514 800 116544
rect 3785 116514 3851 116517
rect 0 116512 3851 116514
rect 0 116456 3790 116512
rect 3846 116456 3851 116512
rect 0 116454 3851 116456
rect 0 116424 800 116454
rect 3785 116451 3851 116454
rect 118417 115834 118483 115837
rect 118417 115832 120090 115834
rect 118417 115776 118422 115832
rect 118478 115776 120090 115832
rect 118417 115774 120090 115776
rect 118417 115771 118483 115774
rect 120030 115600 120090 115774
rect 118417 112706 118483 112709
rect 118417 112704 120060 112706
rect 118417 112648 118422 112704
rect 118478 112648 120060 112704
rect 118417 112646 120060 112648
rect 118417 112643 118483 112646
rect 116945 112026 117011 112029
rect 113804 112024 117011 112026
rect 113804 111968 116950 112024
rect 117006 111968 117011 112024
rect 113804 111966 117011 111968
rect 116945 111963 117011 111966
rect 0 111890 800 111920
rect 3693 111890 3759 111893
rect 0 111888 3759 111890
rect 0 111832 3698 111888
rect 3754 111832 3759 111888
rect 0 111830 3759 111832
rect 0 111800 800 111830
rect 3693 111827 3759 111830
rect 521837 111210 521903 111213
rect 519892 111208 521903 111210
rect 519892 111152 521842 111208
rect 521898 111152 521903 111208
rect 519892 111150 521903 111152
rect 521837 111147 521903 111150
rect 116945 109850 117011 109853
rect 116945 109848 120060 109850
rect 116945 109792 116950 109848
rect 117006 109792 120060 109848
rect 116945 109790 120060 109792
rect 116945 109787 117011 109790
rect 0 107266 800 107296
rect 3601 107266 3667 107269
rect 0 107264 3667 107266
rect 0 107208 3606 107264
rect 3662 107208 3667 107264
rect 0 107206 3667 107208
rect 0 107176 800 107206
rect 3601 107203 3667 107206
rect 118693 106858 118759 106861
rect 118693 106856 120060 106858
rect 118693 106800 118698 106856
rect 118754 106800 120060 106856
rect 118693 106798 120060 106800
rect 118693 106795 118759 106798
rect 117497 104682 117563 104685
rect 117497 104680 120090 104682
rect 117497 104624 117502 104680
rect 117558 104624 120090 104680
rect 117497 104622 120090 104624
rect 117497 104619 117563 104622
rect 120030 104040 120090 104622
rect 521929 103866 521995 103869
rect 519892 103864 521995 103866
rect 519892 103808 521934 103864
rect 521990 103808 521995 103864
rect 519892 103806 521995 103808
rect 521929 103803 521995 103806
rect 0 102778 800 102808
rect 3509 102778 3575 102781
rect 0 102776 3575 102778
rect 0 102720 3514 102776
rect 3570 102720 3575 102776
rect 0 102718 3575 102720
rect 0 102688 800 102718
rect 3509 102715 3575 102718
rect 117865 101826 117931 101829
rect 117865 101824 120090 101826
rect 117865 101768 117870 101824
rect 117926 101768 120090 101824
rect 117865 101766 120090 101768
rect 117865 101763 117931 101766
rect 120030 101184 120090 101766
rect 116301 100602 116367 100605
rect 113804 100600 116367 100602
rect 113804 100544 116306 100600
rect 116362 100544 116367 100600
rect 113804 100542 116367 100544
rect 116301 100539 116367 100542
rect 117037 98834 117103 98837
rect 117037 98832 120090 98834
rect 117037 98776 117042 98832
rect 117098 98776 120090 98832
rect 117037 98774 120090 98776
rect 117037 98771 117103 98774
rect 120030 98192 120090 98774
rect 0 98154 800 98184
rect 3417 98154 3483 98157
rect 0 98152 3483 98154
rect 0 98096 3422 98152
rect 3478 98096 3483 98152
rect 0 98094 3483 98096
rect 0 98064 800 98094
rect 3417 98091 3483 98094
rect 522021 96386 522087 96389
rect 519892 96384 522087 96386
rect 519892 96328 522026 96384
rect 522082 96328 522087 96384
rect 519892 96326 522087 96328
rect 522021 96323 522087 96326
rect 117497 95978 117563 95981
rect 117497 95976 120090 95978
rect 117497 95920 117502 95976
rect 117558 95920 120090 95976
rect 117497 95918 120090 95920
rect 117497 95915 117563 95918
rect 120030 95336 120090 95918
rect 0 93666 800 93696
rect 3693 93666 3759 93669
rect 0 93664 3759 93666
rect 0 93608 3698 93664
rect 3754 93608 3759 93664
rect 0 93606 3759 93608
rect 0 93576 800 93606
rect 3693 93603 3759 93606
rect 118601 92442 118667 92445
rect 118601 92440 120060 92442
rect 118601 92384 118606 92440
rect 118662 92384 120060 92440
rect 118601 92382 120060 92384
rect 118601 92379 118667 92382
rect 118509 89722 118575 89725
rect 118509 89720 120090 89722
rect 118509 89664 118514 89720
rect 118570 89664 120090 89720
rect 118509 89662 120090 89664
rect 118509 89659 118575 89662
rect 120030 89488 120090 89662
rect 116894 89178 116900 89180
rect 113804 89118 116900 89178
rect 116894 89116 116900 89118
rect 116964 89116 116970 89180
rect 0 89042 800 89072
rect 3785 89042 3851 89045
rect 522113 89042 522179 89045
rect 0 89040 3851 89042
rect 0 88984 3790 89040
rect 3846 88984 3851 89040
rect 0 88982 3851 88984
rect 519892 89040 522179 89042
rect 519892 88984 522118 89040
rect 522174 88984 522179 89040
rect 519892 88982 522179 88984
rect 0 88952 800 88982
rect 3785 88979 3851 88982
rect 522113 88979 522179 88982
rect 117313 86866 117379 86869
rect 117313 86864 120090 86866
rect 117313 86808 117318 86864
rect 117374 86808 120090 86864
rect 117313 86806 120090 86808
rect 117313 86803 117379 86806
rect 120030 86632 120090 86806
rect 0 84418 800 84448
rect 3417 84418 3483 84421
rect 0 84416 3483 84418
rect 0 84360 3422 84416
rect 3478 84360 3483 84416
rect 0 84358 3483 84360
rect 0 84328 800 84358
rect 3417 84355 3483 84358
rect 117313 83874 117379 83877
rect 117313 83872 120090 83874
rect 117313 83816 117318 83872
rect 117374 83816 120090 83872
rect 117313 83814 120090 83816
rect 117313 83811 117379 83814
rect 120030 83776 120090 83814
rect 522205 81698 522271 81701
rect 519892 81696 522271 81698
rect 519892 81640 522210 81696
rect 522266 81640 522271 81696
rect 519892 81638 522271 81640
rect 522205 81635 522271 81638
rect 117681 81426 117747 81429
rect 117681 81424 120090 81426
rect 117681 81368 117686 81424
rect 117742 81368 120090 81424
rect 117681 81366 120090 81368
rect 117681 81363 117747 81366
rect 120030 80784 120090 81366
rect 0 79930 800 79960
rect 4061 79930 4127 79933
rect 0 79928 4127 79930
rect 0 79872 4066 79928
rect 4122 79872 4127 79928
rect 0 79870 4127 79872
rect 0 79840 800 79870
rect 4061 79867 4127 79870
rect 117681 78570 117747 78573
rect 117681 78568 120090 78570
rect 117681 78512 117686 78568
rect 117742 78512 120090 78568
rect 117681 78510 120090 78512
rect 117681 78507 117747 78510
rect 120030 77928 120090 78510
rect 116526 77890 116532 77892
rect 113804 77830 116532 77890
rect 116526 77828 116532 77830
rect 116596 77828 116602 77892
rect 118601 75714 118667 75717
rect 118601 75712 120090 75714
rect 118601 75656 118606 75712
rect 118662 75656 120090 75712
rect 118601 75654 120090 75656
rect 118601 75651 118667 75654
rect 0 75306 800 75336
rect 3969 75306 4035 75309
rect 0 75304 4035 75306
rect 0 75248 3974 75304
rect 4030 75248 4035 75304
rect 0 75246 4035 75248
rect 0 75216 800 75246
rect 3969 75243 4035 75246
rect 120030 75072 120090 75654
rect 522297 74218 522363 74221
rect 519892 74216 522363 74218
rect 519892 74160 522302 74216
rect 522358 74160 522363 74216
rect 519892 74158 522363 74160
rect 522297 74155 522363 74158
rect 117313 72722 117379 72725
rect 117313 72720 120090 72722
rect 117313 72664 117318 72720
rect 117374 72664 120090 72720
rect 117313 72662 120090 72664
rect 117313 72659 117379 72662
rect 120030 72080 120090 72662
rect 0 70818 800 70848
rect 3509 70818 3575 70821
rect 0 70816 3575 70818
rect 0 70760 3514 70816
rect 3570 70760 3575 70816
rect 0 70758 3575 70760
rect 0 70728 800 70758
rect 3509 70755 3575 70758
rect 117865 69866 117931 69869
rect 117865 69864 120090 69866
rect 117865 69808 117870 69864
rect 117926 69808 120090 69864
rect 117865 69806 120090 69808
rect 117865 69803 117931 69806
rect 120030 69224 120090 69806
rect 117313 67010 117379 67013
rect 117313 67008 120090 67010
rect 117313 66952 117318 67008
rect 117374 66952 120090 67008
rect 117313 66950 120090 66952
rect 117313 66947 117379 66950
rect 116301 66466 116367 66469
rect 113804 66464 116367 66466
rect 113804 66408 116306 66464
rect 116362 66408 116367 66464
rect 113804 66406 116367 66408
rect 116301 66403 116367 66406
rect 120030 66368 120090 66950
rect 521694 66874 521700 66876
rect 519892 66814 521700 66874
rect 521694 66812 521700 66814
rect 521764 66812 521770 66876
rect 0 66194 800 66224
rect 3601 66194 3667 66197
rect 0 66192 3667 66194
rect 0 66136 3606 66192
rect 3662 66136 3667 66192
rect 0 66134 3667 66136
rect 0 66104 800 66134
rect 3601 66131 3667 66134
rect 117865 63338 117931 63341
rect 117865 63336 120060 63338
rect 117865 63280 117870 63336
rect 117926 63280 120060 63336
rect 117865 63278 120060 63280
rect 117865 63275 117931 63278
rect 0 61570 800 61600
rect 3877 61570 3943 61573
rect 0 61568 3943 61570
rect 0 61512 3882 61568
rect 3938 61512 3943 61568
rect 0 61510 3943 61512
rect 0 61480 800 61510
rect 3877 61507 3943 61510
rect 118601 60482 118667 60485
rect 118601 60480 120060 60482
rect 118601 60424 118606 60480
rect 118662 60424 120060 60480
rect 118601 60422 120060 60424
rect 118601 60419 118667 60422
rect 520222 59530 520228 59532
rect 519862 59470 520228 59530
rect 519862 59364 519922 59470
rect 520222 59468 520228 59470
rect 520292 59468 520298 59532
rect 117313 57626 117379 57629
rect 117313 57624 120060 57626
rect 117313 57568 117318 57624
rect 117374 57568 120060 57624
rect 117313 57566 120060 57568
rect 117313 57563 117379 57566
rect 0 57082 800 57112
rect 3325 57082 3391 57085
rect 0 57080 3391 57082
rect 0 57024 3330 57080
rect 3386 57024 3391 57080
rect 0 57022 3391 57024
rect 0 56992 800 57022
rect 3325 57019 3391 57022
rect 116526 55042 116532 55044
rect 113804 54982 116532 55042
rect 116526 54980 116532 54982
rect 116596 54980 116602 55044
rect 118509 54634 118575 54637
rect 118509 54632 120060 54634
rect 118509 54576 118514 54632
rect 118570 54576 120060 54632
rect 118509 54574 120060 54576
rect 118509 54571 118575 54574
rect 0 52458 800 52488
rect 3233 52458 3299 52461
rect 0 52456 3299 52458
rect 0 52400 3238 52456
rect 3294 52400 3299 52456
rect 0 52398 3299 52400
rect 0 52368 800 52398
rect 3233 52395 3299 52398
rect 522573 52050 522639 52053
rect 519892 52048 522639 52050
rect 519892 51992 522578 52048
rect 522634 51992 522639 52048
rect 519892 51990 522639 51992
rect 522573 51987 522639 51990
rect 117313 51778 117379 51781
rect 117313 51776 120060 51778
rect 117313 51720 117318 51776
rect 117374 51720 120060 51776
rect 117313 51718 120060 51720
rect 117313 51715 117379 51718
rect 117405 48922 117471 48925
rect 117405 48920 120060 48922
rect 117405 48864 117410 48920
rect 117466 48864 120060 48920
rect 117405 48862 120060 48864
rect 117405 48859 117471 48862
rect 0 47970 800 48000
rect 3141 47970 3207 47973
rect 0 47968 3207 47970
rect 0 47912 3146 47968
rect 3202 47912 3207 47968
rect 0 47910 3207 47912
rect 0 47880 800 47910
rect 3141 47907 3207 47910
rect 117313 45930 117379 45933
rect 117313 45928 120060 45930
rect 117313 45872 117318 45928
rect 117374 45872 120060 45928
rect 117313 45870 120060 45872
rect 117313 45867 117379 45870
rect 521694 44706 521700 44708
rect 519892 44646 521700 44706
rect 521694 44644 521700 44646
rect 521764 44644 521770 44708
rect 116894 43754 116900 43756
rect 113804 43694 116900 43754
rect 116894 43692 116900 43694
rect 116964 43692 116970 43756
rect 0 43346 800 43376
rect 3049 43346 3115 43349
rect 0 43344 3115 43346
rect 0 43288 3054 43344
rect 3110 43288 3115 43344
rect 0 43286 3115 43288
rect 0 43256 800 43286
rect 3049 43283 3115 43286
rect 117313 43074 117379 43077
rect 117313 43072 120060 43074
rect 117313 43016 117318 43072
rect 117374 43016 120060 43072
rect 117313 43014 120060 43016
rect 117313 43011 117379 43014
rect 117865 40218 117931 40221
rect 117865 40216 120060 40218
rect 117865 40160 117870 40216
rect 117926 40160 120060 40216
rect 117865 40158 120060 40160
rect 117865 40155 117931 40158
rect 0 38722 800 38752
rect 2957 38722 3023 38725
rect 0 38720 3023 38722
rect 0 38664 2962 38720
rect 3018 38664 3023 38720
rect 0 38662 3023 38664
rect 0 38632 800 38662
rect 2957 38659 3023 38662
rect 117221 37226 117287 37229
rect 520825 37226 520891 37229
rect 117221 37224 120060 37226
rect 117221 37168 117226 37224
rect 117282 37168 120060 37224
rect 117221 37166 120060 37168
rect 519892 37224 520891 37226
rect 519892 37168 520830 37224
rect 520886 37168 520891 37224
rect 519892 37166 520891 37168
rect 117221 37163 117287 37166
rect 520825 37163 520891 37166
rect 117129 34370 117195 34373
rect 117129 34368 120060 34370
rect 117129 34312 117134 34368
rect 117190 34312 120060 34368
rect 117129 34310 120060 34312
rect 117129 34307 117195 34310
rect 0 34234 800 34264
rect 2865 34234 2931 34237
rect 0 34232 2931 34234
rect 0 34176 2870 34232
rect 2926 34176 2931 34232
rect 0 34174 2931 34176
rect 0 34144 800 34174
rect 2865 34171 2931 34174
rect 117037 32330 117103 32333
rect 113804 32328 117103 32330
rect 113804 32272 117042 32328
rect 117098 32272 117103 32328
rect 113804 32270 117103 32272
rect 117037 32267 117103 32270
rect 117313 31514 117379 31517
rect 117313 31512 120060 31514
rect 117313 31456 117318 31512
rect 117374 31456 120060 31512
rect 117313 31454 120060 31456
rect 117313 31451 117379 31454
rect 522062 29882 522068 29884
rect 519892 29822 522068 29882
rect 522062 29820 522068 29822
rect 522132 29820 522138 29884
rect 0 29610 800 29640
rect 3693 29610 3759 29613
rect 0 29608 3759 29610
rect 0 29552 3698 29608
rect 3754 29552 3759 29608
rect 0 29550 3759 29552
rect 0 29520 800 29550
rect 3693 29547 3759 29550
rect 118509 28522 118575 28525
rect 118509 28520 120060 28522
rect 118509 28464 118514 28520
rect 118570 28464 120060 28520
rect 118509 28462 120060 28464
rect 118509 28459 118575 28462
rect 118601 25666 118667 25669
rect 118601 25664 120060 25666
rect 118601 25608 118606 25664
rect 118662 25608 120060 25664
rect 118601 25606 120060 25608
rect 118601 25603 118667 25606
rect 0 25122 800 25152
rect 3785 25122 3851 25125
rect 0 25120 3851 25122
rect 0 25064 3790 25120
rect 3846 25064 3851 25120
rect 0 25062 3851 25064
rect 0 25032 800 25062
rect 3785 25059 3851 25062
rect 117865 22810 117931 22813
rect 117865 22808 120060 22810
rect 117865 22752 117870 22808
rect 117926 22752 120060 22808
rect 117865 22750 120060 22752
rect 117865 22747 117931 22750
rect 522389 22402 522455 22405
rect 519892 22400 522455 22402
rect 519892 22344 522394 22400
rect 522450 22344 522455 22400
rect 519892 22342 522455 22344
rect 522389 22339 522455 22342
rect 116485 20906 116551 20909
rect 113804 20904 116551 20906
rect 113804 20848 116490 20904
rect 116546 20848 116551 20904
rect 113804 20846 116551 20848
rect 116485 20843 116551 20846
rect 0 20498 800 20528
rect 4061 20498 4127 20501
rect 0 20496 4127 20498
rect 0 20440 4066 20496
rect 4122 20440 4127 20496
rect 0 20438 4127 20440
rect 0 20408 800 20438
rect 4061 20435 4127 20438
rect 117773 19818 117839 19821
rect 117773 19816 120060 19818
rect 117773 19760 117778 19816
rect 117834 19760 120060 19816
rect 117773 19758 120060 19760
rect 117773 19755 117839 19758
rect 117497 16962 117563 16965
rect 117497 16960 120060 16962
rect 117497 16904 117502 16960
rect 117558 16904 120060 16960
rect 117497 16902 120060 16904
rect 117497 16899 117563 16902
rect 0 15874 800 15904
rect 3417 15874 3483 15877
rect 0 15872 3483 15874
rect 0 15816 3422 15872
rect 3478 15816 3483 15872
rect 0 15814 3483 15816
rect 0 15784 800 15814
rect 3417 15811 3483 15814
rect 520917 15058 520983 15061
rect 519892 15056 520983 15058
rect 519892 15000 520922 15056
rect 520978 15000 520983 15056
rect 519892 14998 520983 15000
rect 520917 14995 520983 14998
rect 117313 14106 117379 14109
rect 117313 14104 120060 14106
rect 117313 14048 117318 14104
rect 117374 14048 120060 14104
rect 117313 14046 120060 14048
rect 117313 14043 117379 14046
rect 0 11386 800 11416
rect 3969 11386 4035 11389
rect 0 11384 4035 11386
rect 0 11328 3974 11384
rect 4030 11328 4035 11384
rect 0 11326 4035 11328
rect 0 11296 800 11326
rect 3969 11323 4035 11326
rect 117313 11114 117379 11117
rect 117313 11112 120060 11114
rect 117313 11056 117318 11112
rect 117374 11056 120060 11112
rect 117313 11054 120060 11056
rect 117313 11051 117379 11054
rect 116945 9618 117011 9621
rect 113804 9616 117011 9618
rect 113804 9560 116950 9616
rect 117006 9560 117011 9616
rect 113804 9558 117011 9560
rect 116945 9555 117011 9558
rect 117313 8258 117379 8261
rect 117313 8256 120060 8258
rect 117313 8200 117318 8256
rect 117374 8200 120060 8256
rect 117313 8198 120060 8200
rect 117313 8195 117379 8198
rect 522941 7714 523007 7717
rect 519892 7712 523007 7714
rect 519892 7656 522946 7712
rect 523002 7656 523007 7712
rect 519892 7654 523007 7656
rect 522941 7651 523007 7654
rect 0 6762 800 6792
rect 3233 6762 3299 6765
rect 0 6760 3299 6762
rect 0 6704 3238 6760
rect 3294 6704 3299 6760
rect 0 6702 3299 6704
rect 0 6672 800 6702
rect 3233 6699 3299 6702
rect 4981 6082 5047 6085
rect 115013 6082 115079 6085
rect 4981 6080 115079 6082
rect 4981 6024 4986 6080
rect 5042 6024 115018 6080
rect 115074 6024 115079 6080
rect 4981 6022 115079 6024
rect 4981 6019 5047 6022
rect 115013 6019 115079 6022
rect 5441 5946 5507 5949
rect 112529 5946 112595 5949
rect 5441 5944 112595 5946
rect 5441 5888 5446 5944
rect 5502 5888 112534 5944
rect 112590 5888 112595 5944
rect 5441 5886 112595 5888
rect 5441 5883 5507 5886
rect 112529 5883 112595 5886
rect 77250 5750 82186 5810
rect 77250 5538 77310 5750
rect 75870 5478 77310 5538
rect 75870 5130 75930 5478
rect 72374 5070 75930 5130
rect 35850 4798 60750 4858
rect 35850 4589 35910 4798
rect 35801 4584 35910 4589
rect 35801 4528 35806 4584
rect 35862 4528 35910 4584
rect 35801 4526 35910 4528
rect 35801 4523 35867 4526
rect 60690 4450 60750 4798
rect 72374 4589 72434 5070
rect 77250 4934 82002 4994
rect 65977 4586 66043 4589
rect 71957 4586 72023 4589
rect 65977 4584 72023 4586
rect 65977 4528 65982 4584
rect 66038 4528 71962 4584
rect 72018 4528 72023 4584
rect 65977 4526 72023 4528
rect 72374 4584 72483 4589
rect 72374 4528 72422 4584
rect 72478 4528 72483 4584
rect 72374 4526 72483 4528
rect 65977 4523 66043 4526
rect 71957 4523 72023 4526
rect 72417 4523 72483 4526
rect 74901 4586 74967 4589
rect 77250 4586 77310 4934
rect 74901 4584 77310 4586
rect 74901 4528 74906 4584
rect 74962 4528 77310 4584
rect 74901 4526 77310 4528
rect 81942 4589 82002 4934
rect 82126 4589 82186 5750
rect 91050 5750 98010 5810
rect 91050 5266 91110 5750
rect 97950 5674 98010 5750
rect 99330 5750 100770 5810
rect 99330 5674 99390 5750
rect 97950 5614 99390 5674
rect 97950 5478 99390 5538
rect 97950 5266 98010 5478
rect 85622 5206 91110 5266
rect 96570 5206 98010 5266
rect 85622 4722 85682 5206
rect 96570 5130 96630 5206
rect 82632 4662 85682 4722
rect 85806 5070 96630 5130
rect 99330 5130 99390 5478
rect 100710 5266 100770 5750
rect 117313 5402 117379 5405
rect 117313 5400 120060 5402
rect 117313 5344 117318 5400
rect 117374 5344 120060 5400
rect 117313 5342 120060 5344
rect 117313 5339 117379 5342
rect 521745 5266 521811 5269
rect 100710 5264 521811 5266
rect 100710 5208 521750 5264
rect 521806 5208 521811 5264
rect 100710 5206 521811 5208
rect 521745 5203 521811 5206
rect 520457 5130 520523 5133
rect 99330 5128 520523 5130
rect 99330 5072 520462 5128
rect 520518 5072 520523 5128
rect 99330 5070 520523 5072
rect 82632 4589 82692 4662
rect 81942 4584 82051 4589
rect 81942 4528 81990 4584
rect 82046 4528 82051 4584
rect 81942 4526 82051 4528
rect 82126 4584 82235 4589
rect 82126 4528 82174 4584
rect 82230 4528 82235 4584
rect 82126 4526 82235 4528
rect 74901 4523 74967 4526
rect 81985 4523 82051 4526
rect 82169 4523 82235 4526
rect 82629 4584 82695 4589
rect 82629 4528 82634 4584
rect 82690 4528 82695 4584
rect 82629 4523 82695 4528
rect 82813 4586 82879 4589
rect 85806 4586 85866 5070
rect 520457 5067 520523 5070
rect 521929 4994 521995 4997
rect 86910 4992 521995 4994
rect 86910 4936 521934 4992
rect 521990 4936 521995 4992
rect 86910 4934 521995 4936
rect 82813 4584 85866 4586
rect 82813 4528 82818 4584
rect 82874 4528 85866 4584
rect 82813 4526 85866 4528
rect 86401 4586 86467 4589
rect 86910 4586 86970 4934
rect 521929 4931 521995 4934
rect 523033 4858 523099 4861
rect 86401 4584 86970 4586
rect 86401 4528 86406 4584
rect 86462 4528 86970 4584
rect 86401 4526 86970 4528
rect 89670 4856 523099 4858
rect 89670 4800 523038 4856
rect 523094 4800 523099 4856
rect 89670 4798 523099 4800
rect 82813 4523 82879 4526
rect 86401 4523 86467 4526
rect 89670 4450 89730 4798
rect 523033 4795 523099 4798
rect 521653 4722 521719 4725
rect 103470 4720 521719 4722
rect 103470 4664 521658 4720
rect 521714 4664 521719 4720
rect 103470 4662 521719 4664
rect 102685 4586 102751 4589
rect 103470 4586 103530 4662
rect 521653 4659 521719 4662
rect 102685 4584 103530 4586
rect 102685 4528 102690 4584
rect 102746 4528 103530 4584
rect 102685 4526 103530 4528
rect 102685 4523 102751 4526
rect 60690 4390 67650 4450
rect 67590 4178 67650 4390
rect 77250 4390 89730 4450
rect 77250 4178 77310 4390
rect 67590 4118 77310 4178
rect 115197 3090 115263 3093
rect 475009 3090 475075 3093
rect 115197 3088 475075 3090
rect 115197 3032 115202 3088
rect 115258 3032 475014 3088
rect 475070 3032 475075 3088
rect 115197 3030 475075 3032
rect 115197 3027 115263 3030
rect 475009 3027 475075 3030
rect 113909 2954 113975 2957
rect 518065 2954 518131 2957
rect 113909 2952 518131 2954
rect 113909 2896 113914 2952
rect 113970 2896 518070 2952
rect 518126 2896 518131 2952
rect 113909 2894 518131 2896
rect 113909 2891 113975 2894
rect 518065 2891 518131 2894
rect 49325 2818 49391 2821
rect 520273 2818 520339 2821
rect 49325 2816 520339 2818
rect 49325 2760 49330 2816
rect 49386 2760 520278 2816
rect 520334 2760 520339 2816
rect 49325 2758 520339 2760
rect 49325 2755 49391 2758
rect 520273 2755 520339 2758
rect 119613 2682 119679 2685
rect 484393 2682 484459 2685
rect 119613 2680 484459 2682
rect 119613 2624 119618 2680
rect 119674 2624 484398 2680
rect 484454 2624 484459 2680
rect 119613 2622 484459 2624
rect 119613 2619 119679 2622
rect 484393 2619 484459 2622
rect 119981 2546 120047 2549
rect 481173 2546 481239 2549
rect 119981 2544 481239 2546
rect 119981 2488 119986 2544
rect 120042 2488 481178 2544
rect 481234 2488 481239 2544
rect 119981 2486 481239 2488
rect 119981 2483 120047 2486
rect 481173 2483 481239 2486
rect 115473 2410 115539 2413
rect 471973 2410 472039 2413
rect 115473 2408 472039 2410
rect 115473 2352 115478 2408
rect 115534 2352 471978 2408
rect 472034 2352 472039 2408
rect 115473 2350 472039 2352
rect 115473 2347 115539 2350
rect 471973 2347 472039 2350
rect 0 2274 800 2304
rect 2957 2274 3023 2277
rect 0 2272 3023 2274
rect 0 2216 2962 2272
rect 3018 2216 3023 2272
rect 0 2214 3023 2216
rect 0 2184 800 2214
rect 2957 2211 3023 2214
rect 119429 2274 119495 2277
rect 465717 2274 465783 2277
rect 119429 2272 465783 2274
rect 119429 2216 119434 2272
rect 119490 2216 465722 2272
rect 465778 2216 465783 2272
rect 119429 2214 465783 2216
rect 119429 2211 119495 2214
rect 465717 2211 465783 2214
rect 118141 2138 118207 2141
rect 456793 2138 456859 2141
rect 118141 2136 456859 2138
rect 118141 2080 118146 2136
rect 118202 2080 456798 2136
rect 456854 2080 456859 2136
rect 118141 2078 456859 2080
rect 118141 2075 118207 2078
rect 456793 2075 456859 2078
rect 115657 2002 115723 2005
rect 450353 2002 450419 2005
rect 115657 2000 450419 2002
rect 115657 1944 115662 2000
rect 115718 1944 450358 2000
rect 450414 1944 450419 2000
rect 115657 1942 450419 1944
rect 115657 1939 115723 1942
rect 450353 1939 450419 1942
rect 118325 1866 118391 1869
rect 447317 1866 447383 1869
rect 118325 1864 447383 1866
rect 118325 1808 118330 1864
rect 118386 1808 447322 1864
rect 447378 1808 447383 1864
rect 118325 1806 447383 1808
rect 118325 1803 118391 1806
rect 447317 1803 447383 1806
<< via3 >>
rect 116900 89116 116964 89180
rect 116532 77828 116596 77892
rect 521700 66812 521764 66876
rect 520228 59468 520292 59532
rect 116532 54980 116596 55044
rect 521700 44644 521764 44708
rect 116900 43692 116964 43756
rect 522068 29820 522132 29884
<< metal4 >>
rect 4208 154000 4528 157760
rect 9208 154000 9528 157760
rect 14208 154000 14528 157760
rect 19208 154000 19528 157760
rect 24208 154000 24528 157760
rect 29208 154000 29528 157760
rect 34208 154000 34528 157760
rect 39208 154000 39528 157760
rect 44208 154000 44528 157760
rect 49208 154000 49528 157760
rect 54208 154000 54528 157760
rect 59208 154000 59528 157760
rect 64208 154000 64528 157760
rect 69208 154000 69528 157760
rect 74208 154000 74528 157760
rect 79208 154000 79528 157760
rect 84208 154000 84528 157760
rect 89208 154000 89528 157760
rect 94208 154000 94528 157760
rect 99208 154000 99528 157760
rect 104208 154000 104528 157760
rect 109208 154000 109528 157760
rect 114208 154000 114528 157760
rect 119208 154000 119528 157760
rect 124208 154000 124528 157760
rect 129208 154000 129528 157760
rect 134208 154000 134528 157760
rect 139208 154000 139528 157760
rect 144208 154000 144528 157760
rect 149208 154000 149528 157760
rect 154208 154000 154528 157760
rect 159208 154000 159528 157760
rect 164208 154000 164528 157760
rect 169208 154000 169528 157760
rect 174208 154000 174528 157760
rect 179208 154000 179528 157760
rect 184208 154000 184528 157760
rect 189208 154000 189528 157760
rect 194208 154000 194528 157760
rect 199208 154000 199528 157760
rect 204208 154000 204528 157760
rect 209208 154000 209528 157760
rect 214208 154000 214528 157760
rect 219208 154000 219528 157760
rect 224208 154000 224528 157760
rect 229208 154000 229528 157760
rect 234208 154000 234528 157760
rect 239208 154000 239528 157760
rect 244208 154000 244528 157760
rect 249208 154000 249528 157760
rect 254208 154000 254528 157760
rect 259208 154000 259528 157760
rect 264208 154000 264528 157760
rect 269208 154000 269528 157760
rect 274208 154000 274528 157760
rect 279208 154000 279528 157760
rect 284208 154000 284528 157760
rect 289208 154000 289528 157760
rect 294208 154000 294528 157760
rect 299208 154000 299528 157760
rect 304208 154000 304528 157760
rect 309208 154000 309528 157760
rect 314208 154000 314528 157760
rect 319208 154000 319528 157760
rect 324208 154000 324528 157760
rect 329208 154000 329528 157760
rect 334208 154000 334528 157760
rect 339208 154000 339528 157760
rect 344208 154000 344528 157760
rect 349208 154000 349528 157760
rect 354208 154000 354528 157760
rect 359208 154000 359528 157760
rect 364208 154000 364528 157760
rect 369208 154000 369528 157760
rect 374208 154000 374528 157760
rect 379208 154000 379528 157760
rect 384208 154000 384528 157760
rect 389208 154000 389528 157760
rect 394208 154000 394528 157760
rect 399208 154000 399528 157760
rect 404208 154000 404528 157760
rect 409208 154000 409528 157760
rect 414208 154000 414528 157760
rect 419208 154000 419528 157760
rect 424208 154000 424528 157760
rect 429208 154000 429528 157760
rect 434208 154000 434528 157760
rect 439208 154000 439528 157760
rect 444208 154000 444528 157760
rect 449208 154000 449528 157760
rect 454208 154000 454528 157760
rect 459208 154000 459528 157760
rect 464208 154000 464528 157760
rect 469208 154000 469528 157760
rect 474208 154000 474528 157760
rect 479208 154000 479528 157760
rect 484208 154000 484528 157760
rect 489208 154000 489528 157760
rect 494208 154000 494528 157760
rect 499208 154000 499528 157760
rect 504208 154000 504528 157760
rect 509208 154000 509528 157760
rect 514208 154000 514528 157760
rect 519208 154000 519528 157760
rect 524208 135624 524528 157760
rect 524208 135388 524250 135624
rect 524486 135388 524528 135624
rect 524208 109624 524528 135388
rect 524208 109388 524250 109624
rect 524486 109388 524528 109624
rect 116899 89180 116965 89181
rect 116899 89116 116900 89180
rect 116964 89116 116965 89180
rect 116899 89115 116965 89116
rect 116531 77892 116597 77893
rect 116531 77828 116532 77892
rect 116596 77828 116597 77892
rect 116531 77827 116597 77828
rect 116534 62338 116594 77827
rect 116902 73898 116962 89115
rect 524208 83624 524528 109388
rect 524208 83388 524250 83624
rect 524486 83388 524528 83624
rect 521702 66877 521762 75022
rect 521699 66876 521765 66877
rect 521699 66812 521700 66876
rect 521764 66812 521765 66876
rect 521699 66811 521765 66812
rect 512870 59618 512930 62102
rect 524208 57624 524528 83388
rect 524208 57388 524250 57624
rect 524486 57388 524528 57624
rect 116531 55044 116597 55045
rect 116531 54980 116532 55044
rect 116596 54980 116597 55044
rect 116531 54979 116597 54980
rect 116534 20858 116594 54979
rect 521699 44708 521765 44709
rect 521699 44644 521700 44708
rect 521764 44644 521765 44708
rect 521699 44643 521765 44644
rect 116899 43756 116965 43757
rect 116899 43692 116900 43756
rect 116964 43692 116965 43756
rect 116899 43691 116965 43692
rect 116902 22218 116962 43691
rect 512870 21538 512930 23342
rect 521702 21538 521762 44643
rect 524208 31624 524528 57388
rect 524208 31388 524250 31624
rect 524486 31388 524528 31624
rect 522067 29884 522133 29885
rect 522067 29820 522068 29884
rect 522132 29820 522133 29884
rect 522067 29819 522133 29820
rect 522070 23578 522130 29819
rect 524208 5624 524528 31388
rect 524208 5388 524250 5624
rect 524486 5388 524528 5624
rect 524208 2176 524528 5388
rect 529208 148624 529528 157760
rect 529208 148388 529250 148624
rect 529486 148388 529528 148624
rect 529208 122624 529528 148388
rect 529208 122388 529250 122624
rect 529486 122388 529528 122624
rect 529208 96624 529528 122388
rect 529208 96388 529250 96624
rect 529486 96388 529528 96624
rect 529208 70624 529528 96388
rect 529208 70388 529250 70624
rect 529486 70388 529528 70624
rect 529208 44624 529528 70388
rect 529208 44388 529250 44624
rect 529486 44388 529528 44624
rect 529208 18624 529528 44388
rect 529208 18388 529250 18624
rect 529486 18388 529528 18624
rect 529208 2176 529528 18388
rect 534208 135624 534528 157760
rect 534208 135388 534250 135624
rect 534486 135388 534528 135624
rect 534208 109624 534528 135388
rect 534208 109388 534250 109624
rect 534486 109388 534528 109624
rect 534208 83624 534528 109388
rect 534208 83388 534250 83624
rect 534486 83388 534528 83624
rect 534208 57624 534528 83388
rect 534208 57388 534250 57624
rect 534486 57388 534528 57624
rect 534208 31624 534528 57388
rect 534208 31388 534250 31624
rect 534486 31388 534528 31624
rect 534208 5624 534528 31388
rect 534208 5388 534250 5624
rect 534486 5388 534528 5624
rect 534208 2176 534528 5388
rect 539208 148624 539528 157760
rect 539208 148388 539250 148624
rect 539486 148388 539528 148624
rect 539208 122624 539528 148388
rect 539208 122388 539250 122624
rect 539486 122388 539528 122624
rect 539208 96624 539528 122388
rect 539208 96388 539250 96624
rect 539486 96388 539528 96624
rect 539208 70624 539528 96388
rect 539208 70388 539250 70624
rect 539486 70388 539528 70624
rect 539208 44624 539528 70388
rect 539208 44388 539250 44624
rect 539486 44388 539528 44624
rect 539208 18624 539528 44388
rect 539208 18388 539250 18624
rect 539486 18388 539528 18624
rect 539208 2176 539528 18388
rect 544208 135624 544528 157760
rect 544208 135388 544250 135624
rect 544486 135388 544528 135624
rect 544208 109624 544528 135388
rect 544208 109388 544250 109624
rect 544486 109388 544528 109624
rect 544208 83624 544528 109388
rect 544208 83388 544250 83624
rect 544486 83388 544528 83624
rect 544208 57624 544528 83388
rect 544208 57388 544250 57624
rect 544486 57388 544528 57624
rect 544208 31624 544528 57388
rect 544208 31388 544250 31624
rect 544486 31388 544528 31624
rect 544208 5624 544528 31388
rect 544208 5388 544250 5624
rect 544486 5388 544528 5624
rect 544208 2176 544528 5388
rect 549208 148624 549528 157760
rect 549208 148388 549250 148624
rect 549486 148388 549528 148624
rect 549208 122624 549528 148388
rect 549208 122388 549250 122624
rect 549486 122388 549528 122624
rect 549208 96624 549528 122388
rect 549208 96388 549250 96624
rect 549486 96388 549528 96624
rect 549208 70624 549528 96388
rect 549208 70388 549250 70624
rect 549486 70388 549528 70624
rect 549208 44624 549528 70388
rect 549208 44388 549250 44624
rect 549486 44388 549528 44624
rect 549208 18624 549528 44388
rect 549208 18388 549250 18624
rect 549486 18388 549528 18624
rect 549208 2176 549528 18388
rect 554208 135624 554528 157760
rect 554208 135388 554250 135624
rect 554486 135388 554528 135624
rect 554208 109624 554528 135388
rect 554208 109388 554250 109624
rect 554486 109388 554528 109624
rect 554208 83624 554528 109388
rect 554208 83388 554250 83624
rect 554486 83388 554528 83624
rect 554208 57624 554528 83388
rect 554208 57388 554250 57624
rect 554486 57388 554528 57624
rect 554208 31624 554528 57388
rect 554208 31388 554250 31624
rect 554486 31388 554528 31624
rect 554208 5624 554528 31388
rect 554208 5388 554250 5624
rect 554486 5388 554528 5624
rect 554208 2176 554528 5388
rect 559208 148624 559528 157760
rect 559208 148388 559250 148624
rect 559486 148388 559528 148624
rect 559208 122624 559528 148388
rect 559208 122388 559250 122624
rect 559486 122388 559528 122624
rect 559208 96624 559528 122388
rect 559208 96388 559250 96624
rect 559486 96388 559528 96624
rect 559208 70624 559528 96388
rect 559208 70388 559250 70624
rect 559486 70388 559528 70624
rect 559208 44624 559528 70388
rect 559208 44388 559250 44624
rect 559486 44388 559528 44624
rect 559208 18624 559528 44388
rect 559208 18388 559250 18624
rect 559486 18388 559528 18624
rect 559208 2176 559528 18388
rect 564208 135624 564528 157760
rect 564208 135388 564250 135624
rect 564486 135388 564528 135624
rect 564208 109624 564528 135388
rect 564208 109388 564250 109624
rect 564486 109388 564528 109624
rect 564208 83624 564528 109388
rect 564208 83388 564250 83624
rect 564486 83388 564528 83624
rect 564208 57624 564528 83388
rect 564208 57388 564250 57624
rect 564486 57388 564528 57624
rect 564208 31624 564528 57388
rect 564208 31388 564250 31624
rect 564486 31388 564528 31624
rect 564208 5624 564528 31388
rect 564208 5388 564250 5624
rect 564486 5388 564528 5624
rect 564208 2176 564528 5388
rect 569208 148624 569528 157760
rect 569208 148388 569250 148624
rect 569486 148388 569528 148624
rect 569208 122624 569528 148388
rect 569208 122388 569250 122624
rect 569486 122388 569528 122624
rect 569208 96624 569528 122388
rect 569208 96388 569250 96624
rect 569486 96388 569528 96624
rect 569208 70624 569528 96388
rect 569208 70388 569250 70624
rect 569486 70388 569528 70624
rect 569208 44624 569528 70388
rect 569208 44388 569250 44624
rect 569486 44388 569528 44624
rect 569208 18624 569528 44388
rect 569208 18388 569250 18624
rect 569486 18388 569528 18624
rect 569208 2176 569528 18388
rect 574208 135624 574528 157760
rect 574208 135388 574250 135624
rect 574486 135388 574528 135624
rect 574208 109624 574528 135388
rect 574208 109388 574250 109624
rect 574486 109388 574528 109624
rect 574208 83624 574528 109388
rect 574208 83388 574250 83624
rect 574486 83388 574528 83624
rect 574208 57624 574528 83388
rect 574208 57388 574250 57624
rect 574486 57388 574528 57624
rect 574208 31624 574528 57388
rect 574208 31388 574250 31624
rect 574486 31388 574528 31624
rect 574208 5624 574528 31388
rect 574208 5388 574250 5624
rect 574486 5388 574528 5624
rect 574208 2176 574528 5388
<< via4 >>
rect 524250 135388 524486 135624
rect 524250 109388 524486 109624
rect 524250 83388 524486 83624
rect 521614 75022 521850 75258
rect 116814 73662 117050 73898
rect 116446 62102 116682 62338
rect 512782 62102 513018 62338
rect 512782 59382 513018 59618
rect 520142 59532 520378 59618
rect 520142 59468 520228 59532
rect 520228 59468 520292 59532
rect 520292 59468 520378 59532
rect 520142 59382 520378 59468
rect 524250 57388 524486 57624
rect 512782 23342 513018 23578
rect 116814 21982 117050 22218
rect 524250 31388 524486 31624
rect 521982 23342 522218 23578
rect 512782 21302 513018 21538
rect 521614 21302 521850 21538
rect 116446 20622 116682 20858
rect 524250 5388 524486 5624
rect 529250 148388 529486 148624
rect 529250 122388 529486 122624
rect 529250 96388 529486 96624
rect 529250 70388 529486 70624
rect 529250 44388 529486 44624
rect 529250 18388 529486 18624
rect 534250 135388 534486 135624
rect 534250 109388 534486 109624
rect 534250 83388 534486 83624
rect 534250 57388 534486 57624
rect 534250 31388 534486 31624
rect 534250 5388 534486 5624
rect 539250 148388 539486 148624
rect 539250 122388 539486 122624
rect 539250 96388 539486 96624
rect 539250 70388 539486 70624
rect 539250 44388 539486 44624
rect 539250 18388 539486 18624
rect 544250 135388 544486 135624
rect 544250 109388 544486 109624
rect 544250 83388 544486 83624
rect 544250 57388 544486 57624
rect 544250 31388 544486 31624
rect 544250 5388 544486 5624
rect 549250 148388 549486 148624
rect 549250 122388 549486 122624
rect 549250 96388 549486 96624
rect 549250 70388 549486 70624
rect 549250 44388 549486 44624
rect 549250 18388 549486 18624
rect 554250 135388 554486 135624
rect 554250 109388 554486 109624
rect 554250 83388 554486 83624
rect 554250 57388 554486 57624
rect 554250 31388 554486 31624
rect 554250 5388 554486 5624
rect 559250 148388 559486 148624
rect 559250 122388 559486 122624
rect 559250 96388 559486 96624
rect 559250 70388 559486 70624
rect 559250 44388 559486 44624
rect 559250 18388 559486 18624
rect 564250 135388 564486 135624
rect 564250 109388 564486 109624
rect 564250 83388 564486 83624
rect 564250 57388 564486 57624
rect 564250 31388 564486 31624
rect 564250 5388 564486 5624
rect 569250 148388 569486 148624
rect 569250 122388 569486 122624
rect 569250 96388 569486 96624
rect 569250 70388 569486 70624
rect 569250 44388 569486 44624
rect 569250 18388 569486 18624
rect 574250 135388 574486 135624
rect 574250 109388 574486 109624
rect 574250 83388 574486 83624
rect 574250 57388 574486 57624
rect 574250 31388 574486 31624
rect 574250 5388 574486 5624
<< metal5 >>
rect 1104 148346 2000 148666
rect 116000 148346 118000 148666
rect 522000 148624 578864 148666
rect 522000 148388 529250 148624
rect 529486 148388 539250 148624
rect 539486 148388 549250 148624
rect 549486 148388 559250 148624
rect 559486 148388 569250 148624
rect 569486 148388 578864 148624
rect 522000 148346 578864 148388
rect 1104 135346 2000 135666
rect 116000 135346 118000 135666
rect 522000 135624 578864 135666
rect 522000 135388 524250 135624
rect 524486 135388 534250 135624
rect 534486 135388 544250 135624
rect 544486 135388 554250 135624
rect 554486 135388 564250 135624
rect 564486 135388 574250 135624
rect 574486 135388 578864 135624
rect 522000 135346 578864 135388
rect 1104 122346 2000 122666
rect 116000 122346 118000 122666
rect 522000 122624 578864 122666
rect 522000 122388 529250 122624
rect 529486 122388 539250 122624
rect 539486 122388 549250 122624
rect 549486 122388 559250 122624
rect 559486 122388 569250 122624
rect 569486 122388 578864 122624
rect 522000 122346 578864 122388
rect 1104 109346 2000 109666
rect 116000 109346 118000 109666
rect 522000 109624 578864 109666
rect 522000 109388 524250 109624
rect 524486 109388 534250 109624
rect 534486 109388 544250 109624
rect 544486 109388 554250 109624
rect 554486 109388 564250 109624
rect 564486 109388 574250 109624
rect 574486 109388 578864 109624
rect 522000 109346 578864 109388
rect 1104 96346 2000 96666
rect 116000 96346 118000 96666
rect 522000 96624 578864 96666
rect 522000 96388 529250 96624
rect 529486 96388 539250 96624
rect 539486 96388 549250 96624
rect 549486 96388 559250 96624
rect 559486 96388 569250 96624
rect 569486 96388 578864 96624
rect 522000 96346 578864 96388
rect 1104 83346 2000 83666
rect 116000 83346 118000 83666
rect 522000 83624 578864 83666
rect 522000 83388 524250 83624
rect 524486 83388 534250 83624
rect 534486 83388 544250 83624
rect 544486 83388 554250 83624
rect 554486 83388 564250 83624
rect 564486 83388 574250 83624
rect 574486 83388 578864 83624
rect 522000 83346 578864 83388
rect 512556 75258 521892 75300
rect 512556 75022 521614 75258
rect 521850 75022 521892 75258
rect 512556 74980 521892 75022
rect 512556 74620 512876 74980
rect 123212 74300 512876 74620
rect 123212 73940 123532 74300
rect 116772 73898 123532 73940
rect 116772 73662 116814 73898
rect 117050 73662 123532 73898
rect 116772 73620 123532 73662
rect 1104 70346 2000 70666
rect 116000 70346 118000 70666
rect 522000 70624 578864 70666
rect 522000 70388 529250 70624
rect 529486 70388 539250 70624
rect 539486 70388 549250 70624
rect 549486 70388 559250 70624
rect 559486 70388 569250 70624
rect 569486 70388 578864 70624
rect 522000 70346 578864 70388
rect 116404 62338 123532 62380
rect 116404 62102 116446 62338
rect 116682 62102 123532 62338
rect 116404 62060 123532 62102
rect 123212 61700 123532 62060
rect 512740 62338 513060 62380
rect 512740 62102 512782 62338
rect 513018 62102 513060 62338
rect 512740 61700 513060 62102
rect 123212 61380 513060 61700
rect 512740 59618 520420 59660
rect 512740 59382 512782 59618
rect 513018 59382 520142 59618
rect 520378 59382 520420 59618
rect 512740 59340 520420 59382
rect 1104 57346 2000 57666
rect 116000 57346 118000 57666
rect 522000 57624 578864 57666
rect 522000 57388 524250 57624
rect 524486 57388 534250 57624
rect 534486 57388 544250 57624
rect 544486 57388 554250 57624
rect 554486 57388 564250 57624
rect 564486 57388 574250 57624
rect 574486 57388 578864 57624
rect 522000 57346 578864 57388
rect 1104 44346 2000 44666
rect 116000 44346 118000 44666
rect 522000 44624 578864 44666
rect 522000 44388 529250 44624
rect 529486 44388 539250 44624
rect 539486 44388 549250 44624
rect 549486 44388 559250 44624
rect 559486 44388 569250 44624
rect 569486 44388 578864 44624
rect 522000 44346 578864 44388
rect 1104 31346 2000 31666
rect 116000 31346 118000 31666
rect 522000 31624 578864 31666
rect 522000 31388 524250 31624
rect 524486 31388 534250 31624
rect 534486 31388 544250 31624
rect 544486 31388 554250 31624
rect 554486 31388 564250 31624
rect 564486 31388 574250 31624
rect 574486 31388 578864 31624
rect 522000 31346 578864 31388
rect 512740 23578 522260 23620
rect 512740 23342 512782 23578
rect 513018 23342 521982 23578
rect 522218 23342 522260 23578
rect 512740 23300 522260 23342
rect 116772 22218 119668 22260
rect 116772 21982 116814 22218
rect 117050 21982 119668 22218
rect 116772 21940 119668 21982
rect 119348 21580 119668 21940
rect 119348 21538 513060 21580
rect 119348 21302 512782 21538
rect 513018 21302 513060 21538
rect 119348 21260 513060 21302
rect 518720 21538 521892 21580
rect 518720 21302 521614 21538
rect 521850 21302 521892 21538
rect 518720 21260 521892 21302
rect 518720 20900 519040 21260
rect 116404 20858 519040 20900
rect 116404 20622 116446 20858
rect 116682 20622 519040 20858
rect 116404 20580 519040 20622
rect 1104 18346 2000 18666
rect 116000 18346 118000 18666
rect 522000 18624 578864 18666
rect 522000 18388 529250 18624
rect 529486 18388 539250 18624
rect 539486 18388 549250 18624
rect 549486 18388 559250 18624
rect 559486 18388 569250 18624
rect 569486 18388 578864 18624
rect 522000 18346 578864 18388
rect 1104 5346 2000 5666
rect 116000 5346 118000 5666
rect 522000 5624 578864 5666
rect 522000 5388 524250 5624
rect 524486 5388 534250 5624
rect 534486 5388 544250 5624
rect 544486 5388 554250 5624
rect 554486 5388 564250 5624
rect 564486 5388 574250 5624
rect 574486 5388 578864 5624
rect 522000 5346 578864 5388
use mgmt_core  core
timestamp 1638138710
transform 1 0 120000 0 1 4000
box 0 0 400000 148000
use DFFRAM  DFFRAM
timestamp 1638138710
transform 1 0 4000 0 1 4000
box 4 0 110000 148000
<< labels >>
rlabel metal5 s 1104 18346 2000 18666 6 VGND
port 0 nsew ground input
rlabel metal5 s 116000 18346 118000 18666 6 VGND
port 0 nsew ground input
rlabel metal5 s 522000 18346 578864 18666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 44346 2000 44666 6 VGND
port 0 nsew ground input
rlabel metal5 s 116000 44346 118000 44666 6 VGND
port 0 nsew ground input
rlabel metal5 s 522000 44346 578864 44666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 70346 2000 70666 6 VGND
port 0 nsew ground input
rlabel metal5 s 116000 70346 118000 70666 6 VGND
port 0 nsew ground input
rlabel metal5 s 522000 70346 578864 70666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 96346 2000 96666 6 VGND
port 0 nsew ground input
rlabel metal5 s 116000 96346 118000 96666 6 VGND
port 0 nsew ground input
rlabel metal5 s 522000 96346 578864 96666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 122346 2000 122666 6 VGND
port 0 nsew ground input
rlabel metal5 s 116000 122346 118000 122666 6 VGND
port 0 nsew ground input
rlabel metal5 s 522000 122346 578864 122666 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 148346 2000 148666 6 VGND
port 0 nsew ground input
rlabel metal5 s 116000 148346 118000 148666 6 VGND
port 0 nsew ground input
rlabel metal5 s 522000 148346 578864 148666 6 VGND
port 0 nsew ground input
rlabel metal4 s 9208 154000 9528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 19208 154000 19528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 29208 154000 29528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 39208 154000 39528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 49208 154000 49528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 59208 154000 59528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 69208 154000 69528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 79208 154000 79528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 89208 154000 89528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 99208 154000 99528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 109208 154000 109528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 119208 154000 119528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 129208 154000 129528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 139208 154000 139528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 149208 154000 149528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 159208 154000 159528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 169208 154000 169528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 179208 154000 179528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 189208 154000 189528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 199208 154000 199528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 209208 154000 209528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 219208 154000 219528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 229208 154000 229528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 239208 154000 239528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 249208 154000 249528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 259208 154000 259528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 269208 154000 269528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 279208 154000 279528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 289208 154000 289528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 299208 154000 299528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 309208 154000 309528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 319208 154000 319528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 329208 154000 329528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 339208 154000 339528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 349208 154000 349528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 359208 154000 359528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 369208 154000 369528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 379208 154000 379528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 389208 154000 389528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 399208 154000 399528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 409208 154000 409528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 419208 154000 419528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 429208 154000 429528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 439208 154000 439528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 449208 154000 449528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 459208 154000 459528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 469208 154000 469528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 479208 154000 479528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 489208 154000 489528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 499208 154000 499528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 509208 154000 509528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 519208 154000 519528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 529208 2176 529528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 539208 2176 539528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 549208 2176 549528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 559208 2176 559528 157760 6 VGND
port 0 nsew ground input
rlabel metal4 s 569208 2176 569528 157760 6 VGND
port 0 nsew ground input
rlabel metal5 s 1104 5346 2000 5666 6 VPWR
port 1 nsew power input
rlabel metal5 s 116000 5346 118000 5666 6 VPWR
port 1 nsew power input
rlabel metal5 s 522000 5346 578864 5666 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 31346 2000 31666 6 VPWR
port 1 nsew power input
rlabel metal5 s 116000 31346 118000 31666 6 VPWR
port 1 nsew power input
rlabel metal5 s 522000 31346 578864 31666 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 57346 2000 57666 6 VPWR
port 1 nsew power input
rlabel metal5 s 116000 57346 118000 57666 6 VPWR
port 1 nsew power input
rlabel metal5 s 522000 57346 578864 57666 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 83346 2000 83666 6 VPWR
port 1 nsew power input
rlabel metal5 s 116000 83346 118000 83666 6 VPWR
port 1 nsew power input
rlabel metal5 s 522000 83346 578864 83666 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 109346 2000 109666 6 VPWR
port 1 nsew power input
rlabel metal5 s 116000 109346 118000 109666 6 VPWR
port 1 nsew power input
rlabel metal5 s 522000 109346 578864 109666 6 VPWR
port 1 nsew power input
rlabel metal5 s 1104 135346 2000 135666 6 VPWR
port 1 nsew power input
rlabel metal5 s 116000 135346 118000 135666 6 VPWR
port 1 nsew power input
rlabel metal5 s 522000 135346 578864 135666 6 VPWR
port 1 nsew power input
rlabel metal4 s 4208 154000 4528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 14208 154000 14528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 24208 154000 24528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 34208 154000 34528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 44208 154000 44528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 54208 154000 54528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 64208 154000 64528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 74208 154000 74528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 84208 154000 84528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 94208 154000 94528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 104208 154000 104528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 114208 154000 114528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 124208 154000 124528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 134208 154000 134528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 144208 154000 144528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 154208 154000 154528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 164208 154000 164528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 174208 154000 174528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 184208 154000 184528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 194208 154000 194528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 204208 154000 204528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 214208 154000 214528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 224208 154000 224528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 234208 154000 234528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 244208 154000 244528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 254208 154000 254528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 264208 154000 264528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 274208 154000 274528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 284208 154000 284528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 294208 154000 294528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 304208 154000 304528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 314208 154000 314528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 324208 154000 324528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 334208 154000 334528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 344208 154000 344528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 354208 154000 354528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 364208 154000 364528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 374208 154000 374528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 384208 154000 384528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 394208 154000 394528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 404208 154000 404528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 414208 154000 414528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 424208 154000 424528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 434208 154000 434528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 444208 154000 444528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 454208 154000 454528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 464208 154000 464528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 474208 154000 474528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 484208 154000 484528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 494208 154000 494528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 504208 154000 504528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 514208 154000 514528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 524208 2176 524528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 534208 2176 534528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 544208 2176 544528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 554208 2176 554528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 564208 2176 564528 157760 6 VPWR
port 1 nsew power input
rlabel metal4 s 574208 2176 574528 157760 6 VPWR
port 1 nsew power input
rlabel metal2 s 478 159200 534 160000 6 core_clk
port 2 nsew signal input
rlabel metal2 s 1398 159200 1454 160000 6 core_rstn
port 3 nsew signal input
rlabel metal2 s 508042 0 508098 800 6 debug_in
port 4 nsew signal input
rlabel metal2 s 513378 0 513434 800 6 debug_mode
port 5 nsew signal tristate
rlabel metal2 s 523958 0 524014 800 6 debug_oeb
port 6 nsew signal tristate
rlabel metal2 s 518622 0 518678 800 6 debug_out
port 7 nsew signal tristate
rlabel metal2 s 39762 0 39818 800 6 flash_clk
port 8 nsew signal tristate
rlabel metal2 s 34518 0 34574 800 6 flash_csb
port 9 nsew signal tristate
rlabel metal2 s 45098 0 45154 800 6 flash_io0_di
port 10 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 flash_io0_do
port 11 nsew signal tristate
rlabel metal2 s 55770 0 55826 800 6 flash_io0_oeb
port 12 nsew signal tristate
rlabel metal2 s 61106 0 61162 800 6 flash_io1_di
port 13 nsew signal input
rlabel metal2 s 66442 0 66498 800 6 flash_io1_do
port 14 nsew signal tristate
rlabel metal2 s 71686 0 71742 800 6 flash_io1_oeb
port 15 nsew signal tristate
rlabel metal2 s 77022 0 77078 800 6 flash_io2_di
port 16 nsew signal input
rlabel metal2 s 82358 0 82414 800 6 flash_io2_do
port 17 nsew signal tristate
rlabel metal3 s 0 6672 800 6792 6 flash_io2_oeb
port 18 nsew signal tristate
rlabel metal2 s 87694 0 87750 800 6 flash_io3_di
port 19 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 flash_io3_do
port 20 nsew signal tristate
rlabel metal3 s 0 2184 800 2304 6 flash_io3_oeb
port 21 nsew signal tristate
rlabel metal2 s 2594 0 2650 800 6 gpio_in_pad
port 22 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 gpio_inenb_pad
port 23 nsew signal tristate
rlabel metal2 s 13174 0 13230 800 6 gpio_mode0_pad
port 24 nsew signal tristate
rlabel metal2 s 18510 0 18566 800 6 gpio_mode1_pad
port 25 nsew signal tristate
rlabel metal2 s 23846 0 23902 800 6 gpio_out_pad
port 26 nsew signal tristate
rlabel metal2 s 29182 0 29238 800 6 gpio_outenb_pad
port 27 nsew signal tristate
rlabel metal2 s 103610 0 103666 800 6 hk_ack_i
port 28 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 hk_dat_i[0]
port 29 nsew signal input
rlabel metal2 s 167458 0 167514 800 6 hk_dat_i[10]
port 30 nsew signal input
rlabel metal2 s 172794 0 172850 800 6 hk_dat_i[11]
port 31 nsew signal input
rlabel metal2 s 178130 0 178186 800 6 hk_dat_i[12]
port 32 nsew signal input
rlabel metal2 s 183466 0 183522 800 6 hk_dat_i[13]
port 33 nsew signal input
rlabel metal2 s 188802 0 188858 800 6 hk_dat_i[14]
port 34 nsew signal input
rlabel metal2 s 194138 0 194194 800 6 hk_dat_i[15]
port 35 nsew signal input
rlabel metal2 s 199382 0 199438 800 6 hk_dat_i[16]
port 36 nsew signal input
rlabel metal2 s 204718 0 204774 800 6 hk_dat_i[17]
port 37 nsew signal input
rlabel metal2 s 210054 0 210110 800 6 hk_dat_i[18]
port 38 nsew signal input
rlabel metal2 s 215390 0 215446 800 6 hk_dat_i[19]
port 39 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 hk_dat_i[1]
port 40 nsew signal input
rlabel metal2 s 220726 0 220782 800 6 hk_dat_i[20]
port 41 nsew signal input
rlabel metal2 s 226062 0 226118 800 6 hk_dat_i[21]
port 42 nsew signal input
rlabel metal2 s 231306 0 231362 800 6 hk_dat_i[22]
port 43 nsew signal input
rlabel metal2 s 236642 0 236698 800 6 hk_dat_i[23]
port 44 nsew signal input
rlabel metal2 s 241978 0 242034 800 6 hk_dat_i[24]
port 45 nsew signal input
rlabel metal2 s 247314 0 247370 800 6 hk_dat_i[25]
port 46 nsew signal input
rlabel metal2 s 252650 0 252706 800 6 hk_dat_i[26]
port 47 nsew signal input
rlabel metal2 s 257986 0 258042 800 6 hk_dat_i[27]
port 48 nsew signal input
rlabel metal2 s 263230 0 263286 800 6 hk_dat_i[28]
port 49 nsew signal input
rlabel metal2 s 268566 0 268622 800 6 hk_dat_i[29]
port 50 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 hk_dat_i[2]
port 51 nsew signal input
rlabel metal2 s 273902 0 273958 800 6 hk_dat_i[30]
port 52 nsew signal input
rlabel metal2 s 279238 0 279294 800 6 hk_dat_i[31]
port 53 nsew signal input
rlabel metal2 s 130290 0 130346 800 6 hk_dat_i[3]
port 54 nsew signal input
rlabel metal2 s 135534 0 135590 800 6 hk_dat_i[4]
port 55 nsew signal input
rlabel metal2 s 140870 0 140926 800 6 hk_dat_i[5]
port 56 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 hk_dat_i[6]
port 57 nsew signal input
rlabel metal2 s 151542 0 151598 800 6 hk_dat_i[7]
port 58 nsew signal input
rlabel metal2 s 156878 0 156934 800 6 hk_dat_i[8]
port 59 nsew signal input
rlabel metal2 s 162214 0 162270 800 6 hk_dat_i[9]
port 60 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 hk_stb_o
port 61 nsew signal tristate
rlabel metal2 s 574558 159200 574614 160000 6 irq[0]
port 62 nsew signal input
rlabel metal2 s 575570 159200 575626 160000 6 irq[1]
port 63 nsew signal input
rlabel metal2 s 576490 159200 576546 160000 6 irq[2]
port 64 nsew signal input
rlabel metal2 s 577502 159200 577558 160000 6 irq[3]
port 65 nsew signal input
rlabel metal2 s 578422 159200 578478 160000 6 irq[4]
port 66 nsew signal input
rlabel metal2 s 579434 159200 579490 160000 6 irq[5]
port 67 nsew signal input
rlabel metal2 s 2410 159200 2466 160000 6 la_iena[0]
port 68 nsew signal tristate
rlabel metal2 s 392306 159200 392362 160000 6 la_iena[100]
port 69 nsew signal tristate
rlabel metal2 s 396170 159200 396226 160000 6 la_iena[101]
port 70 nsew signal tristate
rlabel metal2 s 400034 159200 400090 160000 6 la_iena[102]
port 71 nsew signal tristate
rlabel metal2 s 403990 159200 404046 160000 6 la_iena[103]
port 72 nsew signal tristate
rlabel metal2 s 407854 159200 407910 160000 6 la_iena[104]
port 73 nsew signal tristate
rlabel metal2 s 411810 159200 411866 160000 6 la_iena[105]
port 74 nsew signal tristate
rlabel metal2 s 415674 159200 415730 160000 6 la_iena[106]
port 75 nsew signal tristate
rlabel metal2 s 419538 159200 419594 160000 6 la_iena[107]
port 76 nsew signal tristate
rlabel metal2 s 423494 159200 423550 160000 6 la_iena[108]
port 77 nsew signal tristate
rlabel metal2 s 427358 159200 427414 160000 6 la_iena[109]
port 78 nsew signal tristate
rlabel metal2 s 41326 159200 41382 160000 6 la_iena[10]
port 79 nsew signal tristate
rlabel metal2 s 431222 159200 431278 160000 6 la_iena[110]
port 80 nsew signal tristate
rlabel metal2 s 435178 159200 435234 160000 6 la_iena[111]
port 81 nsew signal tristate
rlabel metal2 s 439042 159200 439098 160000 6 la_iena[112]
port 82 nsew signal tristate
rlabel metal2 s 442998 159200 443054 160000 6 la_iena[113]
port 83 nsew signal tristate
rlabel metal2 s 446862 159200 446918 160000 6 la_iena[114]
port 84 nsew signal tristate
rlabel metal2 s 450726 159200 450782 160000 6 la_iena[115]
port 85 nsew signal tristate
rlabel metal2 s 454682 159200 454738 160000 6 la_iena[116]
port 86 nsew signal tristate
rlabel metal2 s 458546 159200 458602 160000 6 la_iena[117]
port 87 nsew signal tristate
rlabel metal2 s 462502 159200 462558 160000 6 la_iena[118]
port 88 nsew signal tristate
rlabel metal2 s 466366 159200 466422 160000 6 la_iena[119]
port 89 nsew signal tristate
rlabel metal2 s 45282 159200 45338 160000 6 la_iena[11]
port 90 nsew signal tristate
rlabel metal2 s 470230 159200 470286 160000 6 la_iena[120]
port 91 nsew signal tristate
rlabel metal2 s 474186 159200 474242 160000 6 la_iena[121]
port 92 nsew signal tristate
rlabel metal2 s 478050 159200 478106 160000 6 la_iena[122]
port 93 nsew signal tristate
rlabel metal2 s 481914 159200 481970 160000 6 la_iena[123]
port 94 nsew signal tristate
rlabel metal2 s 485870 159200 485926 160000 6 la_iena[124]
port 95 nsew signal tristate
rlabel metal2 s 489734 159200 489790 160000 6 la_iena[125]
port 96 nsew signal tristate
rlabel metal2 s 493690 159200 493746 160000 6 la_iena[126]
port 97 nsew signal tristate
rlabel metal2 s 497554 159200 497610 160000 6 la_iena[127]
port 98 nsew signal tristate
rlabel metal2 s 49146 159200 49202 160000 6 la_iena[12]
port 99 nsew signal tristate
rlabel metal2 s 53102 159200 53158 160000 6 la_iena[13]
port 100 nsew signal tristate
rlabel metal2 s 56966 159200 57022 160000 6 la_iena[14]
port 101 nsew signal tristate
rlabel metal2 s 60830 159200 60886 160000 6 la_iena[15]
port 102 nsew signal tristate
rlabel metal2 s 64786 159200 64842 160000 6 la_iena[16]
port 103 nsew signal tristate
rlabel metal2 s 68650 159200 68706 160000 6 la_iena[17]
port 104 nsew signal tristate
rlabel metal2 s 72606 159200 72662 160000 6 la_iena[18]
port 105 nsew signal tristate
rlabel metal2 s 76470 159200 76526 160000 6 la_iena[19]
port 106 nsew signal tristate
rlabel metal2 s 6274 159200 6330 160000 6 la_iena[1]
port 107 nsew signal tristate
rlabel metal2 s 80334 159200 80390 160000 6 la_iena[20]
port 108 nsew signal tristate
rlabel metal2 s 84290 159200 84346 160000 6 la_iena[21]
port 109 nsew signal tristate
rlabel metal2 s 88154 159200 88210 160000 6 la_iena[22]
port 110 nsew signal tristate
rlabel metal2 s 92018 159200 92074 160000 6 la_iena[23]
port 111 nsew signal tristate
rlabel metal2 s 95974 159200 96030 160000 6 la_iena[24]
port 112 nsew signal tristate
rlabel metal2 s 99838 159200 99894 160000 6 la_iena[25]
port 113 nsew signal tristate
rlabel metal2 s 103794 159200 103850 160000 6 la_iena[26]
port 114 nsew signal tristate
rlabel metal2 s 107658 159200 107714 160000 6 la_iena[27]
port 115 nsew signal tristate
rlabel metal2 s 111522 159200 111578 160000 6 la_iena[28]
port 116 nsew signal tristate
rlabel metal2 s 115478 159200 115534 160000 6 la_iena[29]
port 117 nsew signal tristate
rlabel metal2 s 10138 159200 10194 160000 6 la_iena[2]
port 118 nsew signal tristate
rlabel metal2 s 119342 159200 119398 160000 6 la_iena[30]
port 119 nsew signal tristate
rlabel metal2 s 123206 159200 123262 160000 6 la_iena[31]
port 120 nsew signal tristate
rlabel metal2 s 127162 159200 127218 160000 6 la_iena[32]
port 121 nsew signal tristate
rlabel metal2 s 131026 159200 131082 160000 6 la_iena[33]
port 122 nsew signal tristate
rlabel metal2 s 134982 159200 135038 160000 6 la_iena[34]
port 123 nsew signal tristate
rlabel metal2 s 138846 159200 138902 160000 6 la_iena[35]
port 124 nsew signal tristate
rlabel metal2 s 142710 159200 142766 160000 6 la_iena[36]
port 125 nsew signal tristate
rlabel metal2 s 146666 159200 146722 160000 6 la_iena[37]
port 126 nsew signal tristate
rlabel metal2 s 150530 159200 150586 160000 6 la_iena[38]
port 127 nsew signal tristate
rlabel metal2 s 154486 159200 154542 160000 6 la_iena[39]
port 128 nsew signal tristate
rlabel metal2 s 14094 159200 14150 160000 6 la_iena[3]
port 129 nsew signal tristate
rlabel metal2 s 158350 159200 158406 160000 6 la_iena[40]
port 130 nsew signal tristate
rlabel metal2 s 162214 159200 162270 160000 6 la_iena[41]
port 131 nsew signal tristate
rlabel metal2 s 166170 159200 166226 160000 6 la_iena[42]
port 132 nsew signal tristate
rlabel metal2 s 170034 159200 170090 160000 6 la_iena[43]
port 133 nsew signal tristate
rlabel metal2 s 173898 159200 173954 160000 6 la_iena[44]
port 134 nsew signal tristate
rlabel metal2 s 177854 159200 177910 160000 6 la_iena[45]
port 135 nsew signal tristate
rlabel metal2 s 181718 159200 181774 160000 6 la_iena[46]
port 136 nsew signal tristate
rlabel metal2 s 185674 159200 185730 160000 6 la_iena[47]
port 137 nsew signal tristate
rlabel metal2 s 189538 159200 189594 160000 6 la_iena[48]
port 138 nsew signal tristate
rlabel metal2 s 193402 159200 193458 160000 6 la_iena[49]
port 139 nsew signal tristate
rlabel metal2 s 17958 159200 18014 160000 6 la_iena[4]
port 140 nsew signal tristate
rlabel metal2 s 197358 159200 197414 160000 6 la_iena[50]
port 141 nsew signal tristate
rlabel metal2 s 201222 159200 201278 160000 6 la_iena[51]
port 142 nsew signal tristate
rlabel metal2 s 205086 159200 205142 160000 6 la_iena[52]
port 143 nsew signal tristate
rlabel metal2 s 209042 159200 209098 160000 6 la_iena[53]
port 144 nsew signal tristate
rlabel metal2 s 212906 159200 212962 160000 6 la_iena[54]
port 145 nsew signal tristate
rlabel metal2 s 216862 159200 216918 160000 6 la_iena[55]
port 146 nsew signal tristate
rlabel metal2 s 220726 159200 220782 160000 6 la_iena[56]
port 147 nsew signal tristate
rlabel metal2 s 224590 159200 224646 160000 6 la_iena[57]
port 148 nsew signal tristate
rlabel metal2 s 228546 159200 228602 160000 6 la_iena[58]
port 149 nsew signal tristate
rlabel metal2 s 232410 159200 232466 160000 6 la_iena[59]
port 150 nsew signal tristate
rlabel metal2 s 21914 159200 21970 160000 6 la_iena[5]
port 151 nsew signal tristate
rlabel metal2 s 236274 159200 236330 160000 6 la_iena[60]
port 152 nsew signal tristate
rlabel metal2 s 240230 159200 240286 160000 6 la_iena[61]
port 153 nsew signal tristate
rlabel metal2 s 244094 159200 244150 160000 6 la_iena[62]
port 154 nsew signal tristate
rlabel metal2 s 248050 159200 248106 160000 6 la_iena[63]
port 155 nsew signal tristate
rlabel metal2 s 251914 159200 251970 160000 6 la_iena[64]
port 156 nsew signal tristate
rlabel metal2 s 255778 159200 255834 160000 6 la_iena[65]
port 157 nsew signal tristate
rlabel metal2 s 259734 159200 259790 160000 6 la_iena[66]
port 158 nsew signal tristate
rlabel metal2 s 263598 159200 263654 160000 6 la_iena[67]
port 159 nsew signal tristate
rlabel metal2 s 267554 159200 267610 160000 6 la_iena[68]
port 160 nsew signal tristate
rlabel metal2 s 271418 159200 271474 160000 6 la_iena[69]
port 161 nsew signal tristate
rlabel metal2 s 25778 159200 25834 160000 6 la_iena[6]
port 162 nsew signal tristate
rlabel metal2 s 275282 159200 275338 160000 6 la_iena[70]
port 163 nsew signal tristate
rlabel metal2 s 279238 159200 279294 160000 6 la_iena[71]
port 164 nsew signal tristate
rlabel metal2 s 283102 159200 283158 160000 6 la_iena[72]
port 165 nsew signal tristate
rlabel metal2 s 286966 159200 287022 160000 6 la_iena[73]
port 166 nsew signal tristate
rlabel metal2 s 290922 159200 290978 160000 6 la_iena[74]
port 167 nsew signal tristate
rlabel metal2 s 294786 159200 294842 160000 6 la_iena[75]
port 168 nsew signal tristate
rlabel metal2 s 298742 159200 298798 160000 6 la_iena[76]
port 169 nsew signal tristate
rlabel metal2 s 302606 159200 302662 160000 6 la_iena[77]
port 170 nsew signal tristate
rlabel metal2 s 306470 159200 306526 160000 6 la_iena[78]
port 171 nsew signal tristate
rlabel metal2 s 310426 159200 310482 160000 6 la_iena[79]
port 172 nsew signal tristate
rlabel metal2 s 29642 159200 29698 160000 6 la_iena[7]
port 173 nsew signal tristate
rlabel metal2 s 314290 159200 314346 160000 6 la_iena[80]
port 174 nsew signal tristate
rlabel metal2 s 318154 159200 318210 160000 6 la_iena[81]
port 175 nsew signal tristate
rlabel metal2 s 322110 159200 322166 160000 6 la_iena[82]
port 176 nsew signal tristate
rlabel metal2 s 325974 159200 326030 160000 6 la_iena[83]
port 177 nsew signal tristate
rlabel metal2 s 329930 159200 329986 160000 6 la_iena[84]
port 178 nsew signal tristate
rlabel metal2 s 333794 159200 333850 160000 6 la_iena[85]
port 179 nsew signal tristate
rlabel metal2 s 337658 159200 337714 160000 6 la_iena[86]
port 180 nsew signal tristate
rlabel metal2 s 341614 159200 341670 160000 6 la_iena[87]
port 181 nsew signal tristate
rlabel metal2 s 345478 159200 345534 160000 6 la_iena[88]
port 182 nsew signal tristate
rlabel metal2 s 349342 159200 349398 160000 6 la_iena[89]
port 183 nsew signal tristate
rlabel metal2 s 33598 159200 33654 160000 6 la_iena[8]
port 184 nsew signal tristate
rlabel metal2 s 353298 159200 353354 160000 6 la_iena[90]
port 185 nsew signal tristate
rlabel metal2 s 357162 159200 357218 160000 6 la_iena[91]
port 186 nsew signal tristate
rlabel metal2 s 361118 159200 361174 160000 6 la_iena[92]
port 187 nsew signal tristate
rlabel metal2 s 364982 159200 365038 160000 6 la_iena[93]
port 188 nsew signal tristate
rlabel metal2 s 368846 159200 368902 160000 6 la_iena[94]
port 189 nsew signal tristate
rlabel metal2 s 372802 159200 372858 160000 6 la_iena[95]
port 190 nsew signal tristate
rlabel metal2 s 376666 159200 376722 160000 6 la_iena[96]
port 191 nsew signal tristate
rlabel metal2 s 380622 159200 380678 160000 6 la_iena[97]
port 192 nsew signal tristate
rlabel metal2 s 384486 159200 384542 160000 6 la_iena[98]
port 193 nsew signal tristate
rlabel metal2 s 388350 159200 388406 160000 6 la_iena[99]
port 194 nsew signal tristate
rlabel metal2 s 37462 159200 37518 160000 6 la_iena[9]
port 195 nsew signal tristate
rlabel metal2 s 3330 159200 3386 160000 6 la_input[0]
port 196 nsew signal input
rlabel metal2 s 393226 159200 393282 160000 6 la_input[100]
port 197 nsew signal input
rlabel metal2 s 397182 159200 397238 160000 6 la_input[101]
port 198 nsew signal input
rlabel metal2 s 401046 159200 401102 160000 6 la_input[102]
port 199 nsew signal input
rlabel metal2 s 404910 159200 404966 160000 6 la_input[103]
port 200 nsew signal input
rlabel metal2 s 408866 159200 408922 160000 6 la_input[104]
port 201 nsew signal input
rlabel metal2 s 412730 159200 412786 160000 6 la_input[105]
port 202 nsew signal input
rlabel metal2 s 416686 159200 416742 160000 6 la_input[106]
port 203 nsew signal input
rlabel metal2 s 420550 159200 420606 160000 6 la_input[107]
port 204 nsew signal input
rlabel metal2 s 424414 159200 424470 160000 6 la_input[108]
port 205 nsew signal input
rlabel metal2 s 428370 159200 428426 160000 6 la_input[109]
port 206 nsew signal input
rlabel metal2 s 42338 159200 42394 160000 6 la_input[10]
port 207 nsew signal input
rlabel metal2 s 432234 159200 432290 160000 6 la_input[110]
port 208 nsew signal input
rlabel metal2 s 436098 159200 436154 160000 6 la_input[111]
port 209 nsew signal input
rlabel metal2 s 440054 159200 440110 160000 6 la_input[112]
port 210 nsew signal input
rlabel metal2 s 443918 159200 443974 160000 6 la_input[113]
port 211 nsew signal input
rlabel metal2 s 447874 159200 447930 160000 6 la_input[114]
port 212 nsew signal input
rlabel metal2 s 451738 159200 451794 160000 6 la_input[115]
port 213 nsew signal input
rlabel metal2 s 455602 159200 455658 160000 6 la_input[116]
port 214 nsew signal input
rlabel metal2 s 459558 159200 459614 160000 6 la_input[117]
port 215 nsew signal input
rlabel metal2 s 463422 159200 463478 160000 6 la_input[118]
port 216 nsew signal input
rlabel metal2 s 467286 159200 467342 160000 6 la_input[119]
port 217 nsew signal input
rlabel metal2 s 46202 159200 46258 160000 6 la_input[11]
port 218 nsew signal input
rlabel metal2 s 471242 159200 471298 160000 6 la_input[120]
port 219 nsew signal input
rlabel metal2 s 475106 159200 475162 160000 6 la_input[121]
port 220 nsew signal input
rlabel metal2 s 479062 159200 479118 160000 6 la_input[122]
port 221 nsew signal input
rlabel metal2 s 482926 159200 482982 160000 6 la_input[123]
port 222 nsew signal input
rlabel metal2 s 486790 159200 486846 160000 6 la_input[124]
port 223 nsew signal input
rlabel metal2 s 490746 159200 490802 160000 6 la_input[125]
port 224 nsew signal input
rlabel metal2 s 494610 159200 494666 160000 6 la_input[126]
port 225 nsew signal input
rlabel metal2 s 498566 159200 498622 160000 6 la_input[127]
port 226 nsew signal input
rlabel metal2 s 50158 159200 50214 160000 6 la_input[12]
port 227 nsew signal input
rlabel metal2 s 54022 159200 54078 160000 6 la_input[13]
port 228 nsew signal input
rlabel metal2 s 57978 159200 58034 160000 6 la_input[14]
port 229 nsew signal input
rlabel metal2 s 61842 159200 61898 160000 6 la_input[15]
port 230 nsew signal input
rlabel metal2 s 65706 159200 65762 160000 6 la_input[16]
port 231 nsew signal input
rlabel metal2 s 69662 159200 69718 160000 6 la_input[17]
port 232 nsew signal input
rlabel metal2 s 73526 159200 73582 160000 6 la_input[18]
port 233 nsew signal input
rlabel metal2 s 77482 159200 77538 160000 6 la_input[19]
port 234 nsew signal input
rlabel metal2 s 7286 159200 7342 160000 6 la_input[1]
port 235 nsew signal input
rlabel metal2 s 81346 159200 81402 160000 6 la_input[20]
port 236 nsew signal input
rlabel metal2 s 85210 159200 85266 160000 6 la_input[21]
port 237 nsew signal input
rlabel metal2 s 89166 159200 89222 160000 6 la_input[22]
port 238 nsew signal input
rlabel metal2 s 93030 159200 93086 160000 6 la_input[23]
port 239 nsew signal input
rlabel metal2 s 96894 159200 96950 160000 6 la_input[24]
port 240 nsew signal input
rlabel metal2 s 100850 159200 100906 160000 6 la_input[25]
port 241 nsew signal input
rlabel metal2 s 104714 159200 104770 160000 6 la_input[26]
port 242 nsew signal input
rlabel metal2 s 108670 159200 108726 160000 6 la_input[27]
port 243 nsew signal input
rlabel metal2 s 112534 159200 112590 160000 6 la_input[28]
port 244 nsew signal input
rlabel metal2 s 116398 159200 116454 160000 6 la_input[29]
port 245 nsew signal input
rlabel metal2 s 11150 159200 11206 160000 6 la_input[2]
port 246 nsew signal input
rlabel metal2 s 120354 159200 120410 160000 6 la_input[30]
port 247 nsew signal input
rlabel metal2 s 124218 159200 124274 160000 6 la_input[31]
port 248 nsew signal input
rlabel metal2 s 128082 159200 128138 160000 6 la_input[32]
port 249 nsew signal input
rlabel metal2 s 132038 159200 132094 160000 6 la_input[33]
port 250 nsew signal input
rlabel metal2 s 135902 159200 135958 160000 6 la_input[34]
port 251 nsew signal input
rlabel metal2 s 139858 159200 139914 160000 6 la_input[35]
port 252 nsew signal input
rlabel metal2 s 143722 159200 143778 160000 6 la_input[36]
port 253 nsew signal input
rlabel metal2 s 147586 159200 147642 160000 6 la_input[37]
port 254 nsew signal input
rlabel metal2 s 151542 159200 151598 160000 6 la_input[38]
port 255 nsew signal input
rlabel metal2 s 155406 159200 155462 160000 6 la_input[39]
port 256 nsew signal input
rlabel metal2 s 15014 159200 15070 160000 6 la_input[3]
port 257 nsew signal input
rlabel metal2 s 159270 159200 159326 160000 6 la_input[40]
port 258 nsew signal input
rlabel metal2 s 163226 159200 163282 160000 6 la_input[41]
port 259 nsew signal input
rlabel metal2 s 167090 159200 167146 160000 6 la_input[42]
port 260 nsew signal input
rlabel metal2 s 171046 159200 171102 160000 6 la_input[43]
port 261 nsew signal input
rlabel metal2 s 174910 159200 174966 160000 6 la_input[44]
port 262 nsew signal input
rlabel metal2 s 178774 159200 178830 160000 6 la_input[45]
port 263 nsew signal input
rlabel metal2 s 182730 159200 182786 160000 6 la_input[46]
port 264 nsew signal input
rlabel metal2 s 186594 159200 186650 160000 6 la_input[47]
port 265 nsew signal input
rlabel metal2 s 190550 159200 190606 160000 6 la_input[48]
port 266 nsew signal input
rlabel metal2 s 194414 159200 194470 160000 6 la_input[49]
port 267 nsew signal input
rlabel metal2 s 18970 159200 19026 160000 6 la_input[4]
port 268 nsew signal input
rlabel metal2 s 198278 159200 198334 160000 6 la_input[50]
port 269 nsew signal input
rlabel metal2 s 202234 159200 202290 160000 6 la_input[51]
port 270 nsew signal input
rlabel metal2 s 206098 159200 206154 160000 6 la_input[52]
port 271 nsew signal input
rlabel metal2 s 209962 159200 210018 160000 6 la_input[53]
port 272 nsew signal input
rlabel metal2 s 213918 159200 213974 160000 6 la_input[54]
port 273 nsew signal input
rlabel metal2 s 217782 159200 217838 160000 6 la_input[55]
port 274 nsew signal input
rlabel metal2 s 221738 159200 221794 160000 6 la_input[56]
port 275 nsew signal input
rlabel metal2 s 225602 159200 225658 160000 6 la_input[57]
port 276 nsew signal input
rlabel metal2 s 229466 159200 229522 160000 6 la_input[58]
port 277 nsew signal input
rlabel metal2 s 233422 159200 233478 160000 6 la_input[59]
port 278 nsew signal input
rlabel metal2 s 22834 159200 22890 160000 6 la_input[5]
port 279 nsew signal input
rlabel metal2 s 237286 159200 237342 160000 6 la_input[60]
port 280 nsew signal input
rlabel metal2 s 241150 159200 241206 160000 6 la_input[61]
port 281 nsew signal input
rlabel metal2 s 245106 159200 245162 160000 6 la_input[62]
port 282 nsew signal input
rlabel metal2 s 248970 159200 249026 160000 6 la_input[63]
port 283 nsew signal input
rlabel metal2 s 252926 159200 252982 160000 6 la_input[64]
port 284 nsew signal input
rlabel metal2 s 256790 159200 256846 160000 6 la_input[65]
port 285 nsew signal input
rlabel metal2 s 260654 159200 260710 160000 6 la_input[66]
port 286 nsew signal input
rlabel metal2 s 264610 159200 264666 160000 6 la_input[67]
port 287 nsew signal input
rlabel metal2 s 268474 159200 268530 160000 6 la_input[68]
port 288 nsew signal input
rlabel metal2 s 272338 159200 272394 160000 6 la_input[69]
port 289 nsew signal input
rlabel metal2 s 26790 159200 26846 160000 6 la_input[6]
port 290 nsew signal input
rlabel metal2 s 276294 159200 276350 160000 6 la_input[70]
port 291 nsew signal input
rlabel metal2 s 280158 159200 280214 160000 6 la_input[71]
port 292 nsew signal input
rlabel metal2 s 284114 159200 284170 160000 6 la_input[72]
port 293 nsew signal input
rlabel metal2 s 287978 159200 288034 160000 6 la_input[73]
port 294 nsew signal input
rlabel metal2 s 291842 159200 291898 160000 6 la_input[74]
port 295 nsew signal input
rlabel metal2 s 295798 159200 295854 160000 6 la_input[75]
port 296 nsew signal input
rlabel metal2 s 299662 159200 299718 160000 6 la_input[76]
port 297 nsew signal input
rlabel metal2 s 303618 159200 303674 160000 6 la_input[77]
port 298 nsew signal input
rlabel metal2 s 307482 159200 307538 160000 6 la_input[78]
port 299 nsew signal input
rlabel metal2 s 311346 159200 311402 160000 6 la_input[79]
port 300 nsew signal input
rlabel metal2 s 30654 159200 30710 160000 6 la_input[7]
port 301 nsew signal input
rlabel metal2 s 315302 159200 315358 160000 6 la_input[80]
port 302 nsew signal input
rlabel metal2 s 319166 159200 319222 160000 6 la_input[81]
port 303 nsew signal input
rlabel metal2 s 323030 159200 323086 160000 6 la_input[82]
port 304 nsew signal input
rlabel metal2 s 326986 159200 327042 160000 6 la_input[83]
port 305 nsew signal input
rlabel metal2 s 330850 159200 330906 160000 6 la_input[84]
port 306 nsew signal input
rlabel metal2 s 334806 159200 334862 160000 6 la_input[85]
port 307 nsew signal input
rlabel metal2 s 338670 159200 338726 160000 6 la_input[86]
port 308 nsew signal input
rlabel metal2 s 342534 159200 342590 160000 6 la_input[87]
port 309 nsew signal input
rlabel metal2 s 346490 159200 346546 160000 6 la_input[88]
port 310 nsew signal input
rlabel metal2 s 350354 159200 350410 160000 6 la_input[89]
port 311 nsew signal input
rlabel metal2 s 34518 159200 34574 160000 6 la_input[8]
port 312 nsew signal input
rlabel metal2 s 354218 159200 354274 160000 6 la_input[90]
port 313 nsew signal input
rlabel metal2 s 358174 159200 358230 160000 6 la_input[91]
port 314 nsew signal input
rlabel metal2 s 362038 159200 362094 160000 6 la_input[92]
port 315 nsew signal input
rlabel metal2 s 365994 159200 366050 160000 6 la_input[93]
port 316 nsew signal input
rlabel metal2 s 369858 159200 369914 160000 6 la_input[94]
port 317 nsew signal input
rlabel metal2 s 373722 159200 373778 160000 6 la_input[95]
port 318 nsew signal input
rlabel metal2 s 377678 159200 377734 160000 6 la_input[96]
port 319 nsew signal input
rlabel metal2 s 381542 159200 381598 160000 6 la_input[97]
port 320 nsew signal input
rlabel metal2 s 385498 159200 385554 160000 6 la_input[98]
port 321 nsew signal input
rlabel metal2 s 389362 159200 389418 160000 6 la_input[99]
port 322 nsew signal input
rlabel metal2 s 38474 159200 38530 160000 6 la_input[9]
port 323 nsew signal input
rlabel metal2 s 4342 159200 4398 160000 6 la_oenb[0]
port 324 nsew signal tristate
rlabel metal2 s 394238 159200 394294 160000 6 la_oenb[100]
port 325 nsew signal tristate
rlabel metal2 s 398102 159200 398158 160000 6 la_oenb[101]
port 326 nsew signal tristate
rlabel metal2 s 402058 159200 402114 160000 6 la_oenb[102]
port 327 nsew signal tristate
rlabel metal2 s 405922 159200 405978 160000 6 la_oenb[103]
port 328 nsew signal tristate
rlabel metal2 s 409786 159200 409842 160000 6 la_oenb[104]
port 329 nsew signal tristate
rlabel metal2 s 413742 159200 413798 160000 6 la_oenb[105]
port 330 nsew signal tristate
rlabel metal2 s 417606 159200 417662 160000 6 la_oenb[106]
port 331 nsew signal tristate
rlabel metal2 s 421562 159200 421618 160000 6 la_oenb[107]
port 332 nsew signal tristate
rlabel metal2 s 425426 159200 425482 160000 6 la_oenb[108]
port 333 nsew signal tristate
rlabel metal2 s 429290 159200 429346 160000 6 la_oenb[109]
port 334 nsew signal tristate
rlabel metal2 s 43350 159200 43406 160000 6 la_oenb[10]
port 335 nsew signal tristate
rlabel metal2 s 433246 159200 433302 160000 6 la_oenb[110]
port 336 nsew signal tristate
rlabel metal2 s 437110 159200 437166 160000 6 la_oenb[111]
port 337 nsew signal tristate
rlabel metal2 s 440974 159200 441030 160000 6 la_oenb[112]
port 338 nsew signal tristate
rlabel metal2 s 444930 159200 444986 160000 6 la_oenb[113]
port 339 nsew signal tristate
rlabel metal2 s 448794 159200 448850 160000 6 la_oenb[114]
port 340 nsew signal tristate
rlabel metal2 s 452750 159200 452806 160000 6 la_oenb[115]
port 341 nsew signal tristate
rlabel metal2 s 456614 159200 456670 160000 6 la_oenb[116]
port 342 nsew signal tristate
rlabel metal2 s 460478 159200 460534 160000 6 la_oenb[117]
port 343 nsew signal tristate
rlabel metal2 s 464434 159200 464490 160000 6 la_oenb[118]
port 344 nsew signal tristate
rlabel metal2 s 468298 159200 468354 160000 6 la_oenb[119]
port 345 nsew signal tristate
rlabel metal2 s 47214 159200 47270 160000 6 la_oenb[11]
port 346 nsew signal tristate
rlabel metal2 s 472162 159200 472218 160000 6 la_oenb[120]
port 347 nsew signal tristate
rlabel metal2 s 476118 159200 476174 160000 6 la_oenb[121]
port 348 nsew signal tristate
rlabel metal2 s 479982 159200 480038 160000 6 la_oenb[122]
port 349 nsew signal tristate
rlabel metal2 s 483938 159200 483994 160000 6 la_oenb[123]
port 350 nsew signal tristate
rlabel metal2 s 487802 159200 487858 160000 6 la_oenb[124]
port 351 nsew signal tristate
rlabel metal2 s 491666 159200 491722 160000 6 la_oenb[125]
port 352 nsew signal tristate
rlabel metal2 s 495622 159200 495678 160000 6 la_oenb[126]
port 353 nsew signal tristate
rlabel metal2 s 499486 159200 499542 160000 6 la_oenb[127]
port 354 nsew signal tristate
rlabel metal2 s 51078 159200 51134 160000 6 la_oenb[12]
port 355 nsew signal tristate
rlabel metal2 s 55034 159200 55090 160000 6 la_oenb[13]
port 356 nsew signal tristate
rlabel metal2 s 58898 159200 58954 160000 6 la_oenb[14]
port 357 nsew signal tristate
rlabel metal2 s 62854 159200 62910 160000 6 la_oenb[15]
port 358 nsew signal tristate
rlabel metal2 s 66718 159200 66774 160000 6 la_oenb[16]
port 359 nsew signal tristate
rlabel metal2 s 70582 159200 70638 160000 6 la_oenb[17]
port 360 nsew signal tristate
rlabel metal2 s 74538 159200 74594 160000 6 la_oenb[18]
port 361 nsew signal tristate
rlabel metal2 s 78402 159200 78458 160000 6 la_oenb[19]
port 362 nsew signal tristate
rlabel metal2 s 8206 159200 8262 160000 6 la_oenb[1]
port 363 nsew signal tristate
rlabel metal2 s 82266 159200 82322 160000 6 la_oenb[20]
port 364 nsew signal tristate
rlabel metal2 s 86222 159200 86278 160000 6 la_oenb[21]
port 365 nsew signal tristate
rlabel metal2 s 90086 159200 90142 160000 6 la_oenb[22]
port 366 nsew signal tristate
rlabel metal2 s 94042 159200 94098 160000 6 la_oenb[23]
port 367 nsew signal tristate
rlabel metal2 s 97906 159200 97962 160000 6 la_oenb[24]
port 368 nsew signal tristate
rlabel metal2 s 101770 159200 101826 160000 6 la_oenb[25]
port 369 nsew signal tristate
rlabel metal2 s 105726 159200 105782 160000 6 la_oenb[26]
port 370 nsew signal tristate
rlabel metal2 s 109590 159200 109646 160000 6 la_oenb[27]
port 371 nsew signal tristate
rlabel metal2 s 113546 159200 113602 160000 6 la_oenb[28]
port 372 nsew signal tristate
rlabel metal2 s 117410 159200 117466 160000 6 la_oenb[29]
port 373 nsew signal tristate
rlabel metal2 s 12162 159200 12218 160000 6 la_oenb[2]
port 374 nsew signal tristate
rlabel metal2 s 121274 159200 121330 160000 6 la_oenb[30]
port 375 nsew signal tristate
rlabel metal2 s 125230 159200 125286 160000 6 la_oenb[31]
port 376 nsew signal tristate
rlabel metal2 s 129094 159200 129150 160000 6 la_oenb[32]
port 377 nsew signal tristate
rlabel metal2 s 132958 159200 133014 160000 6 la_oenb[33]
port 378 nsew signal tristate
rlabel metal2 s 136914 159200 136970 160000 6 la_oenb[34]
port 379 nsew signal tristate
rlabel metal2 s 140778 159200 140834 160000 6 la_oenb[35]
port 380 nsew signal tristate
rlabel metal2 s 144734 159200 144790 160000 6 la_oenb[36]
port 381 nsew signal tristate
rlabel metal2 s 148598 159200 148654 160000 6 la_oenb[37]
port 382 nsew signal tristate
rlabel metal2 s 152462 159200 152518 160000 6 la_oenb[38]
port 383 nsew signal tristate
rlabel metal2 s 156418 159200 156474 160000 6 la_oenb[39]
port 384 nsew signal tristate
rlabel metal2 s 16026 159200 16082 160000 6 la_oenb[3]
port 385 nsew signal tristate
rlabel metal2 s 160282 159200 160338 160000 6 la_oenb[40]
port 386 nsew signal tristate
rlabel metal2 s 164146 159200 164202 160000 6 la_oenb[41]
port 387 nsew signal tristate
rlabel metal2 s 168102 159200 168158 160000 6 la_oenb[42]
port 388 nsew signal tristate
rlabel metal2 s 171966 159200 172022 160000 6 la_oenb[43]
port 389 nsew signal tristate
rlabel metal2 s 175922 159200 175978 160000 6 la_oenb[44]
port 390 nsew signal tristate
rlabel metal2 s 179786 159200 179842 160000 6 la_oenb[45]
port 391 nsew signal tristate
rlabel metal2 s 183650 159200 183706 160000 6 la_oenb[46]
port 392 nsew signal tristate
rlabel metal2 s 187606 159200 187662 160000 6 la_oenb[47]
port 393 nsew signal tristate
rlabel metal2 s 191470 159200 191526 160000 6 la_oenb[48]
port 394 nsew signal tristate
rlabel metal2 s 195334 159200 195390 160000 6 la_oenb[49]
port 395 nsew signal tristate
rlabel metal2 s 19890 159200 19946 160000 6 la_oenb[4]
port 396 nsew signal tristate
rlabel metal2 s 199290 159200 199346 160000 6 la_oenb[50]
port 397 nsew signal tristate
rlabel metal2 s 203154 159200 203210 160000 6 la_oenb[51]
port 398 nsew signal tristate
rlabel metal2 s 207110 159200 207166 160000 6 la_oenb[52]
port 399 nsew signal tristate
rlabel metal2 s 210974 159200 211030 160000 6 la_oenb[53]
port 400 nsew signal tristate
rlabel metal2 s 214838 159200 214894 160000 6 la_oenb[54]
port 401 nsew signal tristate
rlabel metal2 s 218794 159200 218850 160000 6 la_oenb[55]
port 402 nsew signal tristate
rlabel metal2 s 222658 159200 222714 160000 6 la_oenb[56]
port 403 nsew signal tristate
rlabel metal2 s 226614 159200 226670 160000 6 la_oenb[57]
port 404 nsew signal tristate
rlabel metal2 s 230478 159200 230534 160000 6 la_oenb[58]
port 405 nsew signal tristate
rlabel metal2 s 234342 159200 234398 160000 6 la_oenb[59]
port 406 nsew signal tristate
rlabel metal2 s 23846 159200 23902 160000 6 la_oenb[5]
port 407 nsew signal tristate
rlabel metal2 s 238298 159200 238354 160000 6 la_oenb[60]
port 408 nsew signal tristate
rlabel metal2 s 242162 159200 242218 160000 6 la_oenb[61]
port 409 nsew signal tristate
rlabel metal2 s 246026 159200 246082 160000 6 la_oenb[62]
port 410 nsew signal tristate
rlabel metal2 s 249982 159200 250038 160000 6 la_oenb[63]
port 411 nsew signal tristate
rlabel metal2 s 253846 159200 253902 160000 6 la_oenb[64]
port 412 nsew signal tristate
rlabel metal2 s 257802 159200 257858 160000 6 la_oenb[65]
port 413 nsew signal tristate
rlabel metal2 s 261666 159200 261722 160000 6 la_oenb[66]
port 414 nsew signal tristate
rlabel metal2 s 265530 159200 265586 160000 6 la_oenb[67]
port 415 nsew signal tristate
rlabel metal2 s 269486 159200 269542 160000 6 la_oenb[68]
port 416 nsew signal tristate
rlabel metal2 s 273350 159200 273406 160000 6 la_oenb[69]
port 417 nsew signal tristate
rlabel metal2 s 27710 159200 27766 160000 6 la_oenb[6]
port 418 nsew signal tristate
rlabel metal2 s 277214 159200 277270 160000 6 la_oenb[70]
port 419 nsew signal tristate
rlabel metal2 s 281170 159200 281226 160000 6 la_oenb[71]
port 420 nsew signal tristate
rlabel metal2 s 285034 159200 285090 160000 6 la_oenb[72]
port 421 nsew signal tristate
rlabel metal2 s 288990 159200 289046 160000 6 la_oenb[73]
port 422 nsew signal tristate
rlabel metal2 s 292854 159200 292910 160000 6 la_oenb[74]
port 423 nsew signal tristate
rlabel metal2 s 296718 159200 296774 160000 6 la_oenb[75]
port 424 nsew signal tristate
rlabel metal2 s 300674 159200 300730 160000 6 la_oenb[76]
port 425 nsew signal tristate
rlabel metal2 s 304538 159200 304594 160000 6 la_oenb[77]
port 426 nsew signal tristate
rlabel metal2 s 308494 159200 308550 160000 6 la_oenb[78]
port 427 nsew signal tristate
rlabel metal2 s 312358 159200 312414 160000 6 la_oenb[79]
port 428 nsew signal tristate
rlabel metal2 s 31666 159200 31722 160000 6 la_oenb[7]
port 429 nsew signal tristate
rlabel metal2 s 316222 159200 316278 160000 6 la_oenb[80]
port 430 nsew signal tristate
rlabel metal2 s 320178 159200 320234 160000 6 la_oenb[81]
port 431 nsew signal tristate
rlabel metal2 s 324042 159200 324098 160000 6 la_oenb[82]
port 432 nsew signal tristate
rlabel metal2 s 327906 159200 327962 160000 6 la_oenb[83]
port 433 nsew signal tristate
rlabel metal2 s 331862 159200 331918 160000 6 la_oenb[84]
port 434 nsew signal tristate
rlabel metal2 s 335726 159200 335782 160000 6 la_oenb[85]
port 435 nsew signal tristate
rlabel metal2 s 339682 159200 339738 160000 6 la_oenb[86]
port 436 nsew signal tristate
rlabel metal2 s 343546 159200 343602 160000 6 la_oenb[87]
port 437 nsew signal tristate
rlabel metal2 s 347410 159200 347466 160000 6 la_oenb[88]
port 438 nsew signal tristate
rlabel metal2 s 351366 159200 351422 160000 6 la_oenb[89]
port 439 nsew signal tristate
rlabel metal2 s 35530 159200 35586 160000 6 la_oenb[8]
port 440 nsew signal tristate
rlabel metal2 s 355230 159200 355286 160000 6 la_oenb[90]
port 441 nsew signal tristate
rlabel metal2 s 359094 159200 359150 160000 6 la_oenb[91]
port 442 nsew signal tristate
rlabel metal2 s 363050 159200 363106 160000 6 la_oenb[92]
port 443 nsew signal tristate
rlabel metal2 s 366914 159200 366970 160000 6 la_oenb[93]
port 444 nsew signal tristate
rlabel metal2 s 370870 159200 370926 160000 6 la_oenb[94]
port 445 nsew signal tristate
rlabel metal2 s 374734 159200 374790 160000 6 la_oenb[95]
port 446 nsew signal tristate
rlabel metal2 s 378598 159200 378654 160000 6 la_oenb[96]
port 447 nsew signal tristate
rlabel metal2 s 382554 159200 382610 160000 6 la_oenb[97]
port 448 nsew signal tristate
rlabel metal2 s 386418 159200 386474 160000 6 la_oenb[98]
port 449 nsew signal tristate
rlabel metal2 s 390282 159200 390338 160000 6 la_oenb[99]
port 450 nsew signal tristate
rlabel metal2 s 39394 159200 39450 160000 6 la_oenb[9]
port 451 nsew signal tristate
rlabel metal2 s 5262 159200 5318 160000 6 la_output[0]
port 452 nsew signal tristate
rlabel metal2 s 395158 159200 395214 160000 6 la_output[100]
port 453 nsew signal tristate
rlabel metal2 s 399114 159200 399170 160000 6 la_output[101]
port 454 nsew signal tristate
rlabel metal2 s 402978 159200 403034 160000 6 la_output[102]
port 455 nsew signal tristate
rlabel metal2 s 406934 159200 406990 160000 6 la_output[103]
port 456 nsew signal tristate
rlabel metal2 s 410798 159200 410854 160000 6 la_output[104]
port 457 nsew signal tristate
rlabel metal2 s 414662 159200 414718 160000 6 la_output[105]
port 458 nsew signal tristate
rlabel metal2 s 418618 159200 418674 160000 6 la_output[106]
port 459 nsew signal tristate
rlabel metal2 s 422482 159200 422538 160000 6 la_output[107]
port 460 nsew signal tristate
rlabel metal2 s 426346 159200 426402 160000 6 la_output[108]
port 461 nsew signal tristate
rlabel metal2 s 430302 159200 430358 160000 6 la_output[109]
port 462 nsew signal tristate
rlabel metal2 s 44270 159200 44326 160000 6 la_output[10]
port 463 nsew signal tristate
rlabel metal2 s 434166 159200 434222 160000 6 la_output[110]
port 464 nsew signal tristate
rlabel metal2 s 438122 159200 438178 160000 6 la_output[111]
port 465 nsew signal tristate
rlabel metal2 s 441986 159200 442042 160000 6 la_output[112]
port 466 nsew signal tristate
rlabel metal2 s 445850 159200 445906 160000 6 la_output[113]
port 467 nsew signal tristate
rlabel metal2 s 449806 159200 449862 160000 6 la_output[114]
port 468 nsew signal tristate
rlabel metal2 s 453670 159200 453726 160000 6 la_output[115]
port 469 nsew signal tristate
rlabel metal2 s 457626 159200 457682 160000 6 la_output[116]
port 470 nsew signal tristate
rlabel metal2 s 461490 159200 461546 160000 6 la_output[117]
port 471 nsew signal tristate
rlabel metal2 s 465354 159200 465410 160000 6 la_output[118]
port 472 nsew signal tristate
rlabel metal2 s 469310 159200 469366 160000 6 la_output[119]
port 473 nsew signal tristate
rlabel metal2 s 48226 159200 48282 160000 6 la_output[11]
port 474 nsew signal tristate
rlabel metal2 s 473174 159200 473230 160000 6 la_output[120]
port 475 nsew signal tristate
rlabel metal2 s 477038 159200 477094 160000 6 la_output[121]
port 476 nsew signal tristate
rlabel metal2 s 480994 159200 481050 160000 6 la_output[122]
port 477 nsew signal tristate
rlabel metal2 s 484858 159200 484914 160000 6 la_output[123]
port 478 nsew signal tristate
rlabel metal2 s 488814 159200 488870 160000 6 la_output[124]
port 479 nsew signal tristate
rlabel metal2 s 492678 159200 492734 160000 6 la_output[125]
port 480 nsew signal tristate
rlabel metal2 s 496542 159200 496598 160000 6 la_output[126]
port 481 nsew signal tristate
rlabel metal2 s 500498 159200 500554 160000 6 la_output[127]
port 482 nsew signal tristate
rlabel metal2 s 52090 159200 52146 160000 6 la_output[12]
port 483 nsew signal tristate
rlabel metal2 s 55954 159200 56010 160000 6 la_output[13]
port 484 nsew signal tristate
rlabel metal2 s 59910 159200 59966 160000 6 la_output[14]
port 485 nsew signal tristate
rlabel metal2 s 63774 159200 63830 160000 6 la_output[15]
port 486 nsew signal tristate
rlabel metal2 s 67730 159200 67786 160000 6 la_output[16]
port 487 nsew signal tristate
rlabel metal2 s 71594 159200 71650 160000 6 la_output[17]
port 488 nsew signal tristate
rlabel metal2 s 75458 159200 75514 160000 6 la_output[18]
port 489 nsew signal tristate
rlabel metal2 s 79414 159200 79470 160000 6 la_output[19]
port 490 nsew signal tristate
rlabel metal2 s 9218 159200 9274 160000 6 la_output[1]
port 491 nsew signal tristate
rlabel metal2 s 83278 159200 83334 160000 6 la_output[20]
port 492 nsew signal tristate
rlabel metal2 s 87142 159200 87198 160000 6 la_output[21]
port 493 nsew signal tristate
rlabel metal2 s 91098 159200 91154 160000 6 la_output[22]
port 494 nsew signal tristate
rlabel metal2 s 94962 159200 95018 160000 6 la_output[23]
port 495 nsew signal tristate
rlabel metal2 s 98918 159200 98974 160000 6 la_output[24]
port 496 nsew signal tristate
rlabel metal2 s 102782 159200 102838 160000 6 la_output[25]
port 497 nsew signal tristate
rlabel metal2 s 106646 159200 106702 160000 6 la_output[26]
port 498 nsew signal tristate
rlabel metal2 s 110602 159200 110658 160000 6 la_output[27]
port 499 nsew signal tristate
rlabel metal2 s 114466 159200 114522 160000 6 la_output[28]
port 500 nsew signal tristate
rlabel metal2 s 118330 159200 118386 160000 6 la_output[29]
port 501 nsew signal tristate
rlabel metal2 s 13082 159200 13138 160000 6 la_output[2]
port 502 nsew signal tristate
rlabel metal2 s 122286 159200 122342 160000 6 la_output[30]
port 503 nsew signal tristate
rlabel metal2 s 126150 159200 126206 160000 6 la_output[31]
port 504 nsew signal tristate
rlabel metal2 s 130106 159200 130162 160000 6 la_output[32]
port 505 nsew signal tristate
rlabel metal2 s 133970 159200 134026 160000 6 la_output[33]
port 506 nsew signal tristate
rlabel metal2 s 137834 159200 137890 160000 6 la_output[34]
port 507 nsew signal tristate
rlabel metal2 s 141790 159200 141846 160000 6 la_output[35]
port 508 nsew signal tristate
rlabel metal2 s 145654 159200 145710 160000 6 la_output[36]
port 509 nsew signal tristate
rlabel metal2 s 149610 159200 149666 160000 6 la_output[37]
port 510 nsew signal tristate
rlabel metal2 s 153474 159200 153530 160000 6 la_output[38]
port 511 nsew signal tristate
rlabel metal2 s 157338 159200 157394 160000 6 la_output[39]
port 512 nsew signal tristate
rlabel metal2 s 17038 159200 17094 160000 6 la_output[3]
port 513 nsew signal tristate
rlabel metal2 s 161294 159200 161350 160000 6 la_output[40]
port 514 nsew signal tristate
rlabel metal2 s 165158 159200 165214 160000 6 la_output[41]
port 515 nsew signal tristate
rlabel metal2 s 169022 159200 169078 160000 6 la_output[42]
port 516 nsew signal tristate
rlabel metal2 s 172978 159200 173034 160000 6 la_output[43]
port 517 nsew signal tristate
rlabel metal2 s 176842 159200 176898 160000 6 la_output[44]
port 518 nsew signal tristate
rlabel metal2 s 180798 159200 180854 160000 6 la_output[45]
port 519 nsew signal tristate
rlabel metal2 s 184662 159200 184718 160000 6 la_output[46]
port 520 nsew signal tristate
rlabel metal2 s 188526 159200 188582 160000 6 la_output[47]
port 521 nsew signal tristate
rlabel metal2 s 192482 159200 192538 160000 6 la_output[48]
port 522 nsew signal tristate
rlabel metal2 s 196346 159200 196402 160000 6 la_output[49]
port 523 nsew signal tristate
rlabel metal2 s 20902 159200 20958 160000 6 la_output[4]
port 524 nsew signal tristate
rlabel metal2 s 200210 159200 200266 160000 6 la_output[50]
port 525 nsew signal tristate
rlabel metal2 s 204166 159200 204222 160000 6 la_output[51]
port 526 nsew signal tristate
rlabel metal2 s 208030 159200 208086 160000 6 la_output[52]
port 527 nsew signal tristate
rlabel metal2 s 211986 159200 212042 160000 6 la_output[53]
port 528 nsew signal tristate
rlabel metal2 s 215850 159200 215906 160000 6 la_output[54]
port 529 nsew signal tristate
rlabel metal2 s 219714 159200 219770 160000 6 la_output[55]
port 530 nsew signal tristate
rlabel metal2 s 223670 159200 223726 160000 6 la_output[56]
port 531 nsew signal tristate
rlabel metal2 s 227534 159200 227590 160000 6 la_output[57]
port 532 nsew signal tristate
rlabel metal2 s 231490 159200 231546 160000 6 la_output[58]
port 533 nsew signal tristate
rlabel metal2 s 235354 159200 235410 160000 6 la_output[59]
port 534 nsew signal tristate
rlabel metal2 s 24766 159200 24822 160000 6 la_output[5]
port 535 nsew signal tristate
rlabel metal2 s 239218 159200 239274 160000 6 la_output[60]
port 536 nsew signal tristate
rlabel metal2 s 243174 159200 243230 160000 6 la_output[61]
port 537 nsew signal tristate
rlabel metal2 s 247038 159200 247094 160000 6 la_output[62]
port 538 nsew signal tristate
rlabel metal2 s 250902 159200 250958 160000 6 la_output[63]
port 539 nsew signal tristate
rlabel metal2 s 254858 159200 254914 160000 6 la_output[64]
port 540 nsew signal tristate
rlabel metal2 s 258722 159200 258778 160000 6 la_output[65]
port 541 nsew signal tristate
rlabel metal2 s 262678 159200 262734 160000 6 la_output[66]
port 542 nsew signal tristate
rlabel metal2 s 266542 159200 266598 160000 6 la_output[67]
port 543 nsew signal tristate
rlabel metal2 s 270406 159200 270462 160000 6 la_output[68]
port 544 nsew signal tristate
rlabel metal2 s 274362 159200 274418 160000 6 la_output[69]
port 545 nsew signal tristate
rlabel metal2 s 28722 159200 28778 160000 6 la_output[6]
port 546 nsew signal tristate
rlabel metal2 s 278226 159200 278282 160000 6 la_output[70]
port 547 nsew signal tristate
rlabel metal2 s 282090 159200 282146 160000 6 la_output[71]
port 548 nsew signal tristate
rlabel metal2 s 286046 159200 286102 160000 6 la_output[72]
port 549 nsew signal tristate
rlabel metal2 s 289910 159200 289966 160000 6 la_output[73]
port 550 nsew signal tristate
rlabel metal2 s 293866 159200 293922 160000 6 la_output[74]
port 551 nsew signal tristate
rlabel metal2 s 297730 159200 297786 160000 6 la_output[75]
port 552 nsew signal tristate
rlabel metal2 s 301594 159200 301650 160000 6 la_output[76]
port 553 nsew signal tristate
rlabel metal2 s 305550 159200 305606 160000 6 la_output[77]
port 554 nsew signal tristate
rlabel metal2 s 309414 159200 309470 160000 6 la_output[78]
port 555 nsew signal tristate
rlabel metal2 s 313278 159200 313334 160000 6 la_output[79]
port 556 nsew signal tristate
rlabel metal2 s 32586 159200 32642 160000 6 la_output[7]
port 557 nsew signal tristate
rlabel metal2 s 317234 159200 317290 160000 6 la_output[80]
port 558 nsew signal tristate
rlabel metal2 s 321098 159200 321154 160000 6 la_output[81]
port 559 nsew signal tristate
rlabel metal2 s 325054 159200 325110 160000 6 la_output[82]
port 560 nsew signal tristate
rlabel metal2 s 328918 159200 328974 160000 6 la_output[83]
port 561 nsew signal tristate
rlabel metal2 s 332782 159200 332838 160000 6 la_output[84]
port 562 nsew signal tristate
rlabel metal2 s 336738 159200 336794 160000 6 la_output[85]
port 563 nsew signal tristate
rlabel metal2 s 340602 159200 340658 160000 6 la_output[86]
port 564 nsew signal tristate
rlabel metal2 s 344558 159200 344614 160000 6 la_output[87]
port 565 nsew signal tristate
rlabel metal2 s 348422 159200 348478 160000 6 la_output[88]
port 566 nsew signal tristate
rlabel metal2 s 352286 159200 352342 160000 6 la_output[89]
port 567 nsew signal tristate
rlabel metal2 s 36542 159200 36598 160000 6 la_output[8]
port 568 nsew signal tristate
rlabel metal2 s 356242 159200 356298 160000 6 la_output[90]
port 569 nsew signal tristate
rlabel metal2 s 360106 159200 360162 160000 6 la_output[91]
port 570 nsew signal tristate
rlabel metal2 s 363970 159200 364026 160000 6 la_output[92]
port 571 nsew signal tristate
rlabel metal2 s 367926 159200 367982 160000 6 la_output[93]
port 572 nsew signal tristate
rlabel metal2 s 371790 159200 371846 160000 6 la_output[94]
port 573 nsew signal tristate
rlabel metal2 s 375746 159200 375802 160000 6 la_output[95]
port 574 nsew signal tristate
rlabel metal2 s 379610 159200 379666 160000 6 la_output[96]
port 575 nsew signal tristate
rlabel metal2 s 383474 159200 383530 160000 6 la_output[97]
port 576 nsew signal tristate
rlabel metal2 s 387430 159200 387486 160000 6 la_output[98]
port 577 nsew signal tristate
rlabel metal2 s 391294 159200 391350 160000 6 la_output[99]
port 578 nsew signal tristate
rlabel metal2 s 40406 159200 40462 160000 6 la_output[9]
port 579 nsew signal tristate
rlabel metal3 s 0 157496 800 157616 6 mprj_ack_i
port 580 nsew signal input
rlabel metal2 s 504362 159200 504418 160000 6 mprj_adr_o[0]
port 581 nsew signal tristate
rlabel metal2 s 527730 159200 527786 160000 6 mprj_adr_o[10]
port 582 nsew signal tristate
rlabel metal2 s 529754 159200 529810 160000 6 mprj_adr_o[11]
port 583 nsew signal tristate
rlabel metal2 s 531686 159200 531742 160000 6 mprj_adr_o[12]
port 584 nsew signal tristate
rlabel metal2 s 533618 159200 533674 160000 6 mprj_adr_o[13]
port 585 nsew signal tristate
rlabel metal2 s 535550 159200 535606 160000 6 mprj_adr_o[14]
port 586 nsew signal tristate
rlabel metal2 s 537482 159200 537538 160000 6 mprj_adr_o[15]
port 587 nsew signal tristate
rlabel metal2 s 539506 159200 539562 160000 6 mprj_adr_o[16]
port 588 nsew signal tristate
rlabel metal2 s 541438 159200 541494 160000 6 mprj_adr_o[17]
port 589 nsew signal tristate
rlabel metal2 s 543370 159200 543426 160000 6 mprj_adr_o[18]
port 590 nsew signal tristate
rlabel metal2 s 545302 159200 545358 160000 6 mprj_adr_o[19]
port 591 nsew signal tristate
rlabel metal2 s 507306 159200 507362 160000 6 mprj_adr_o[1]
port 592 nsew signal tristate
rlabel metal2 s 547234 159200 547290 160000 6 mprj_adr_o[20]
port 593 nsew signal tristate
rlabel metal2 s 549166 159200 549222 160000 6 mprj_adr_o[21]
port 594 nsew signal tristate
rlabel metal2 s 551190 159200 551246 160000 6 mprj_adr_o[22]
port 595 nsew signal tristate
rlabel metal2 s 553122 159200 553178 160000 6 mprj_adr_o[23]
port 596 nsew signal tristate
rlabel metal2 s 555054 159200 555110 160000 6 mprj_adr_o[24]
port 597 nsew signal tristate
rlabel metal2 s 556986 159200 557042 160000 6 mprj_adr_o[25]
port 598 nsew signal tristate
rlabel metal2 s 558918 159200 558974 160000 6 mprj_adr_o[26]
port 599 nsew signal tristate
rlabel metal2 s 560942 159200 560998 160000 6 mprj_adr_o[27]
port 600 nsew signal tristate
rlabel metal2 s 562874 159200 562930 160000 6 mprj_adr_o[28]
port 601 nsew signal tristate
rlabel metal2 s 564806 159200 564862 160000 6 mprj_adr_o[29]
port 602 nsew signal tristate
rlabel metal2 s 510250 159200 510306 160000 6 mprj_adr_o[2]
port 603 nsew signal tristate
rlabel metal2 s 566738 159200 566794 160000 6 mprj_adr_o[30]
port 604 nsew signal tristate
rlabel metal2 s 568670 159200 568726 160000 6 mprj_adr_o[31]
port 605 nsew signal tristate
rlabel metal2 s 513102 159200 513158 160000 6 mprj_adr_o[3]
port 606 nsew signal tristate
rlabel metal2 s 516046 159200 516102 160000 6 mprj_adr_o[4]
port 607 nsew signal tristate
rlabel metal2 s 517978 159200 518034 160000 6 mprj_adr_o[5]
port 608 nsew signal tristate
rlabel metal2 s 520002 159200 520058 160000 6 mprj_adr_o[6]
port 609 nsew signal tristate
rlabel metal2 s 521934 159200 521990 160000 6 mprj_adr_o[7]
port 610 nsew signal tristate
rlabel metal2 s 523866 159200 523922 160000 6 mprj_adr_o[8]
port 611 nsew signal tristate
rlabel metal2 s 525798 159200 525854 160000 6 mprj_adr_o[9]
port 612 nsew signal tristate
rlabel metal2 s 501418 159200 501474 160000 6 mprj_cyc_o
port 613 nsew signal tristate
rlabel metal3 s 0 11296 800 11416 6 mprj_dat_i[0]
port 614 nsew signal input
rlabel metal3 s 0 56992 800 57112 6 mprj_dat_i[10]
port 615 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 mprj_dat_i[11]
port 616 nsew signal input
rlabel metal3 s 0 66104 800 66224 6 mprj_dat_i[12]
port 617 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 mprj_dat_i[13]
port 618 nsew signal input
rlabel metal3 s 0 75216 800 75336 6 mprj_dat_i[14]
port 619 nsew signal input
rlabel metal3 s 0 79840 800 79960 6 mprj_dat_i[15]
port 620 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 mprj_dat_i[16]
port 621 nsew signal input
rlabel metal3 s 0 88952 800 89072 6 mprj_dat_i[17]
port 622 nsew signal input
rlabel metal3 s 0 93576 800 93696 6 mprj_dat_i[18]
port 623 nsew signal input
rlabel metal3 s 0 98064 800 98184 6 mprj_dat_i[19]
port 624 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 mprj_dat_i[1]
port 625 nsew signal input
rlabel metal3 s 0 102688 800 102808 6 mprj_dat_i[20]
port 626 nsew signal input
rlabel metal3 s 0 107176 800 107296 6 mprj_dat_i[21]
port 627 nsew signal input
rlabel metal3 s 0 111800 800 111920 6 mprj_dat_i[22]
port 628 nsew signal input
rlabel metal3 s 0 116424 800 116544 6 mprj_dat_i[23]
port 629 nsew signal input
rlabel metal3 s 0 120912 800 121032 6 mprj_dat_i[24]
port 630 nsew signal input
rlabel metal3 s 0 125536 800 125656 6 mprj_dat_i[25]
port 631 nsew signal input
rlabel metal3 s 0 130024 800 130144 6 mprj_dat_i[26]
port 632 nsew signal input
rlabel metal3 s 0 134648 800 134768 6 mprj_dat_i[27]
port 633 nsew signal input
rlabel metal3 s 0 139272 800 139392 6 mprj_dat_i[28]
port 634 nsew signal input
rlabel metal3 s 0 143760 800 143880 6 mprj_dat_i[29]
port 635 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 mprj_dat_i[2]
port 636 nsew signal input
rlabel metal3 s 0 148384 800 148504 6 mprj_dat_i[30]
port 637 nsew signal input
rlabel metal3 s 0 152872 800 152992 6 mprj_dat_i[31]
port 638 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 mprj_dat_i[3]
port 639 nsew signal input
rlabel metal3 s 0 29520 800 29640 6 mprj_dat_i[4]
port 640 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 mprj_dat_i[5]
port 641 nsew signal input
rlabel metal3 s 0 38632 800 38752 6 mprj_dat_i[6]
port 642 nsew signal input
rlabel metal3 s 0 43256 800 43376 6 mprj_dat_i[7]
port 643 nsew signal input
rlabel metal3 s 0 47880 800 48000 6 mprj_dat_i[8]
port 644 nsew signal input
rlabel metal3 s 0 52368 800 52488 6 mprj_dat_i[9]
port 645 nsew signal input
rlabel metal2 s 505374 159200 505430 160000 6 mprj_dat_o[0]
port 646 nsew signal tristate
rlabel metal2 s 528742 159200 528798 160000 6 mprj_dat_o[10]
port 647 nsew signal tristate
rlabel metal2 s 530674 159200 530730 160000 6 mprj_dat_o[11]
port 648 nsew signal tristate
rlabel metal2 s 532606 159200 532662 160000 6 mprj_dat_o[12]
port 649 nsew signal tristate
rlabel metal2 s 534630 159200 534686 160000 6 mprj_dat_o[13]
port 650 nsew signal tristate
rlabel metal2 s 536562 159200 536618 160000 6 mprj_dat_o[14]
port 651 nsew signal tristate
rlabel metal2 s 538494 159200 538550 160000 6 mprj_dat_o[15]
port 652 nsew signal tristate
rlabel metal2 s 540426 159200 540482 160000 6 mprj_dat_o[16]
port 653 nsew signal tristate
rlabel metal2 s 542358 159200 542414 160000 6 mprj_dat_o[17]
port 654 nsew signal tristate
rlabel metal2 s 544290 159200 544346 160000 6 mprj_dat_o[18]
port 655 nsew signal tristate
rlabel metal2 s 546314 159200 546370 160000 6 mprj_dat_o[19]
port 656 nsew signal tristate
rlabel metal2 s 508226 159200 508282 160000 6 mprj_dat_o[1]
port 657 nsew signal tristate
rlabel metal2 s 548246 159200 548302 160000 6 mprj_dat_o[20]
port 658 nsew signal tristate
rlabel metal2 s 550178 159200 550234 160000 6 mprj_dat_o[21]
port 659 nsew signal tristate
rlabel metal2 s 552110 159200 552166 160000 6 mprj_dat_o[22]
port 660 nsew signal tristate
rlabel metal2 s 554042 159200 554098 160000 6 mprj_dat_o[23]
port 661 nsew signal tristate
rlabel metal2 s 556066 159200 556122 160000 6 mprj_dat_o[24]
port 662 nsew signal tristate
rlabel metal2 s 557998 159200 558054 160000 6 mprj_dat_o[25]
port 663 nsew signal tristate
rlabel metal2 s 559930 159200 559986 160000 6 mprj_dat_o[26]
port 664 nsew signal tristate
rlabel metal2 s 561862 159200 561918 160000 6 mprj_dat_o[27]
port 665 nsew signal tristate
rlabel metal2 s 563794 159200 563850 160000 6 mprj_dat_o[28]
port 666 nsew signal tristate
rlabel metal2 s 565818 159200 565874 160000 6 mprj_dat_o[29]
port 667 nsew signal tristate
rlabel metal2 s 511170 159200 511226 160000 6 mprj_dat_o[2]
port 668 nsew signal tristate
rlabel metal2 s 567750 159200 567806 160000 6 mprj_dat_o[30]
port 669 nsew signal tristate
rlabel metal2 s 569682 159200 569738 160000 6 mprj_dat_o[31]
port 670 nsew signal tristate
rlabel metal2 s 514114 159200 514170 160000 6 mprj_dat_o[3]
port 671 nsew signal tristate
rlabel metal2 s 517058 159200 517114 160000 6 mprj_dat_o[4]
port 672 nsew signal tristate
rlabel metal2 s 518990 159200 519046 160000 6 mprj_dat_o[5]
port 673 nsew signal tristate
rlabel metal2 s 520922 159200 520978 160000 6 mprj_dat_o[6]
port 674 nsew signal tristate
rlabel metal2 s 522854 159200 522910 160000 6 mprj_dat_o[7]
port 675 nsew signal tristate
rlabel metal2 s 524878 159200 524934 160000 6 mprj_dat_o[8]
port 676 nsew signal tristate
rlabel metal2 s 526810 159200 526866 160000 6 mprj_dat_o[9]
port 677 nsew signal tristate
rlabel metal2 s 506294 159200 506350 160000 6 mprj_sel_o[0]
port 678 nsew signal tristate
rlabel metal2 s 509238 159200 509294 160000 6 mprj_sel_o[1]
port 679 nsew signal tristate
rlabel metal2 s 512182 159200 512238 160000 6 mprj_sel_o[2]
port 680 nsew signal tristate
rlabel metal2 s 515126 159200 515182 160000 6 mprj_sel_o[3]
port 681 nsew signal tristate
rlabel metal2 s 502430 159200 502486 160000 6 mprj_stb_o
port 682 nsew signal tristate
rlabel metal2 s 570694 159200 570750 160000 6 mprj_wb_iena
port 683 nsew signal tristate
rlabel metal2 s 503350 159200 503406 160000 6 mprj_we_o
port 684 nsew signal tristate
rlabel metal2 s 98366 0 98422 800 6 qspi_enabled
port 685 nsew signal tristate
rlabel metal2 s 577226 0 577282 800 6 ser_rx
port 686 nsew signal input
rlabel metal2 s 566554 0 566610 800 6 ser_tx
port 687 nsew signal tristate
rlabel metal2 s 529294 0 529350 800 6 spi_csb
port 688 nsew signal tristate
rlabel metal2 s 534630 0 534686 800 6 spi_enabled
port 689 nsew signal tristate
rlabel metal2 s 539966 0 540022 800 6 spi_sck
port 690 nsew signal tristate
rlabel metal2 s 545302 0 545358 800 6 spi_sdi
port 691 nsew signal input
rlabel metal2 s 550546 0 550602 800 6 spi_sdo
port 692 nsew signal tristate
rlabel metal2 s 555882 0 555938 800 6 spi_sdoenb
port 693 nsew signal tristate
rlabel metal2 s 295154 0 295210 800 6 sram_ro_addr[0]
port 694 nsew signal input
rlabel metal2 s 300490 0 300546 800 6 sram_ro_addr[1]
port 695 nsew signal input
rlabel metal2 s 305826 0 305882 800 6 sram_ro_addr[2]
port 696 nsew signal input
rlabel metal2 s 311162 0 311218 800 6 sram_ro_addr[3]
port 697 nsew signal input
rlabel metal2 s 316498 0 316554 800 6 sram_ro_addr[4]
port 698 nsew signal input
rlabel metal2 s 321834 0 321890 800 6 sram_ro_addr[5]
port 699 nsew signal input
rlabel metal2 s 327078 0 327134 800 6 sram_ro_addr[6]
port 700 nsew signal input
rlabel metal2 s 332414 0 332470 800 6 sram_ro_addr[7]
port 701 nsew signal input
rlabel metal2 s 284574 0 284630 800 6 sram_ro_clk
port 702 nsew signal input
rlabel metal2 s 289910 0 289966 800 6 sram_ro_csb
port 703 nsew signal input
rlabel metal2 s 337750 0 337806 800 6 sram_ro_data[0]
port 704 nsew signal tristate
rlabel metal2 s 390926 0 390982 800 6 sram_ro_data[10]
port 705 nsew signal tristate
rlabel metal2 s 396262 0 396318 800 6 sram_ro_data[11]
port 706 nsew signal tristate
rlabel metal2 s 401598 0 401654 800 6 sram_ro_data[12]
port 707 nsew signal tristate
rlabel metal2 s 406934 0 406990 800 6 sram_ro_data[13]
port 708 nsew signal tristate
rlabel metal2 s 412270 0 412326 800 6 sram_ro_data[14]
port 709 nsew signal tristate
rlabel metal2 s 417606 0 417662 800 6 sram_ro_data[15]
port 710 nsew signal tristate
rlabel metal2 s 422850 0 422906 800 6 sram_ro_data[16]
port 711 nsew signal tristate
rlabel metal2 s 428186 0 428242 800 6 sram_ro_data[17]
port 712 nsew signal tristate
rlabel metal2 s 433522 0 433578 800 6 sram_ro_data[18]
port 713 nsew signal tristate
rlabel metal2 s 438858 0 438914 800 6 sram_ro_data[19]
port 714 nsew signal tristate
rlabel metal2 s 343086 0 343142 800 6 sram_ro_data[1]
port 715 nsew signal tristate
rlabel metal2 s 444194 0 444250 800 6 sram_ro_data[20]
port 716 nsew signal tristate
rlabel metal2 s 449530 0 449586 800 6 sram_ro_data[21]
port 717 nsew signal tristate
rlabel metal2 s 454774 0 454830 800 6 sram_ro_data[22]
port 718 nsew signal tristate
rlabel metal2 s 460110 0 460166 800 6 sram_ro_data[23]
port 719 nsew signal tristate
rlabel metal2 s 465446 0 465502 800 6 sram_ro_data[24]
port 720 nsew signal tristate
rlabel metal2 s 470782 0 470838 800 6 sram_ro_data[25]
port 721 nsew signal tristate
rlabel metal2 s 476118 0 476174 800 6 sram_ro_data[26]
port 722 nsew signal tristate
rlabel metal2 s 481454 0 481510 800 6 sram_ro_data[27]
port 723 nsew signal tristate
rlabel metal2 s 486698 0 486754 800 6 sram_ro_data[28]
port 724 nsew signal tristate
rlabel metal2 s 492034 0 492090 800 6 sram_ro_data[29]
port 725 nsew signal tristate
rlabel metal2 s 348422 0 348478 800 6 sram_ro_data[2]
port 726 nsew signal tristate
rlabel metal2 s 497370 0 497426 800 6 sram_ro_data[30]
port 727 nsew signal tristate
rlabel metal2 s 502706 0 502762 800 6 sram_ro_data[31]
port 728 nsew signal tristate
rlabel metal2 s 353758 0 353814 800 6 sram_ro_data[3]
port 729 nsew signal tristate
rlabel metal2 s 359002 0 359058 800 6 sram_ro_data[4]
port 730 nsew signal tristate
rlabel metal2 s 364338 0 364394 800 6 sram_ro_data[5]
port 731 nsew signal tristate
rlabel metal2 s 369674 0 369730 800 6 sram_ro_data[6]
port 732 nsew signal tristate
rlabel metal2 s 375010 0 375066 800 6 sram_ro_data[7]
port 733 nsew signal tristate
rlabel metal2 s 380346 0 380402 800 6 sram_ro_data[8]
port 734 nsew signal tristate
rlabel metal2 s 385682 0 385738 800 6 sram_ro_data[9]
port 735 nsew signal tristate
rlabel metal2 s 561218 0 561274 800 6 trap
port 736 nsew signal tristate
rlabel metal2 s 571890 0 571946 800 6 uart_enabled
port 737 nsew signal tristate
rlabel metal2 s 571614 159200 571670 160000 6 user_irq_ena[0]
port 738 nsew signal tristate
rlabel metal2 s 572626 159200 572682 160000 6 user_irq_ena[1]
port 739 nsew signal tristate
rlabel metal2 s 573546 159200 573602 160000 6 user_irq_ena[2]
port 740 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 580000 160000
<< end >>
